magic
tech sky130A
timestamp 1730994170
<< metal1 >>
rect 6400 12130 10050 12150
rect 6400 12070 9670 12130
rect 9730 12070 9770 12130
rect 9830 12070 9870 12130
rect 9930 12070 9970 12130
rect 10030 12070 10050 12130
rect 6400 12050 10050 12070
<< via1 >>
rect 9670 12070 9730 12130
rect 9770 12070 9830 12130
rect 9870 12070 9930 12130
rect 9970 12070 10030 12130
<< metal2 >>
rect 6900 12630 7000 12650
rect 6900 12570 6920 12630
rect 6980 12570 7000 12630
rect 6900 12530 7000 12570
rect 6900 12470 6920 12530
rect 6980 12470 7000 12530
rect 6900 12430 7000 12470
rect 6900 12370 6920 12430
rect 6980 12370 7000 12430
rect 6900 12330 7000 12370
rect 6900 12270 6920 12330
rect 6980 12270 7000 12330
rect 6900 12250 7000 12270
rect 7100 12630 7200 12650
rect 7100 12570 7120 12630
rect 7180 12570 7200 12630
rect 7100 12530 7200 12570
rect 7100 12470 7120 12530
rect 7180 12470 7200 12530
rect 7100 12430 7200 12470
rect 7100 12370 7120 12430
rect 7180 12370 7200 12430
rect 7100 12330 7200 12370
rect 7100 12270 7120 12330
rect 7180 12270 7200 12330
rect 7100 12250 7200 12270
rect 9650 12130 10050 12150
rect 9650 12070 9670 12130
rect 9730 12070 9770 12130
rect 9830 12070 9870 12130
rect 9930 12070 9970 12130
rect 10030 12070 10050 12130
rect 9650 12050 10050 12070
rect 9450 11730 10050 11750
rect 9450 11670 9670 11730
rect 9730 11670 9770 11730
rect 9830 11670 9870 11730
rect 9930 11670 9970 11730
rect 10030 11670 10050 11730
rect 9450 11650 10050 11670
rect 9500 11480 10050 11500
rect 9500 11420 9670 11480
rect 9730 11420 9770 11480
rect 9830 11420 9870 11480
rect 9930 11420 9970 11480
rect 10030 11420 10050 11480
rect 9500 11400 10050 11420
<< via2 >>
rect 6920 12570 6980 12630
rect 6920 12470 6980 12530
rect 6920 12370 6980 12430
rect 6920 12270 6980 12330
rect 7120 12570 7180 12630
rect 7120 12470 7180 12530
rect 7120 12370 7180 12430
rect 7120 12270 7180 12330
rect 9670 12070 9730 12130
rect 9770 12070 9830 12130
rect 9870 12070 9930 12130
rect 9970 12070 10030 12130
rect 9670 11670 9730 11730
rect 9770 11670 9830 11730
rect 9870 11670 9930 11730
rect 9970 11670 10030 11730
rect 9670 11420 9730 11480
rect 9770 11420 9830 11480
rect 9870 11420 9930 11480
rect 9970 11420 10030 11480
<< metal3 >>
rect 6900 12630 7000 12650
rect 6900 12570 6920 12630
rect 6980 12570 7000 12630
rect 6900 12530 7000 12570
rect 6900 12470 6920 12530
rect 6980 12470 7000 12530
rect 6900 12430 7000 12470
rect 6900 12370 6920 12430
rect 6980 12370 7000 12430
rect 6900 12330 7000 12370
rect 6900 12270 6920 12330
rect 6980 12270 7000 12330
rect 6900 12250 7000 12270
rect 7100 12630 7200 12650
rect 7100 12570 7120 12630
rect 7180 12570 7200 12630
rect 7100 12530 7200 12570
rect 7100 12470 7120 12530
rect 7180 12470 7200 12530
rect 7100 12430 7200 12470
rect 7100 12370 7120 12430
rect 7180 12370 7200 12430
rect 7100 12330 7200 12370
rect 7100 12270 7120 12330
rect 7180 12270 7200 12330
rect 7100 12250 7200 12270
rect 9650 12130 10050 12150
rect 9650 12070 9670 12130
rect 9730 12070 9770 12130
rect 9830 12070 9870 12130
rect 9930 12070 9970 12130
rect 10030 12070 10050 12130
rect 9650 12050 10050 12070
rect 9650 11730 10050 11750
rect 9650 11670 9670 11730
rect 9730 11670 9770 11730
rect 9830 11670 9870 11730
rect 9930 11670 9970 11730
rect 10030 11670 10050 11730
rect 9650 11650 10050 11670
rect 100 11450 300 11500
rect 100 11350 150 11450
rect 250 11350 300 11450
rect 9650 11480 10050 11500
rect 9650 11420 9670 11480
rect 9730 11420 9770 11480
rect 9830 11420 9870 11480
rect 9930 11420 9970 11480
rect 10030 11420 10050 11480
rect 9650 11400 10050 11420
rect 100 11250 300 11350
rect 100 11150 150 11250
rect 250 11200 300 11250
rect 250 11150 1600 11200
rect 100 11050 850 11150
rect 950 11050 1050 11150
rect 1150 11050 1250 11150
rect 1350 11050 1450 11150
rect 1550 11050 1600 11150
rect 100 10950 150 11050
rect 250 11000 1600 11050
rect 250 10950 300 11000
rect 100 10850 300 10950
rect 100 10750 150 10850
rect 250 10750 300 10850
rect 100 10700 300 10750
<< via3 >>
rect 6920 12570 6980 12630
rect 6920 12470 6980 12530
rect 6920 12370 6980 12430
rect 6920 12270 6980 12330
rect 7120 12570 7180 12630
rect 7120 12470 7180 12530
rect 7120 12370 7180 12430
rect 7120 12270 7180 12330
rect 9670 12070 9730 12130
rect 9770 12070 9830 12130
rect 9870 12070 9930 12130
rect 9970 12070 10030 12130
rect 9670 11670 9730 11730
rect 9770 11670 9830 11730
rect 9870 11670 9930 11730
rect 9970 11670 10030 11730
rect 150 11350 250 11450
rect 9670 11420 9730 11480
rect 9770 11420 9830 11480
rect 9870 11420 9930 11480
rect 9970 11420 10030 11480
rect 150 11150 250 11250
rect 850 11050 950 11150
rect 1050 11050 1150 11150
rect 1250 11050 1350 11150
rect 1450 11050 1550 11150
rect 150 10950 250 11050
rect 150 10750 250 10850
<< metal4 >>
rect 3067 22476 3097 22576
rect 3343 22476 3373 22576
rect 3619 22476 3649 22576
rect 3895 22476 3925 22576
rect 4171 22476 4201 22576
rect 4447 22476 4477 22576
rect 4723 22476 4753 22576
rect 4999 22476 5029 22576
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22476 6961 22576
rect 7207 22476 7237 22576
rect 7483 22476 7513 22576
rect 7759 22476 7789 22576
rect 8035 22476 8065 22576
rect 8311 22476 8341 22576
rect 8587 22476 8617 22576
rect 8863 22476 8893 22576
rect 9139 22500 9169 22576
rect 9415 22500 9445 22576
rect 100 11450 300 22076
rect 100 11350 150 11450
rect 250 11350 300 11450
rect 100 11250 300 11350
rect 100 11150 150 11250
rect 250 11150 300 11250
rect 100 11050 300 11150
rect 100 10950 150 11050
rect 250 10950 300 11050
rect 100 10850 300 10950
rect 100 10750 150 10850
rect 250 10750 300 10850
rect 100 500 300 10750
rect 400 12100 600 22076
rect 9050 13150 9200 22500
rect 6900 13000 9200 13150
rect 6900 12630 7000 13000
rect 9350 12850 9500 22500
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22480 13861 22576
rect 13825 22450 13870 22480
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 6900 12570 6920 12630
rect 6980 12570 7000 12630
rect 6900 12530 7000 12570
rect 6900 12470 6920 12530
rect 6980 12470 7000 12530
rect 6900 12430 7000 12470
rect 6900 12370 6920 12430
rect 6980 12370 7000 12430
rect 6900 12330 7000 12370
rect 6900 12270 6920 12330
rect 6980 12270 7000 12330
rect 6900 12250 7000 12270
rect 7100 12700 9500 12850
rect 7100 12630 7200 12700
rect 7100 12570 7120 12630
rect 7180 12570 7200 12630
rect 7100 12530 7200 12570
rect 7100 12470 7120 12530
rect 7180 12470 7200 12530
rect 7100 12430 7200 12470
rect 7100 12370 7120 12430
rect 7180 12370 7200 12430
rect 7100 12330 7200 12370
rect 7100 12270 7120 12330
rect 7180 12270 7200 12330
rect 7100 12250 7200 12270
rect 13750 12150 13900 22450
rect 9650 12130 13900 12150
rect 400 11900 6100 12100
rect 9650 12070 9670 12130
rect 9730 12070 9770 12130
rect 9830 12070 9870 12130
rect 9930 12070 9970 12130
rect 10030 12070 13900 12130
rect 9650 12050 13900 12070
rect 400 500 600 11900
rect 9650 11730 15300 11750
rect 9650 11670 9670 11730
rect 9730 11670 9770 11730
rect 9830 11670 9870 11730
rect 9930 11670 9970 11730
rect 10030 11670 15300 11730
rect 9650 11650 15300 11670
rect 9650 11480 13350 11500
rect 9650 11420 9670 11480
rect 9730 11420 9770 11480
rect 9830 11420 9870 11480
rect 9930 11420 9970 11480
rect 10030 11420 13350 11480
rect 9650 11400 13350 11420
rect 800 11150 6500 11200
rect 800 11050 850 11150
rect 950 11050 1050 11150
rect 1150 11050 1250 11150
rect 1350 11050 1450 11150
rect 1550 11050 6500 11150
rect 800 11000 6500 11050
rect 13200 100 13350 11400
rect 15150 100 15300 11650
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13249 0 13339 100
rect 15181 0 15271 100
use FAMILY  FAMILY_0 ~/dev/personal/chacha-silicon/tt09-analog-switch
timestamp 1730992266
transform 1 0 2000 0 1 1000
box 0 0 9990 7500
use SWTCH_UNIT2  SWTCH_UNIT2_0 design/SWTCH_UNIT2_SKY130NM
timestamp 1730931062
transform 1 0 7000 0 1 12300
box -1000 -1300 2600 -50
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 100 500 300 22076 1 FreeSans 1 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 1 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
