magic
tech sky130A
magscale 1 2
timestamp 1730924699
<< locali >>
rect -2020 940 -1060 1040
rect -1660 880 -1400 940
rect -1840 460 -1740 640
rect -1520 460 -1420 640
rect -1940 -500 -1840 -300
rect -1640 -500 -1540 -300
rect -1520 -500 -1420 -300
rect -1220 -500 -1120 -300
rect -1660 -920 -1400 -860
rect -2020 -1020 -1060 -920
<< metal1 >>
rect -2020 740 -1640 840
rect -1580 740 -1320 840
rect -2020 220 -1920 740
rect -1580 600 -1480 740
rect -1640 500 -1480 600
rect -1320 500 -1060 600
rect -1580 380 -1480 500
rect -1740 220 -1640 380
rect -2020 120 -1640 220
rect -2020 -720 -1920 120
rect -1740 -40 -1640 120
rect -1580 280 -1320 380
rect -1580 60 -1480 280
rect -1580 -40 -1220 60
rect -1720 -360 -1700 -340
rect -1720 -440 -1700 -420
rect -1580 -360 -1480 -40
rect -1580 -420 -1560 -360
rect -1500 -420 -1480 -360
rect -1580 -720 -1480 -420
rect -1360 -360 -1280 -340
rect -1360 -420 -1340 -360
rect -1360 -440 -1280 -420
rect -1160 -360 -1060 500
rect -1160 -420 -1140 -360
rect -1080 -420 -1060 -360
rect -1160 -440 -1060 -420
rect -2020 -820 -1740 -720
rect -1580 -820 -1320 -720
<< via1 >>
rect -1760 -420 -1700 -360
rect -1560 -420 -1500 -360
rect -1340 -420 -1280 -360
rect -1140 -420 -1080 -360
<< metal2 >>
rect -1780 -360 -1480 -340
rect -1780 -420 -1760 -360
rect -1700 -420 -1560 -360
rect -1500 -420 -1480 -360
rect -1780 -440 -1480 -420
rect -1360 -360 -1060 -340
rect -1360 -420 -1340 -360
rect -1280 -420 -1140 -360
rect -1080 -420 -1060 -360
rect -1360 -440 -1060 -420
use sky130_fd_pr__nfet_01v8_NRQ53D  sky130_fd_pr__nfet_01v8_NRQ53D_0
timestamp 1730922800
transform 1 0 -1689 0 1 560
box -211 -360 211 360
use sky130_fd_pr__nfet_01v8_NRQ53D  sky130_fd_pr__nfet_01v8_NRQ53D_2
timestamp 1730922800
transform 1 0 -1373 0 1 560
box -211 -360 211 360
use sky130_fd_pr__pfet_01v8_XW3LHL  sky130_fd_pr__pfet_01v8_XW3LHL_0
timestamp 1730922800
transform 1 0 -1317 0 1 -381
box -263 -519 263 519
use sky130_fd_pr__pfet_01v8_XW3LHL  sky130_fd_pr__pfet_01v8_XW3LHL_1
timestamp 1730922800
transform 1 0 -1737 0 1 -381
box -263 -519 263 519
<< labels >>
rlabel locali -2020 -1020 -1920 -920 1 VPWR
port 1 n
rlabel locali -2020 940 -1920 1040 1 VGND
port 2 n
rlabel metal1 -2020 120 -1920 220 1 IN
port 3 n
rlabel metal1 -1160 120 -1060 220 1 Q_P
port 4 n
rlabel metal1 -1580 120 -1480 220 1 Q_N
port 5 n
<< end >>
