magic
tech sky130A
timestamp 1730992266
<< locali >>
rect 2250 7490 3300 7500
rect 2250 7480 3300 7490
rect 2250 7470 3300 7480
rect 2250 7460 3300 7470
rect 2250 7450 3300 7460
rect 2200 7440 3300 7450
rect 2200 7430 3300 7440
rect 2200 7420 3300 7430
rect 2200 7410 3300 7420
rect 2200 7400 3300 7410
rect 2150 7390 3300 7400
rect 2150 7380 3300 7390
rect 2150 7370 3300 7380
rect 2150 7360 3300 7370
rect 2150 7350 3300 7360
rect 2100 7340 3300 7350
rect 2100 7330 3300 7340
rect 2100 7320 3300 7330
rect 2100 7310 3300 7320
rect 2100 7300 3300 7310
rect 2100 7290 2500 7300
rect 2550 7290 3300 7300
rect 2100 7280 2500 7290
rect 2550 7280 3300 7290
rect 2100 7270 2500 7280
rect 2550 7270 3300 7280
rect 2100 7260 2500 7270
rect 2550 7260 3300 7270
rect 2100 7250 2500 7260
rect 2550 7250 3300 7260
rect 2050 7240 2400 7250
rect 2450 7240 2500 7250
rect 2550 7240 3300 7250
rect 2050 7230 2400 7240
rect 2450 7230 2500 7240
rect 2550 7230 3300 7240
rect 2050 7220 2400 7230
rect 2450 7220 2500 7230
rect 2550 7220 3300 7230
rect 2050 7210 2400 7220
rect 2450 7210 2500 7220
rect 2550 7210 3300 7220
rect 2050 7200 2400 7210
rect 2450 7200 2500 7210
rect 2550 7200 3300 7210
rect 2050 7190 2100 7200
rect 2300 7190 3300 7200
rect 2050 7180 2100 7190
rect 2300 7180 3300 7190
rect 2050 7170 2100 7180
rect 2300 7170 3300 7180
rect 2050 7160 2100 7170
rect 2300 7160 3300 7170
rect 2050 7150 2100 7160
rect 2300 7150 3300 7160
rect 2250 7140 3300 7150
rect 2250 7130 3300 7140
rect 2250 7120 3300 7130
rect 2250 7110 3300 7120
rect 2250 7100 3300 7110
rect 2150 7090 2250 7100
rect 2400 7090 3400 7100
rect 9850 7090 9950 7100
rect 2150 7080 2250 7090
rect 2400 7080 3400 7090
rect 9850 7080 9950 7090
rect 2150 7070 2250 7080
rect 2400 7070 3400 7080
rect 9850 7070 9950 7080
rect 2150 7060 2250 7070
rect 2400 7060 3400 7070
rect 9850 7060 9950 7070
rect 2150 7050 2250 7060
rect 2400 7050 3400 7060
rect 9850 7050 9950 7060
rect 2100 7040 2200 7050
rect 3250 7040 3450 7050
rect 9850 7040 9900 7050
rect 2100 7030 2200 7040
rect 3250 7030 3450 7040
rect 9850 7030 9900 7040
rect 2100 7020 2200 7030
rect 3250 7020 3450 7030
rect 9850 7020 9900 7030
rect 2100 7010 2200 7020
rect 3250 7010 3450 7020
rect 9850 7010 9900 7020
rect 2100 7000 2200 7010
rect 3250 7000 3450 7010
rect 9850 7000 9900 7010
rect 2050 6990 2150 7000
rect 3400 6990 3500 7000
rect 9900 6990 9990 7000
rect 2050 6980 2150 6990
rect 3400 6980 3500 6990
rect 9900 6980 9990 6990
rect 2050 6970 2150 6980
rect 3400 6970 3500 6980
rect 9900 6970 9990 6980
rect 2050 6960 2150 6970
rect 3400 6960 3500 6970
rect 9900 6960 9990 6970
rect 2050 6950 2150 6960
rect 3400 6950 3500 6960
rect 9900 6950 9990 6960
rect 2000 6940 2200 6950
rect 9850 6940 9990 6950
rect 2000 6930 2200 6940
rect 9850 6930 9990 6940
rect 2000 6920 2200 6930
rect 9850 6920 9990 6930
rect 2000 6910 2200 6920
rect 9850 6910 9990 6920
rect 2000 6900 2200 6910
rect 9850 6900 9990 6910
rect 1950 6890 2250 6900
rect 9850 6890 9990 6900
rect 1950 6880 2250 6890
rect 9850 6880 9990 6890
rect 1950 6870 2250 6880
rect 9850 6870 9990 6880
rect 1950 6860 2250 6870
rect 9850 6860 9990 6870
rect 1950 6850 2250 6860
rect 9850 6850 9990 6860
rect 2000 6840 2300 6850
rect 2000 6830 2300 6840
rect 2000 6820 2300 6830
rect 2000 6810 2300 6820
rect 2000 6800 2300 6810
rect 2050 6790 2250 6800
rect 9850 6790 9900 6800
rect 2050 6780 2250 6790
rect 9850 6780 9900 6790
rect 2050 6770 2250 6780
rect 9850 6770 9900 6780
rect 2050 6760 2250 6770
rect 9850 6760 9900 6770
rect 2050 6750 2250 6760
rect 9850 6750 9900 6760
rect 2000 6740 2200 6750
rect 2600 6740 2800 6750
rect 9850 6740 9950 6750
rect 2000 6730 2200 6740
rect 2600 6730 2800 6740
rect 9850 6730 9950 6740
rect 2000 6720 2200 6730
rect 2600 6720 2800 6730
rect 9850 6720 9950 6730
rect 2000 6710 2200 6720
rect 2600 6710 2800 6720
rect 9850 6710 9950 6720
rect 2000 6700 2200 6710
rect 2600 6700 2800 6710
rect 9850 6700 9950 6710
rect 1950 6690 2200 6700
rect 2650 6690 3200 6700
rect 1950 6680 2200 6690
rect 2650 6680 3200 6690
rect 1950 6670 2200 6680
rect 2650 6670 3200 6680
rect 1950 6660 2200 6670
rect 2650 6660 3200 6670
rect 1950 6650 2200 6660
rect 2650 6650 3200 6660
rect 1900 6640 2100 6650
rect 2650 6640 3450 6650
rect 1900 6630 2100 6640
rect 2650 6630 3450 6640
rect 1900 6620 2100 6630
rect 2650 6620 3450 6630
rect 1900 6610 2100 6620
rect 2650 6610 3450 6620
rect 1900 6600 2100 6610
rect 2650 6600 3450 6610
rect 1850 6590 2000 6600
rect 2700 6590 3600 6600
rect 1850 6580 2000 6590
rect 2700 6580 3600 6590
rect 1850 6570 2000 6580
rect 2700 6570 3600 6580
rect 1850 6560 2000 6570
rect 2700 6560 3600 6570
rect 1850 6550 2000 6560
rect 2700 6550 3600 6560
rect 1900 6540 2000 6550
rect 2650 6540 3700 6550
rect 1900 6530 2000 6540
rect 2650 6530 3700 6540
rect 1900 6520 2000 6530
rect 2650 6520 3700 6530
rect 1900 6510 2000 6520
rect 2650 6510 3700 6520
rect 1900 6500 2000 6510
rect 2650 6500 3700 6510
rect 1450 6490 1550 6500
rect 2600 6490 3800 6500
rect 1450 6480 1550 6490
rect 2600 6480 3800 6490
rect 1450 6470 1550 6480
rect 2600 6470 3800 6480
rect 1450 6460 1550 6470
rect 2600 6460 3800 6470
rect 1450 6450 1550 6460
rect 2600 6450 3800 6460
rect 1500 6440 1550 6450
rect 2600 6440 3900 6450
rect 9850 6440 9900 6450
rect 1500 6430 1550 6440
rect 2600 6430 3900 6440
rect 9850 6430 9900 6440
rect 1500 6420 1550 6430
rect 2600 6420 3900 6430
rect 9850 6420 9900 6430
rect 1500 6410 1550 6420
rect 2600 6410 3900 6420
rect 9850 6410 9900 6420
rect 1500 6400 1550 6410
rect 2600 6400 3900 6410
rect 9850 6400 9900 6410
rect 1500 6390 1550 6400
rect 2500 6390 4000 6400
rect 9850 6390 9900 6400
rect 1500 6380 1550 6390
rect 2500 6380 4000 6390
rect 9850 6380 9900 6390
rect 1500 6370 1550 6380
rect 2500 6370 4000 6380
rect 9850 6370 9900 6380
rect 1500 6360 1550 6370
rect 2500 6360 4000 6370
rect 9850 6360 9900 6370
rect 1500 6350 1550 6360
rect 2500 6350 4000 6360
rect 9850 6350 9900 6360
rect 1500 6340 1550 6350
rect 2500 6340 4050 6350
rect 1500 6330 1550 6340
rect 2500 6330 4050 6340
rect 1500 6320 1550 6330
rect 2500 6320 4050 6330
rect 1500 6310 1550 6320
rect 2500 6310 4050 6320
rect 1500 6300 1550 6310
rect 2500 6300 4050 6310
rect 1450 6290 1550 6300
rect 2500 6290 4100 6300
rect 9700 6290 9800 6300
rect 1450 6280 1550 6290
rect 2500 6280 4100 6290
rect 9700 6280 9800 6290
rect 1450 6270 1550 6280
rect 2500 6270 4100 6280
rect 9700 6270 9800 6280
rect 1450 6260 1550 6270
rect 2500 6260 4100 6270
rect 9700 6260 9800 6270
rect 1450 6250 1550 6260
rect 2500 6250 4100 6260
rect 9700 6250 9800 6260
rect 1450 6240 1550 6250
rect 2500 6240 4150 6250
rect 9700 6240 9750 6250
rect 1450 6230 1550 6240
rect 2500 6230 4150 6240
rect 9700 6230 9750 6240
rect 1450 6220 1550 6230
rect 2500 6220 4150 6230
rect 9700 6220 9750 6230
rect 1450 6210 1550 6220
rect 2500 6210 4150 6220
rect 9700 6210 9750 6220
rect 1450 6200 1550 6210
rect 2500 6200 4150 6210
rect 9700 6200 9750 6210
rect 1450 6190 1550 6200
rect 2450 6190 4200 6200
rect 9500 6190 9550 6200
rect 1450 6180 1550 6190
rect 2450 6180 4200 6190
rect 9500 6180 9550 6190
rect 1450 6170 1550 6180
rect 2450 6170 4200 6180
rect 9500 6170 9550 6180
rect 1450 6160 1550 6170
rect 2450 6160 4200 6170
rect 9500 6160 9550 6170
rect 1450 6150 1550 6160
rect 2450 6150 4200 6160
rect 9500 6150 9550 6160
rect 1450 6140 1600 6150
rect 2500 6140 3850 6150
rect 4000 6140 4250 6150
rect 9500 6140 9600 6150
rect 9700 6140 9800 6150
rect 1450 6130 1600 6140
rect 2500 6130 3850 6140
rect 4000 6130 4250 6140
rect 9500 6130 9600 6140
rect 9700 6130 9800 6140
rect 1450 6120 1600 6130
rect 2500 6120 3850 6130
rect 4000 6120 4250 6130
rect 9500 6120 9600 6130
rect 9700 6120 9800 6130
rect 1450 6110 1600 6120
rect 2500 6110 3850 6120
rect 4000 6110 4250 6120
rect 9500 6110 9600 6120
rect 9700 6110 9800 6120
rect 1450 6100 1600 6110
rect 2500 6100 3850 6110
rect 4000 6100 4250 6110
rect 9500 6100 9600 6110
rect 9700 6100 9800 6110
rect 1450 6090 1550 6100
rect 2500 6090 3750 6100
rect 4050 6090 4250 6100
rect 5300 6090 5350 6100
rect 9550 6090 9600 6100
rect 9750 6090 9800 6100
rect 1450 6080 1550 6090
rect 2500 6080 3750 6090
rect 4050 6080 4250 6090
rect 5300 6080 5350 6090
rect 9550 6080 9600 6090
rect 9750 6080 9800 6090
rect 1450 6070 1550 6080
rect 2500 6070 3750 6080
rect 4050 6070 4250 6080
rect 5300 6070 5350 6080
rect 9550 6070 9600 6080
rect 9750 6070 9800 6080
rect 1450 6060 1550 6070
rect 2500 6060 3750 6070
rect 4050 6060 4250 6070
rect 5300 6060 5350 6070
rect 9550 6060 9600 6070
rect 9750 6060 9800 6070
rect 1450 6050 1550 6060
rect 2500 6050 3750 6060
rect 4050 6050 4250 6060
rect 5300 6050 5350 6060
rect 9550 6050 9600 6060
rect 9750 6050 9800 6060
rect 1350 6040 1600 6050
rect 2550 6040 3150 6050
rect 3300 6040 3750 6050
rect 4100 6040 4300 6050
rect 9550 6040 9650 6050
rect 9750 6040 9800 6050
rect 1350 6030 1600 6040
rect 2550 6030 3150 6040
rect 3300 6030 3750 6040
rect 4100 6030 4300 6040
rect 9550 6030 9650 6040
rect 9750 6030 9800 6040
rect 1350 6020 1600 6030
rect 2550 6020 3150 6030
rect 3300 6020 3750 6030
rect 4100 6020 4300 6030
rect 9550 6020 9650 6030
rect 9750 6020 9800 6030
rect 1350 6010 1600 6020
rect 2550 6010 3150 6020
rect 3300 6010 3750 6020
rect 4100 6010 4300 6020
rect 9550 6010 9650 6020
rect 9750 6010 9800 6020
rect 1350 6000 1600 6010
rect 2550 6000 3150 6010
rect 3300 6000 3750 6010
rect 4100 6000 4300 6010
rect 9550 6000 9650 6010
rect 9750 6000 9800 6010
rect 1350 5990 1600 6000
rect 2600 5990 3100 6000
rect 3300 5990 3700 6000
rect 4200 5990 4300 6000
rect 5250 5990 5300 6000
rect 9550 5990 9650 6000
rect 9750 5990 9850 6000
rect 1350 5980 1600 5990
rect 2600 5980 3100 5990
rect 3300 5980 3700 5990
rect 4200 5980 4300 5990
rect 5250 5980 5300 5990
rect 9550 5980 9650 5990
rect 9750 5980 9850 5990
rect 1350 5970 1600 5980
rect 2600 5970 3100 5980
rect 3300 5970 3700 5980
rect 4200 5970 4300 5980
rect 5250 5970 5300 5980
rect 9550 5970 9650 5980
rect 9750 5970 9850 5980
rect 1350 5960 1600 5970
rect 2600 5960 3100 5970
rect 3300 5960 3700 5970
rect 4200 5960 4300 5970
rect 5250 5960 5300 5970
rect 9550 5960 9650 5970
rect 9750 5960 9850 5970
rect 1350 5950 1600 5960
rect 2600 5950 3100 5960
rect 3300 5950 3700 5960
rect 4200 5950 4300 5960
rect 5250 5950 5300 5960
rect 9550 5950 9650 5960
rect 9750 5950 9850 5960
rect 1200 5940 1650 5950
rect 2650 5940 3050 5950
rect 3300 5940 3700 5950
rect 5200 5940 5300 5950
rect 9550 5940 9700 5950
rect 9750 5940 9850 5950
rect 1200 5930 1650 5940
rect 2650 5930 3050 5940
rect 3300 5930 3700 5940
rect 5200 5930 5300 5940
rect 9550 5930 9700 5940
rect 9750 5930 9850 5940
rect 1200 5920 1650 5930
rect 2650 5920 3050 5930
rect 3300 5920 3700 5930
rect 5200 5920 5300 5930
rect 9550 5920 9700 5930
rect 9750 5920 9850 5930
rect 1200 5910 1650 5920
rect 2650 5910 3050 5920
rect 3300 5910 3700 5920
rect 5200 5910 5300 5920
rect 9550 5910 9700 5920
rect 9750 5910 9850 5920
rect 1200 5900 1650 5910
rect 2650 5900 3050 5910
rect 3300 5900 3700 5910
rect 5200 5900 5300 5910
rect 9550 5900 9700 5910
rect 9750 5900 9850 5910
rect 1050 5890 1700 5900
rect 2700 5890 2900 5900
rect 3300 5890 3700 5900
rect 5200 5890 5300 5900
rect 9450 5890 9850 5900
rect 1050 5880 1700 5890
rect 2700 5880 2900 5890
rect 3300 5880 3700 5890
rect 5200 5880 5300 5890
rect 9450 5880 9850 5890
rect 1050 5870 1700 5880
rect 2700 5870 2900 5880
rect 3300 5870 3700 5880
rect 5200 5870 5300 5880
rect 9450 5870 9850 5880
rect 1050 5860 1700 5870
rect 2700 5860 2900 5870
rect 3300 5860 3700 5870
rect 5200 5860 5300 5870
rect 9450 5860 9850 5870
rect 1050 5850 1700 5860
rect 2700 5850 2900 5860
rect 3300 5850 3700 5860
rect 5200 5850 5300 5860
rect 9450 5850 9850 5860
rect 1000 5840 1800 5850
rect 3300 5840 3700 5850
rect 5150 5840 5250 5850
rect 9350 5840 9900 5850
rect 1000 5830 1800 5840
rect 3300 5830 3700 5840
rect 5150 5830 5250 5840
rect 9350 5830 9900 5840
rect 1000 5820 1800 5830
rect 3300 5820 3700 5830
rect 5150 5820 5250 5830
rect 9350 5820 9900 5830
rect 1000 5810 1800 5820
rect 3300 5810 3700 5820
rect 5150 5810 5250 5820
rect 9350 5810 9900 5820
rect 1000 5800 1800 5810
rect 3300 5800 3700 5810
rect 5150 5800 5250 5810
rect 9350 5800 9900 5810
rect 950 5790 1800 5800
rect 3300 5790 3700 5800
rect 5150 5790 5250 5800
rect 9250 5790 9900 5800
rect 950 5780 1800 5790
rect 3300 5780 3700 5790
rect 5150 5780 5250 5790
rect 9250 5780 9900 5790
rect 950 5770 1800 5780
rect 3300 5770 3700 5780
rect 5150 5770 5250 5780
rect 9250 5770 9900 5780
rect 950 5760 1800 5770
rect 3300 5760 3700 5770
rect 5150 5760 5250 5770
rect 9250 5760 9900 5770
rect 950 5750 1800 5760
rect 3300 5750 3700 5760
rect 5150 5750 5250 5760
rect 9250 5750 9900 5760
rect 900 5740 1100 5750
rect 1250 5740 1800 5750
rect 3350 5740 3700 5750
rect 5150 5740 5250 5750
rect 9050 5740 9900 5750
rect 900 5730 1100 5740
rect 1250 5730 1800 5740
rect 3350 5730 3700 5740
rect 5150 5730 5250 5740
rect 9050 5730 9900 5740
rect 900 5720 1100 5730
rect 1250 5720 1800 5730
rect 3350 5720 3700 5730
rect 5150 5720 5250 5730
rect 9050 5720 9900 5730
rect 900 5710 1100 5720
rect 1250 5710 1800 5720
rect 3350 5710 3700 5720
rect 5150 5710 5250 5720
rect 9050 5710 9900 5720
rect 900 5700 1100 5710
rect 1250 5700 1800 5710
rect 3350 5700 3700 5710
rect 5150 5700 5250 5710
rect 9050 5700 9900 5710
rect 850 5690 1050 5700
rect 1250 5690 1850 5700
rect 3350 5690 3650 5700
rect 5150 5690 5250 5700
rect 8800 5690 8950 5700
rect 9000 5690 9950 5700
rect 850 5680 1050 5690
rect 1250 5680 1850 5690
rect 3350 5680 3650 5690
rect 5150 5680 5250 5690
rect 8800 5680 8950 5690
rect 9000 5680 9950 5690
rect 850 5670 1050 5680
rect 1250 5670 1850 5680
rect 3350 5670 3650 5680
rect 5150 5670 5250 5680
rect 8800 5670 8950 5680
rect 9000 5670 9950 5680
rect 850 5660 1050 5670
rect 1250 5660 1850 5670
rect 3350 5660 3650 5670
rect 5150 5660 5250 5670
rect 8800 5660 8950 5670
rect 9000 5660 9950 5670
rect 850 5650 1050 5660
rect 1250 5650 1850 5660
rect 3350 5650 3650 5660
rect 5150 5650 5250 5660
rect 8800 5650 8950 5660
rect 9000 5650 9950 5660
rect 850 5640 1850 5650
rect 3300 5640 3400 5650
rect 3450 5640 3650 5650
rect 5150 5640 5250 5650
rect 8550 5640 8900 5650
rect 9100 5640 9950 5650
rect 850 5630 1850 5640
rect 3300 5630 3400 5640
rect 3450 5630 3650 5640
rect 5150 5630 5250 5640
rect 8550 5630 8900 5640
rect 9100 5630 9950 5640
rect 850 5620 1850 5630
rect 3300 5620 3400 5630
rect 3450 5620 3650 5630
rect 5150 5620 5250 5630
rect 8550 5620 8900 5630
rect 9100 5620 9950 5630
rect 850 5610 1850 5620
rect 3300 5610 3400 5620
rect 3450 5610 3650 5620
rect 5150 5610 5250 5620
rect 8550 5610 8900 5620
rect 9100 5610 9950 5620
rect 850 5600 1850 5610
rect 3300 5600 3400 5610
rect 3450 5600 3650 5610
rect 5150 5600 5250 5610
rect 8550 5600 8900 5610
rect 9100 5600 9950 5610
rect 750 5590 1850 5600
rect 3350 5590 3400 5600
rect 3500 5590 3600 5600
rect 5150 5590 5200 5600
rect 8500 5590 8750 5600
rect 9150 5590 9950 5600
rect 750 5580 1850 5590
rect 3350 5580 3400 5590
rect 3500 5580 3600 5590
rect 5150 5580 5200 5590
rect 8500 5580 8750 5590
rect 9150 5580 9950 5590
rect 750 5570 1850 5580
rect 3350 5570 3400 5580
rect 3500 5570 3600 5580
rect 5150 5570 5200 5580
rect 8500 5570 8750 5580
rect 9150 5570 9950 5580
rect 750 5560 1850 5570
rect 3350 5560 3400 5570
rect 3500 5560 3600 5570
rect 5150 5560 5200 5570
rect 8500 5560 8750 5570
rect 9150 5560 9950 5570
rect 750 5550 1850 5560
rect 3350 5550 3400 5560
rect 3500 5550 3600 5560
rect 5150 5550 5200 5560
rect 8500 5550 8750 5560
rect 9150 5550 9950 5560
rect 700 5540 900 5550
rect 1000 5540 1850 5550
rect 3350 5540 3450 5550
rect 3550 5540 3600 5550
rect 5150 5540 5200 5550
rect 8350 5540 8600 5550
rect 9150 5540 9990 5550
rect 700 5530 900 5540
rect 1000 5530 1850 5540
rect 3350 5530 3450 5540
rect 3550 5530 3600 5540
rect 5150 5530 5200 5540
rect 8350 5530 8600 5540
rect 9150 5530 9990 5540
rect 700 5520 900 5530
rect 1000 5520 1850 5530
rect 3350 5520 3450 5530
rect 3550 5520 3600 5530
rect 5150 5520 5200 5530
rect 8350 5520 8600 5530
rect 9150 5520 9990 5530
rect 700 5510 900 5520
rect 1000 5510 1850 5520
rect 3350 5510 3450 5520
rect 3550 5510 3600 5520
rect 5150 5510 5200 5520
rect 8350 5510 8600 5520
rect 9150 5510 9990 5520
rect 700 5500 900 5510
rect 1000 5500 1850 5510
rect 3350 5500 3450 5510
rect 3550 5500 3600 5510
rect 5150 5500 5200 5510
rect 8350 5500 8600 5510
rect 9150 5500 9990 5510
rect 650 5490 900 5500
rect 1000 5490 1900 5500
rect 3350 5490 3550 5500
rect 5150 5490 5200 5500
rect 6250 5490 6350 5500
rect 8200 5490 8400 5500
rect 9150 5490 9990 5500
rect 650 5480 900 5490
rect 1000 5480 1900 5490
rect 3350 5480 3550 5490
rect 5150 5480 5200 5490
rect 6250 5480 6350 5490
rect 8200 5480 8400 5490
rect 9150 5480 9990 5490
rect 650 5470 900 5480
rect 1000 5470 1900 5480
rect 3350 5470 3550 5480
rect 5150 5470 5200 5480
rect 6250 5470 6350 5480
rect 8200 5470 8400 5480
rect 9150 5470 9990 5480
rect 650 5460 900 5470
rect 1000 5460 1900 5470
rect 3350 5460 3550 5470
rect 5150 5460 5200 5470
rect 6250 5460 6350 5470
rect 8200 5460 8400 5470
rect 9150 5460 9990 5470
rect 650 5450 900 5460
rect 1000 5450 1900 5460
rect 3350 5450 3550 5460
rect 5150 5450 5200 5460
rect 6250 5450 6350 5460
rect 8200 5450 8400 5460
rect 9150 5450 9990 5460
rect 650 5440 1900 5450
rect 2450 5440 2550 5450
rect 3300 5440 3550 5450
rect 5150 5440 5200 5450
rect 5750 5440 5800 5450
rect 6250 5440 6400 5450
rect 8150 5440 8250 5450
rect 9150 5440 9400 5450
rect 9650 5440 9990 5450
rect 650 5430 1900 5440
rect 2450 5430 2550 5440
rect 3300 5430 3550 5440
rect 5150 5430 5200 5440
rect 5750 5430 5800 5440
rect 6250 5430 6400 5440
rect 8150 5430 8250 5440
rect 9150 5430 9400 5440
rect 9650 5430 9990 5440
rect 650 5420 1900 5430
rect 2450 5420 2550 5430
rect 3300 5420 3550 5430
rect 5150 5420 5200 5430
rect 5750 5420 5800 5430
rect 6250 5420 6400 5430
rect 8150 5420 8250 5430
rect 9150 5420 9400 5430
rect 9650 5420 9990 5430
rect 650 5410 1900 5420
rect 2450 5410 2550 5420
rect 3300 5410 3550 5420
rect 5150 5410 5200 5420
rect 5750 5410 5800 5420
rect 6250 5410 6400 5420
rect 8150 5410 8250 5420
rect 9150 5410 9400 5420
rect 9650 5410 9990 5420
rect 650 5400 1900 5410
rect 2450 5400 2550 5410
rect 3300 5400 3550 5410
rect 5150 5400 5200 5410
rect 5750 5400 5800 5410
rect 6250 5400 6400 5410
rect 8150 5400 8250 5410
rect 9150 5400 9400 5410
rect 9650 5400 9990 5410
rect 600 5390 1900 5400
rect 2500 5390 2550 5400
rect 3200 5390 3500 5400
rect 5150 5390 5200 5400
rect 5750 5390 5800 5400
rect 6250 5390 6550 5400
rect 9100 5390 9250 5400
rect 9650 5390 9990 5400
rect 600 5380 1900 5390
rect 2500 5380 2550 5390
rect 3200 5380 3500 5390
rect 5150 5380 5200 5390
rect 5750 5380 5800 5390
rect 6250 5380 6550 5390
rect 9100 5380 9250 5390
rect 9650 5380 9990 5390
rect 600 5370 1900 5380
rect 2500 5370 2550 5380
rect 3200 5370 3500 5380
rect 5150 5370 5200 5380
rect 5750 5370 5800 5380
rect 6250 5370 6550 5380
rect 9100 5370 9250 5380
rect 9650 5370 9990 5380
rect 600 5360 1900 5370
rect 2500 5360 2550 5370
rect 3200 5360 3500 5370
rect 5150 5360 5200 5370
rect 5750 5360 5800 5370
rect 6250 5360 6550 5370
rect 9100 5360 9250 5370
rect 9650 5360 9990 5370
rect 600 5350 1900 5360
rect 2500 5350 2550 5360
rect 3200 5350 3500 5360
rect 5150 5350 5200 5360
rect 5750 5350 5800 5360
rect 6250 5350 6550 5360
rect 9100 5350 9250 5360
rect 9650 5350 9990 5360
rect 600 5340 1900 5350
rect 3050 5340 3500 5350
rect 7750 5340 7800 5350
rect 8950 5340 9000 5350
rect 9650 5340 9900 5350
rect 600 5330 1900 5340
rect 3050 5330 3500 5340
rect 7750 5330 7800 5340
rect 8950 5330 9000 5340
rect 9650 5330 9900 5340
rect 600 5320 1900 5330
rect 3050 5320 3500 5330
rect 7750 5320 7800 5330
rect 8950 5320 9000 5330
rect 9650 5320 9900 5330
rect 600 5310 1900 5320
rect 3050 5310 3500 5320
rect 7750 5310 7800 5320
rect 8950 5310 9000 5320
rect 9650 5310 9900 5320
rect 600 5300 1900 5310
rect 3050 5300 3500 5310
rect 7750 5300 7800 5310
rect 8950 5300 9000 5310
rect 9650 5300 9900 5310
rect 650 5290 1950 5300
rect 3000 5290 3450 5300
rect 7700 5290 7850 5300
rect 8750 5290 8800 5300
rect 9650 5290 9700 5300
rect 650 5280 1950 5290
rect 3000 5280 3450 5290
rect 7700 5280 7850 5290
rect 8750 5280 8800 5290
rect 9650 5280 9700 5290
rect 650 5270 1950 5280
rect 3000 5270 3450 5280
rect 7700 5270 7850 5280
rect 8750 5270 8800 5280
rect 9650 5270 9700 5280
rect 650 5260 1950 5270
rect 3000 5260 3450 5270
rect 7700 5260 7850 5270
rect 8750 5260 8800 5270
rect 9650 5260 9700 5270
rect 650 5250 1950 5260
rect 3000 5250 3450 5260
rect 7700 5250 7850 5260
rect 8750 5250 8800 5260
rect 9650 5250 9700 5260
rect 700 5240 1950 5250
rect 3000 5240 3450 5250
rect 7450 5240 7550 5250
rect 7650 5240 7850 5250
rect 700 5230 1950 5240
rect 3000 5230 3450 5240
rect 7450 5230 7550 5240
rect 7650 5230 7850 5240
rect 700 5220 1950 5230
rect 3000 5220 3450 5230
rect 7450 5220 7550 5230
rect 7650 5220 7850 5230
rect 700 5210 1950 5220
rect 3000 5210 3450 5220
rect 7450 5210 7550 5220
rect 7650 5210 7850 5220
rect 700 5200 1950 5210
rect 3000 5200 3450 5210
rect 7450 5200 7550 5210
rect 7650 5200 7850 5210
rect 750 5190 1800 5200
rect 1850 5190 1950 5200
rect 3050 5190 3400 5200
rect 7450 5190 7550 5200
rect 7650 5190 7850 5200
rect 750 5180 1800 5190
rect 1850 5180 1950 5190
rect 3050 5180 3400 5190
rect 7450 5180 7550 5190
rect 7650 5180 7850 5190
rect 750 5170 1800 5180
rect 1850 5170 1950 5180
rect 3050 5170 3400 5180
rect 7450 5170 7550 5180
rect 7650 5170 7850 5180
rect 750 5160 1800 5170
rect 1850 5160 1950 5170
rect 3050 5160 3400 5170
rect 7450 5160 7550 5170
rect 7650 5160 7850 5170
rect 750 5150 1800 5160
rect 1850 5150 1950 5160
rect 3050 5150 3400 5160
rect 7450 5150 7550 5160
rect 7650 5150 7850 5160
rect 750 5140 1800 5150
rect 1900 5140 1950 5150
rect 3050 5140 3400 5150
rect 7450 5140 7850 5150
rect 8550 5140 8600 5150
rect 750 5130 1800 5140
rect 1900 5130 1950 5140
rect 3050 5130 3400 5140
rect 7450 5130 7850 5140
rect 8550 5130 8600 5140
rect 750 5120 1800 5130
rect 1900 5120 1950 5130
rect 3050 5120 3400 5130
rect 7450 5120 7850 5130
rect 8550 5120 8600 5130
rect 750 5110 1800 5120
rect 1900 5110 1950 5120
rect 3050 5110 3400 5120
rect 7450 5110 7850 5120
rect 8550 5110 8600 5120
rect 750 5100 1800 5110
rect 1900 5100 1950 5110
rect 3050 5100 3400 5110
rect 7450 5100 7850 5110
rect 8550 5100 8600 5110
rect 750 5090 1750 5100
rect 1900 5090 1950 5100
rect 3050 5090 3350 5100
rect 7450 5090 7850 5100
rect 8550 5090 8600 5100
rect 9900 5090 9990 5100
rect 750 5080 1750 5090
rect 1900 5080 1950 5090
rect 3050 5080 3350 5090
rect 7450 5080 7850 5090
rect 8550 5080 8600 5090
rect 9900 5080 9990 5090
rect 750 5070 1750 5080
rect 1900 5070 1950 5080
rect 3050 5070 3350 5080
rect 7450 5070 7850 5080
rect 8550 5070 8600 5080
rect 9900 5070 9990 5080
rect 750 5060 1750 5070
rect 1900 5060 1950 5070
rect 3050 5060 3350 5070
rect 7450 5060 7850 5070
rect 8550 5060 8600 5070
rect 9900 5060 9990 5070
rect 750 5050 1750 5060
rect 1900 5050 1950 5060
rect 3050 5050 3350 5060
rect 7450 5050 7850 5060
rect 8550 5050 8600 5060
rect 9900 5050 9990 5060
rect 600 5040 1750 5050
rect 1900 5040 2000 5050
rect 3050 5040 3350 5050
rect 7450 5040 7850 5050
rect 8600 5040 8650 5050
rect 9700 5040 9990 5050
rect 600 5030 1750 5040
rect 1900 5030 2000 5040
rect 3050 5030 3350 5040
rect 7450 5030 7850 5040
rect 8600 5030 8650 5040
rect 9700 5030 9990 5040
rect 600 5020 1750 5030
rect 1900 5020 2000 5030
rect 3050 5020 3350 5030
rect 7450 5020 7850 5030
rect 8600 5020 8650 5030
rect 9700 5020 9990 5030
rect 600 5010 1750 5020
rect 1900 5010 2000 5020
rect 3050 5010 3350 5020
rect 7450 5010 7850 5020
rect 8600 5010 8650 5020
rect 9700 5010 9990 5020
rect 600 5000 1750 5010
rect 1900 5000 2000 5010
rect 3050 5000 3350 5010
rect 7450 5000 7850 5010
rect 8600 5000 8650 5010
rect 9700 5000 9990 5010
rect 550 4990 1800 5000
rect 1850 4990 2050 5000
rect 3000 4990 3300 5000
rect 7400 4990 7750 5000
rect 9750 4990 9990 5000
rect 550 4980 1800 4990
rect 1850 4980 2050 4990
rect 3000 4980 3300 4990
rect 7400 4980 7750 4990
rect 9750 4980 9990 4990
rect 550 4970 1800 4980
rect 1850 4970 2050 4980
rect 3000 4970 3300 4980
rect 7400 4970 7750 4980
rect 9750 4970 9990 4980
rect 550 4960 1800 4970
rect 1850 4960 2050 4970
rect 3000 4960 3300 4970
rect 7400 4960 7750 4970
rect 9750 4960 9990 4970
rect 550 4950 1800 4960
rect 1850 4950 2050 4960
rect 3000 4950 3300 4960
rect 7400 4950 7750 4960
rect 9750 4950 9990 4960
rect 700 4940 2100 4950
rect 2900 4940 3300 4950
rect 7400 4940 7650 4950
rect 9750 4940 9990 4950
rect 700 4930 2100 4940
rect 2900 4930 3300 4940
rect 7400 4930 7650 4940
rect 9750 4930 9990 4940
rect 700 4920 2100 4930
rect 2900 4920 3300 4930
rect 7400 4920 7650 4930
rect 9750 4920 9990 4930
rect 700 4910 2100 4920
rect 2900 4910 3300 4920
rect 7400 4910 7650 4920
rect 9750 4910 9990 4920
rect 700 4900 2100 4910
rect 2900 4900 3300 4910
rect 7400 4900 7650 4910
rect 9750 4900 9990 4910
rect 750 4890 1050 4900
rect 1100 4890 2150 4900
rect 2850 4890 3100 4900
rect 3200 4890 3250 4900
rect 4200 4890 4450 4900
rect 7400 4890 7650 4900
rect 9800 4890 9990 4900
rect 750 4880 1050 4890
rect 1100 4880 2150 4890
rect 2850 4880 3100 4890
rect 3200 4880 3250 4890
rect 4200 4880 4450 4890
rect 7400 4880 7650 4890
rect 9800 4880 9990 4890
rect 750 4870 1050 4880
rect 1100 4870 2150 4880
rect 2850 4870 3100 4880
rect 3200 4870 3250 4880
rect 4200 4870 4450 4880
rect 7400 4870 7650 4880
rect 9800 4870 9990 4880
rect 750 4860 1050 4870
rect 1100 4860 2150 4870
rect 2850 4860 3100 4870
rect 3200 4860 3250 4870
rect 4200 4860 4450 4870
rect 7400 4860 7650 4870
rect 9800 4860 9990 4870
rect 750 4850 1050 4860
rect 1100 4850 2150 4860
rect 2850 4850 3100 4860
rect 3200 4850 3250 4860
rect 4200 4850 4450 4860
rect 7400 4850 7650 4860
rect 9800 4850 9990 4860
rect 850 4840 1000 4850
rect 1100 4840 2300 4850
rect 2850 4840 3050 4850
rect 4050 4840 4850 4850
rect 7400 4840 7650 4850
rect 9800 4840 9990 4850
rect 850 4830 1000 4840
rect 1100 4830 2300 4840
rect 2850 4830 3050 4840
rect 4050 4830 4850 4840
rect 7400 4830 7650 4840
rect 9800 4830 9990 4840
rect 850 4820 1000 4830
rect 1100 4820 2300 4830
rect 2850 4820 3050 4830
rect 4050 4820 4850 4830
rect 7400 4820 7650 4830
rect 9800 4820 9990 4830
rect 850 4810 1000 4820
rect 1100 4810 2300 4820
rect 2850 4810 3050 4820
rect 4050 4810 4850 4820
rect 7400 4810 7650 4820
rect 9800 4810 9990 4820
rect 850 4800 1000 4810
rect 1100 4800 2300 4810
rect 2850 4800 3050 4810
rect 4050 4800 4850 4810
rect 7400 4800 7650 4810
rect 9800 4800 9990 4810
rect 400 4790 500 4800
rect 950 4790 1050 4800
rect 1150 4790 2350 4800
rect 3150 4790 3200 4800
rect 3650 4790 3800 4800
rect 3950 4790 4950 4800
rect 7400 4790 7650 4800
rect 9750 4790 9850 4800
rect 400 4780 500 4790
rect 950 4780 1050 4790
rect 1150 4780 2350 4790
rect 3150 4780 3200 4790
rect 3650 4780 3800 4790
rect 3950 4780 4950 4790
rect 7400 4780 7650 4790
rect 9750 4780 9850 4790
rect 400 4770 500 4780
rect 950 4770 1050 4780
rect 1150 4770 2350 4780
rect 3150 4770 3200 4780
rect 3650 4770 3800 4780
rect 3950 4770 4950 4780
rect 7400 4770 7650 4780
rect 9750 4770 9850 4780
rect 400 4760 500 4770
rect 950 4760 1050 4770
rect 1150 4760 2350 4770
rect 3150 4760 3200 4770
rect 3650 4760 3800 4770
rect 3950 4760 4950 4770
rect 7400 4760 7650 4770
rect 9750 4760 9850 4770
rect 400 4750 500 4760
rect 950 4750 1050 4760
rect 1150 4750 2350 4760
rect 3150 4750 3200 4760
rect 3650 4750 3800 4760
rect 3950 4750 4950 4760
rect 7400 4750 7650 4760
rect 9750 4750 9850 4760
rect 450 4740 550 4750
rect 1150 4740 2400 4750
rect 3600 4740 3800 4750
rect 3850 4740 5050 4750
rect 7450 4740 7600 4750
rect 8450 4740 8500 4750
rect 8700 4740 8750 4750
rect 9500 4740 9800 4750
rect 450 4730 550 4740
rect 1150 4730 2400 4740
rect 3600 4730 3800 4740
rect 3850 4730 5050 4740
rect 7450 4730 7600 4740
rect 8450 4730 8500 4740
rect 8700 4730 8750 4740
rect 9500 4730 9800 4740
rect 450 4720 550 4730
rect 1150 4720 2400 4730
rect 3600 4720 3800 4730
rect 3850 4720 5050 4730
rect 7450 4720 7600 4730
rect 8450 4720 8500 4730
rect 8700 4720 8750 4730
rect 9500 4720 9800 4730
rect 450 4710 550 4720
rect 1150 4710 2400 4720
rect 3600 4710 3800 4720
rect 3850 4710 5050 4720
rect 7450 4710 7600 4720
rect 8450 4710 8500 4720
rect 8700 4710 8750 4720
rect 9500 4710 9800 4720
rect 450 4700 550 4710
rect 1150 4700 2400 4710
rect 3600 4700 3800 4710
rect 3850 4700 5050 4710
rect 7450 4700 7600 4710
rect 8450 4700 8500 4710
rect 8700 4700 8750 4710
rect 9500 4700 9800 4710
rect 550 4690 750 4700
rect 1200 4690 2450 4700
rect 3550 4690 5050 4700
rect 8400 4690 8450 4700
rect 8700 4690 8750 4700
rect 9350 4690 9750 4700
rect 550 4680 750 4690
rect 1200 4680 2450 4690
rect 3550 4680 5050 4690
rect 8400 4680 8450 4690
rect 8700 4680 8750 4690
rect 9350 4680 9750 4690
rect 550 4670 750 4680
rect 1200 4670 2450 4680
rect 3550 4670 5050 4680
rect 8400 4670 8450 4680
rect 8700 4670 8750 4680
rect 9350 4670 9750 4680
rect 550 4660 750 4670
rect 1200 4660 2450 4670
rect 3550 4660 5050 4670
rect 8400 4660 8450 4670
rect 8700 4660 8750 4670
rect 9350 4660 9750 4670
rect 550 4650 750 4660
rect 1200 4650 2450 4660
rect 3550 4650 5050 4660
rect 8400 4650 8450 4660
rect 8700 4650 8750 4660
rect 9350 4650 9750 4660
rect 650 4640 850 4650
rect 1200 4640 2550 4650
rect 3500 4640 5100 4650
rect 8700 4640 8750 4650
rect 9300 4640 9700 4650
rect 650 4630 850 4640
rect 1200 4630 2550 4640
rect 3500 4630 5100 4640
rect 8700 4630 8750 4640
rect 9300 4630 9700 4640
rect 650 4620 850 4630
rect 1200 4620 2550 4630
rect 3500 4620 5100 4630
rect 8700 4620 8750 4630
rect 9300 4620 9700 4630
rect 650 4610 850 4620
rect 1200 4610 2550 4620
rect 3500 4610 5100 4620
rect 8700 4610 8750 4620
rect 9300 4610 9700 4620
rect 650 4600 850 4610
rect 1200 4600 2550 4610
rect 3500 4600 5100 4610
rect 8700 4600 8750 4610
rect 9300 4600 9700 4610
rect 700 4590 900 4600
rect 1250 4590 3000 4600
rect 3050 4590 3100 4600
rect 3500 4590 5200 4600
rect 5700 4590 5750 4600
rect 6350 4590 6450 4600
rect 8700 4590 8800 4600
rect 9300 4590 9650 4600
rect 700 4580 900 4590
rect 1250 4580 3000 4590
rect 3050 4580 3100 4590
rect 3500 4580 5200 4590
rect 5700 4580 5750 4590
rect 6350 4580 6450 4590
rect 8700 4580 8800 4590
rect 9300 4580 9650 4590
rect 700 4570 900 4580
rect 1250 4570 3000 4580
rect 3050 4570 3100 4580
rect 3500 4570 5200 4580
rect 5700 4570 5750 4580
rect 6350 4570 6450 4580
rect 8700 4570 8800 4580
rect 9300 4570 9650 4580
rect 700 4560 900 4570
rect 1250 4560 3000 4570
rect 3050 4560 3100 4570
rect 3500 4560 5200 4570
rect 5700 4560 5750 4570
rect 6350 4560 6450 4570
rect 8700 4560 8800 4570
rect 9300 4560 9650 4570
rect 700 4550 900 4560
rect 1250 4550 3000 4560
rect 3050 4550 3100 4560
rect 3500 4550 5200 4560
rect 5700 4550 5750 4560
rect 6350 4550 6450 4560
rect 8700 4550 8800 4560
rect 9300 4550 9650 4560
rect 750 4540 950 4550
rect 1200 4540 2950 4550
rect 3100 4540 3150 4550
rect 3500 4540 3850 4550
rect 3950 4540 5200 4550
rect 6350 4540 6400 4550
rect 8700 4540 8900 4550
rect 9300 4540 9600 4550
rect 750 4530 950 4540
rect 1200 4530 2950 4540
rect 3100 4530 3150 4540
rect 3500 4530 3850 4540
rect 3950 4530 5200 4540
rect 6350 4530 6400 4540
rect 8700 4530 8900 4540
rect 9300 4530 9600 4540
rect 750 4520 950 4530
rect 1200 4520 2950 4530
rect 3100 4520 3150 4530
rect 3500 4520 3850 4530
rect 3950 4520 5200 4530
rect 6350 4520 6400 4530
rect 8700 4520 8900 4530
rect 9300 4520 9600 4530
rect 750 4510 950 4520
rect 1200 4510 2950 4520
rect 3100 4510 3150 4520
rect 3500 4510 3850 4520
rect 3950 4510 5200 4520
rect 6350 4510 6400 4520
rect 8700 4510 8900 4520
rect 9300 4510 9600 4520
rect 750 4500 950 4510
rect 1200 4500 2950 4510
rect 3100 4500 3150 4510
rect 3500 4500 3850 4510
rect 3950 4500 5200 4510
rect 6350 4500 6400 4510
rect 8700 4500 8900 4510
rect 9300 4500 9600 4510
rect 650 4490 1000 4500
rect 1200 4490 2800 4500
rect 2900 4490 2950 4500
rect 3450 4490 3850 4500
rect 3950 4490 5250 4500
rect 6300 4490 6350 4500
rect 7550 4490 7700 4500
rect 8450 4490 8850 4500
rect 9250 4490 9550 4500
rect 650 4480 1000 4490
rect 1200 4480 2800 4490
rect 2900 4480 2950 4490
rect 3450 4480 3850 4490
rect 3950 4480 5250 4490
rect 6300 4480 6350 4490
rect 7550 4480 7700 4490
rect 8450 4480 8850 4490
rect 9250 4480 9550 4490
rect 650 4470 1000 4480
rect 1200 4470 2800 4480
rect 2900 4470 2950 4480
rect 3450 4470 3850 4480
rect 3950 4470 5250 4480
rect 6300 4470 6350 4480
rect 7550 4470 7700 4480
rect 8450 4470 8850 4480
rect 9250 4470 9550 4480
rect 650 4460 1000 4470
rect 1200 4460 2800 4470
rect 2900 4460 2950 4470
rect 3450 4460 3850 4470
rect 3950 4460 5250 4470
rect 6300 4460 6350 4470
rect 7550 4460 7700 4470
rect 8450 4460 8850 4470
rect 9250 4460 9550 4470
rect 650 4450 1000 4460
rect 1200 4450 2800 4460
rect 2900 4450 2950 4460
rect 3450 4450 3850 4460
rect 3950 4450 5250 4460
rect 6300 4450 6350 4460
rect 7550 4450 7700 4460
rect 8450 4450 8850 4460
rect 9250 4450 9550 4460
rect 450 4440 1050 4450
rect 1150 4440 2800 4450
rect 2900 4440 2950 4450
rect 3450 4440 3850 4450
rect 3950 4440 4250 4450
rect 4300 4440 4600 4450
rect 4750 4440 5250 4450
rect 7450 4440 7750 4450
rect 8350 4440 8650 4450
rect 8750 4440 8800 4450
rect 9250 4440 9500 4450
rect 9950 4440 9990 4450
rect 450 4430 1050 4440
rect 1150 4430 2800 4440
rect 2900 4430 2950 4440
rect 3450 4430 3850 4440
rect 3950 4430 4250 4440
rect 4300 4430 4600 4440
rect 4750 4430 5250 4440
rect 7450 4430 7750 4440
rect 8350 4430 8650 4440
rect 8750 4430 8800 4440
rect 9250 4430 9500 4440
rect 9950 4430 9990 4440
rect 450 4420 1050 4430
rect 1150 4420 2800 4430
rect 2900 4420 2950 4430
rect 3450 4420 3850 4430
rect 3950 4420 4250 4430
rect 4300 4420 4600 4430
rect 4750 4420 5250 4430
rect 7450 4420 7750 4430
rect 8350 4420 8650 4430
rect 8750 4420 8800 4430
rect 9250 4420 9500 4430
rect 9950 4420 9990 4430
rect 450 4410 1050 4420
rect 1150 4410 2800 4420
rect 2900 4410 2950 4420
rect 3450 4410 3850 4420
rect 3950 4410 4250 4420
rect 4300 4410 4600 4420
rect 4750 4410 5250 4420
rect 7450 4410 7750 4420
rect 8350 4410 8650 4420
rect 8750 4410 8800 4420
rect 9250 4410 9500 4420
rect 9950 4410 9990 4420
rect 450 4400 1050 4410
rect 1150 4400 2800 4410
rect 2900 4400 2950 4410
rect 3450 4400 3850 4410
rect 3950 4400 4250 4410
rect 4300 4400 4600 4410
rect 4750 4400 5250 4410
rect 7450 4400 7750 4410
rect 8350 4400 8650 4410
rect 8750 4400 8800 4410
rect 9250 4400 9500 4410
rect 9950 4400 9990 4410
rect 250 4390 2800 4400
rect 3400 4390 3800 4400
rect 3950 4390 4250 4400
rect 4350 4390 4550 4400
rect 4950 4390 5300 4400
rect 7450 4390 7750 4400
rect 8200 4390 8450 4400
rect 8750 4390 8800 4400
rect 9250 4390 9450 4400
rect 250 4380 2800 4390
rect 3400 4380 3800 4390
rect 3950 4380 4250 4390
rect 4350 4380 4550 4390
rect 4950 4380 5300 4390
rect 7450 4380 7750 4390
rect 8200 4380 8450 4390
rect 8750 4380 8800 4390
rect 9250 4380 9450 4390
rect 250 4370 2800 4380
rect 3400 4370 3800 4380
rect 3950 4370 4250 4380
rect 4350 4370 4550 4380
rect 4950 4370 5300 4380
rect 7450 4370 7750 4380
rect 8200 4370 8450 4380
rect 8750 4370 8800 4380
rect 9250 4370 9450 4380
rect 250 4360 2800 4370
rect 3400 4360 3800 4370
rect 3950 4360 4250 4370
rect 4350 4360 4550 4370
rect 4950 4360 5300 4370
rect 7450 4360 7750 4370
rect 8200 4360 8450 4370
rect 8750 4360 8800 4370
rect 9250 4360 9450 4370
rect 250 4350 2800 4360
rect 3400 4350 3800 4360
rect 3950 4350 4250 4360
rect 4350 4350 4550 4360
rect 4950 4350 5300 4360
rect 7450 4350 7750 4360
rect 8200 4350 8450 4360
rect 8750 4350 8800 4360
rect 9250 4350 9450 4360
rect 250 4340 2800 4350
rect 3400 4340 4150 4350
rect 4350 4340 4500 4350
rect 4950 4340 5300 4350
rect 7450 4340 7800 4350
rect 7900 4340 8150 4350
rect 8200 4340 8400 4350
rect 9250 4340 9400 4350
rect 250 4330 2800 4340
rect 3400 4330 4150 4340
rect 4350 4330 4500 4340
rect 4950 4330 5300 4340
rect 7450 4330 7800 4340
rect 7900 4330 8150 4340
rect 8200 4330 8400 4340
rect 9250 4330 9400 4340
rect 250 4320 2800 4330
rect 3400 4320 4150 4330
rect 4350 4320 4500 4330
rect 4950 4320 5300 4330
rect 7450 4320 7800 4330
rect 7900 4320 8150 4330
rect 8200 4320 8400 4330
rect 9250 4320 9400 4330
rect 250 4310 2800 4320
rect 3400 4310 4150 4320
rect 4350 4310 4500 4320
rect 4950 4310 5300 4320
rect 7450 4310 7800 4320
rect 7900 4310 8150 4320
rect 8200 4310 8400 4320
rect 9250 4310 9400 4320
rect 250 4300 2800 4310
rect 3400 4300 4150 4310
rect 4350 4300 4500 4310
rect 4950 4300 5300 4310
rect 7450 4300 7800 4310
rect 7900 4300 8150 4310
rect 8200 4300 8400 4310
rect 9250 4300 9400 4310
rect 100 4290 2800 4300
rect 3300 4290 4100 4300
rect 4350 4290 4450 4300
rect 5000 4290 5300 4300
rect 7450 4290 8150 4300
rect 8200 4290 8400 4300
rect 8750 4290 8800 4300
rect 9250 4290 9350 4300
rect 100 4280 2800 4290
rect 3300 4280 4100 4290
rect 4350 4280 4450 4290
rect 5000 4280 5300 4290
rect 7450 4280 8150 4290
rect 8200 4280 8400 4290
rect 8750 4280 8800 4290
rect 9250 4280 9350 4290
rect 100 4270 2800 4280
rect 3300 4270 4100 4280
rect 4350 4270 4450 4280
rect 5000 4270 5300 4280
rect 7450 4270 8150 4280
rect 8200 4270 8400 4280
rect 8750 4270 8800 4280
rect 9250 4270 9350 4280
rect 100 4260 2800 4270
rect 3300 4260 4100 4270
rect 4350 4260 4450 4270
rect 5000 4260 5300 4270
rect 7450 4260 8150 4270
rect 8200 4260 8400 4270
rect 8750 4260 8800 4270
rect 9250 4260 9350 4270
rect 100 4250 2800 4260
rect 3300 4250 4100 4260
rect 4350 4250 4450 4260
rect 5000 4250 5300 4260
rect 7450 4250 8150 4260
rect 8200 4250 8400 4260
rect 8750 4250 8800 4260
rect 9250 4250 9350 4260
rect 150 4240 2750 4250
rect 3300 4240 4100 4250
rect 5050 4240 5350 4250
rect 7500 4240 8150 4250
rect 8200 4240 8400 4250
rect 8550 4240 8800 4250
rect 150 4230 2750 4240
rect 3300 4230 4100 4240
rect 5050 4230 5350 4240
rect 7500 4230 8150 4240
rect 8200 4230 8400 4240
rect 8550 4230 8800 4240
rect 150 4220 2750 4230
rect 3300 4220 4100 4230
rect 5050 4220 5350 4230
rect 7500 4220 8150 4230
rect 8200 4220 8400 4230
rect 8550 4220 8800 4230
rect 150 4210 2750 4220
rect 3300 4210 4100 4220
rect 5050 4210 5350 4220
rect 7500 4210 8150 4220
rect 8200 4210 8400 4220
rect 8550 4210 8800 4220
rect 150 4200 2750 4210
rect 3300 4200 4100 4210
rect 5050 4200 5350 4210
rect 7500 4200 8150 4210
rect 8200 4200 8400 4210
rect 8550 4200 8800 4210
rect 150 4190 2550 4200
rect 3300 4190 4050 4200
rect 5050 4190 5350 4200
rect 7500 4190 8750 4200
rect 150 4180 2550 4190
rect 3300 4180 4050 4190
rect 5050 4180 5350 4190
rect 7500 4180 8750 4190
rect 150 4170 2550 4180
rect 3300 4170 4050 4180
rect 5050 4170 5350 4180
rect 7500 4170 8750 4180
rect 150 4160 2550 4170
rect 3300 4160 4050 4170
rect 5050 4160 5350 4170
rect 7500 4160 8750 4170
rect 150 4150 2550 4160
rect 3300 4150 4050 4160
rect 5050 4150 5350 4160
rect 7500 4150 8750 4160
rect 0 4140 50 4150
rect 150 4140 2600 4150
rect 3350 4140 4050 4150
rect 5150 4140 5400 4150
rect 7550 4140 8750 4150
rect 0 4130 50 4140
rect 150 4130 2600 4140
rect 3350 4130 4050 4140
rect 5150 4130 5400 4140
rect 7550 4130 8750 4140
rect 0 4120 50 4130
rect 150 4120 2600 4130
rect 3350 4120 4050 4130
rect 5150 4120 5400 4130
rect 7550 4120 8750 4130
rect 0 4110 50 4120
rect 150 4110 2600 4120
rect 3350 4110 4050 4120
rect 5150 4110 5400 4120
rect 7550 4110 8750 4120
rect 0 4100 50 4110
rect 150 4100 2600 4110
rect 3350 4100 4050 4110
rect 5150 4100 5400 4110
rect 7550 4100 8750 4110
rect 0 4090 100 4100
rect 150 4090 2600 4100
rect 3300 4090 4000 4100
rect 5150 4090 5400 4100
rect 5550 4090 5600 4100
rect 7300 4090 7450 4100
rect 7700 4090 8550 4100
rect 8700 4090 8750 4100
rect 0 4080 100 4090
rect 150 4080 2600 4090
rect 3300 4080 4000 4090
rect 5150 4080 5400 4090
rect 5550 4080 5600 4090
rect 7300 4080 7450 4090
rect 7700 4080 8550 4090
rect 8700 4080 8750 4090
rect 0 4070 100 4080
rect 150 4070 2600 4080
rect 3300 4070 4000 4080
rect 5150 4070 5400 4080
rect 5550 4070 5600 4080
rect 7300 4070 7450 4080
rect 7700 4070 8550 4080
rect 8700 4070 8750 4080
rect 0 4060 100 4070
rect 150 4060 2600 4070
rect 3300 4060 4000 4070
rect 5150 4060 5400 4070
rect 5550 4060 5600 4070
rect 7300 4060 7450 4070
rect 7700 4060 8550 4070
rect 8700 4060 8750 4070
rect 0 4050 100 4060
rect 150 4050 2600 4060
rect 3300 4050 4000 4060
rect 5150 4050 5400 4060
rect 5550 4050 5600 4060
rect 7300 4050 7450 4060
rect 7700 4050 8550 4060
rect 8700 4050 8750 4060
rect 0 4040 2600 4050
rect 3300 4040 4000 4050
rect 5200 4040 5350 4050
rect 5550 4040 5650 4050
rect 7250 4040 7600 4050
rect 7850 4040 8300 4050
rect 0 4030 2600 4040
rect 3300 4030 4000 4040
rect 5200 4030 5350 4040
rect 5550 4030 5650 4040
rect 7250 4030 7600 4040
rect 7850 4030 8300 4040
rect 0 4020 2600 4030
rect 3300 4020 4000 4030
rect 5200 4020 5350 4030
rect 5550 4020 5650 4030
rect 7250 4020 7600 4030
rect 7850 4020 8300 4030
rect 0 4010 2600 4020
rect 3300 4010 4000 4020
rect 5200 4010 5350 4020
rect 5550 4010 5650 4020
rect 7250 4010 7600 4020
rect 7850 4010 8300 4020
rect 0 4000 2600 4010
rect 3300 4000 4000 4010
rect 5200 4000 5350 4010
rect 5550 4000 5650 4010
rect 7250 4000 7600 4010
rect 7850 4000 8300 4010
rect 0 3990 2600 4000
rect 3300 3990 3900 4000
rect 5200 3990 5350 4000
rect 5550 3990 5750 4000
rect 7200 3990 7750 4000
rect 7950 3990 8100 4000
rect 0 3980 2600 3990
rect 3300 3980 3900 3990
rect 5200 3980 5350 3990
rect 5550 3980 5750 3990
rect 7200 3980 7750 3990
rect 7950 3980 8100 3990
rect 0 3970 2600 3980
rect 3300 3970 3900 3980
rect 5200 3970 5350 3980
rect 5550 3970 5750 3980
rect 7200 3970 7750 3980
rect 7950 3970 8100 3980
rect 0 3960 2600 3970
rect 3300 3960 3900 3970
rect 5200 3960 5350 3970
rect 5550 3960 5750 3970
rect 7200 3960 7750 3970
rect 7950 3960 8100 3970
rect 0 3950 2600 3960
rect 3300 3950 3900 3960
rect 5200 3950 5350 3960
rect 5550 3950 5750 3960
rect 7200 3950 7750 3960
rect 7950 3950 8100 3960
rect 0 3940 2600 3950
rect 3300 3940 3850 3950
rect 5250 3940 5400 3950
rect 5500 3940 5900 3950
rect 7200 3940 7850 3950
rect 0 3930 2600 3940
rect 3300 3930 3850 3940
rect 5250 3930 5400 3940
rect 5500 3930 5900 3940
rect 7200 3930 7850 3940
rect 0 3920 2600 3930
rect 3300 3920 3850 3930
rect 5250 3920 5400 3930
rect 5500 3920 5900 3930
rect 7200 3920 7850 3930
rect 0 3910 2600 3920
rect 3300 3910 3850 3920
rect 5250 3910 5400 3920
rect 5500 3910 5900 3920
rect 7200 3910 7850 3920
rect 0 3900 2600 3910
rect 3300 3900 3850 3910
rect 5250 3900 5400 3910
rect 5500 3900 5900 3910
rect 7200 3900 7850 3910
rect 0 3890 2550 3900
rect 3350 3890 3850 3900
rect 5300 3890 6000 3900
rect 7200 3890 7950 3900
rect 8100 3890 8150 3900
rect 0 3880 2550 3890
rect 3350 3880 3850 3890
rect 5300 3880 6000 3890
rect 7200 3880 7950 3890
rect 8100 3880 8150 3890
rect 0 3870 2550 3880
rect 3350 3870 3850 3880
rect 5300 3870 6000 3880
rect 7200 3870 7950 3880
rect 8100 3870 8150 3880
rect 0 3860 2550 3870
rect 3350 3860 3850 3870
rect 5300 3860 6000 3870
rect 7200 3860 7950 3870
rect 8100 3860 8150 3870
rect 0 3850 2550 3860
rect 3350 3850 3850 3860
rect 5300 3850 6000 3860
rect 7200 3850 7950 3860
rect 8100 3850 8150 3860
rect 0 3840 2400 3850
rect 2450 3840 2550 3850
rect 3300 3840 3850 3850
rect 4150 3840 4200 3850
rect 5300 3840 5950 3850
rect 7150 3840 8000 3850
rect 0 3830 2400 3840
rect 2450 3830 2550 3840
rect 3300 3830 3850 3840
rect 4150 3830 4200 3840
rect 5300 3830 5950 3840
rect 7150 3830 8000 3840
rect 0 3820 2400 3830
rect 2450 3820 2550 3830
rect 3300 3820 3850 3830
rect 4150 3820 4200 3830
rect 5300 3820 5950 3830
rect 7150 3820 8000 3830
rect 0 3810 2400 3820
rect 2450 3810 2550 3820
rect 3300 3810 3850 3820
rect 4150 3810 4200 3820
rect 5300 3810 5950 3820
rect 7150 3810 8000 3820
rect 0 3800 2400 3810
rect 2450 3800 2550 3810
rect 3300 3800 3850 3810
rect 4150 3800 4200 3810
rect 5300 3800 5950 3810
rect 7150 3800 8000 3810
rect 0 3790 2550 3800
rect 3350 3790 3850 3800
rect 5300 3790 6000 3800
rect 7100 3790 8100 3800
rect 0 3780 2550 3790
rect 3350 3780 3850 3790
rect 5300 3780 6000 3790
rect 7100 3780 8100 3790
rect 0 3770 2550 3780
rect 3350 3770 3850 3780
rect 5300 3770 6000 3780
rect 7100 3770 8100 3780
rect 0 3760 2550 3770
rect 3350 3760 3850 3770
rect 5300 3760 6000 3770
rect 7100 3760 8100 3770
rect 0 3750 2550 3760
rect 3350 3750 3850 3760
rect 5300 3750 6000 3760
rect 7100 3750 8100 3760
rect 0 3740 1600 3750
rect 1700 3740 2700 3750
rect 3350 3740 3850 3750
rect 5350 3740 6050 3750
rect 7100 3740 8150 3750
rect 0 3730 1600 3740
rect 1700 3730 2700 3740
rect 3350 3730 3850 3740
rect 5350 3730 6050 3740
rect 7100 3730 8150 3740
rect 0 3720 1600 3730
rect 1700 3720 2700 3730
rect 3350 3720 3850 3730
rect 5350 3720 6050 3730
rect 7100 3720 8150 3730
rect 0 3710 1600 3720
rect 1700 3710 2700 3720
rect 3350 3710 3850 3720
rect 5350 3710 6050 3720
rect 7100 3710 8150 3720
rect 0 3700 1600 3710
rect 1700 3700 2700 3710
rect 3350 3700 3850 3710
rect 5350 3700 6050 3710
rect 7100 3700 8150 3710
rect 50 3690 1600 3700
rect 1700 3690 2850 3700
rect 3350 3690 3850 3700
rect 5350 3690 6050 3700
rect 7050 3690 8150 3700
rect 50 3680 1600 3690
rect 1700 3680 2850 3690
rect 3350 3680 3850 3690
rect 5350 3680 6050 3690
rect 7050 3680 8150 3690
rect 50 3670 1600 3680
rect 1700 3670 2850 3680
rect 3350 3670 3850 3680
rect 5350 3670 6050 3680
rect 7050 3670 8150 3680
rect 50 3660 1600 3670
rect 1700 3660 2850 3670
rect 3350 3660 3850 3670
rect 5350 3660 6050 3670
rect 7050 3660 8150 3670
rect 50 3650 1600 3660
rect 1700 3650 2850 3660
rect 3350 3650 3850 3660
rect 5350 3650 6050 3660
rect 7050 3650 8150 3660
rect 0 3640 3050 3650
rect 3400 3640 3900 3650
rect 5350 3640 6150 3650
rect 7000 3640 8200 3650
rect 0 3630 3050 3640
rect 3400 3630 3900 3640
rect 5350 3630 6150 3640
rect 7000 3630 8200 3640
rect 0 3620 3050 3630
rect 3400 3620 3900 3630
rect 5350 3620 6150 3630
rect 7000 3620 8200 3630
rect 0 3610 3050 3620
rect 3400 3610 3900 3620
rect 5350 3610 6150 3620
rect 7000 3610 8200 3620
rect 0 3600 3050 3610
rect 3400 3600 3900 3610
rect 5350 3600 6150 3610
rect 7000 3600 8200 3610
rect 0 3590 3200 3600
rect 3450 3590 3900 3600
rect 5350 3590 6150 3600
rect 7000 3590 8250 3600
rect 0 3580 3200 3590
rect 3450 3580 3900 3590
rect 5350 3580 6150 3590
rect 7000 3580 8250 3590
rect 0 3570 3200 3580
rect 3450 3570 3900 3580
rect 5350 3570 6150 3580
rect 7000 3570 8250 3580
rect 0 3560 3200 3570
rect 3450 3560 3900 3570
rect 5350 3560 6150 3570
rect 7000 3560 8250 3570
rect 0 3550 3200 3560
rect 3450 3550 3900 3560
rect 5350 3550 6150 3560
rect 7000 3550 8250 3560
rect 0 3540 1400 3550
rect 1500 3540 2400 3550
rect 2750 3540 3250 3550
rect 3450 3540 3900 3550
rect 5400 3540 6150 3550
rect 6950 3540 8300 3550
rect 0 3530 1400 3540
rect 1500 3530 2400 3540
rect 2750 3530 3250 3540
rect 3450 3530 3900 3540
rect 5400 3530 6150 3540
rect 6950 3530 8300 3540
rect 0 3520 1400 3530
rect 1500 3520 2400 3530
rect 2750 3520 3250 3530
rect 3450 3520 3900 3530
rect 5400 3520 6150 3530
rect 6950 3520 8300 3530
rect 0 3510 1400 3520
rect 1500 3510 2400 3520
rect 2750 3510 3250 3520
rect 3450 3510 3900 3520
rect 5400 3510 6150 3520
rect 6950 3510 8300 3520
rect 0 3500 1400 3510
rect 1500 3500 2400 3510
rect 2750 3500 3250 3510
rect 3450 3500 3900 3510
rect 5400 3500 6150 3510
rect 6950 3500 8300 3510
rect 0 3490 1400 3500
rect 1450 3490 2250 3500
rect 2900 3490 3300 3500
rect 3450 3490 3900 3500
rect 5400 3490 6150 3500
rect 6900 3490 8350 3500
rect 0 3480 1400 3490
rect 1450 3480 2250 3490
rect 2900 3480 3300 3490
rect 3450 3480 3900 3490
rect 5400 3480 6150 3490
rect 6900 3480 8350 3490
rect 0 3470 1400 3480
rect 1450 3470 2250 3480
rect 2900 3470 3300 3480
rect 3450 3470 3900 3480
rect 5400 3470 6150 3480
rect 6900 3470 8350 3480
rect 0 3460 1400 3470
rect 1450 3460 2250 3470
rect 2900 3460 3300 3470
rect 3450 3460 3900 3470
rect 5400 3460 6150 3470
rect 6900 3460 8350 3470
rect 0 3450 1400 3460
rect 1450 3450 2250 3460
rect 2900 3450 3300 3460
rect 3450 3450 3900 3460
rect 5400 3450 6150 3460
rect 6900 3450 8350 3460
rect 0 3440 1350 3450
rect 1450 3440 2200 3450
rect 3050 3440 3350 3450
rect 3450 3440 3900 3450
rect 5350 3440 5850 3450
rect 6050 3440 6100 3450
rect 6850 3440 8400 3450
rect 0 3430 1350 3440
rect 1450 3430 2200 3440
rect 3050 3430 3350 3440
rect 3450 3430 3900 3440
rect 5350 3430 5850 3440
rect 6050 3430 6100 3440
rect 6850 3430 8400 3440
rect 0 3420 1350 3430
rect 1450 3420 2200 3430
rect 3050 3420 3350 3430
rect 3450 3420 3900 3430
rect 5350 3420 5850 3430
rect 6050 3420 6100 3430
rect 6850 3420 8400 3430
rect 0 3410 1350 3420
rect 1450 3410 2200 3420
rect 3050 3410 3350 3420
rect 3450 3410 3900 3420
rect 5350 3410 5850 3420
rect 6050 3410 6100 3420
rect 6850 3410 8400 3420
rect 0 3400 1350 3410
rect 1450 3400 2200 3410
rect 3050 3400 3350 3410
rect 3450 3400 3900 3410
rect 5350 3400 5850 3410
rect 6050 3400 6100 3410
rect 6850 3400 8400 3410
rect 0 3390 1350 3400
rect 1450 3390 2100 3400
rect 3100 3390 3450 3400
rect 3600 3390 3950 3400
rect 5350 3390 5650 3400
rect 5750 3390 5850 3400
rect 6050 3390 6100 3400
rect 6800 3390 8450 3400
rect 0 3380 1350 3390
rect 1450 3380 2100 3390
rect 3100 3380 3450 3390
rect 3600 3380 3950 3390
rect 5350 3380 5650 3390
rect 5750 3380 5850 3390
rect 6050 3380 6100 3390
rect 6800 3380 8450 3390
rect 0 3370 1350 3380
rect 1450 3370 2100 3380
rect 3100 3370 3450 3380
rect 3600 3370 3950 3380
rect 5350 3370 5650 3380
rect 5750 3370 5850 3380
rect 6050 3370 6100 3380
rect 6800 3370 8450 3380
rect 0 3360 1350 3370
rect 1450 3360 2100 3370
rect 3100 3360 3450 3370
rect 3600 3360 3950 3370
rect 5350 3360 5650 3370
rect 5750 3360 5850 3370
rect 6050 3360 6100 3370
rect 6800 3360 8450 3370
rect 0 3350 1350 3360
rect 1450 3350 2100 3360
rect 3100 3350 3450 3360
rect 3600 3350 3950 3360
rect 5350 3350 5650 3360
rect 5750 3350 5850 3360
rect 6050 3350 6100 3360
rect 6800 3350 8450 3360
rect 0 3340 1300 3350
rect 1400 3340 2100 3350
rect 3150 3340 3450 3350
rect 3650 3340 3950 3350
rect 5350 3340 5600 3350
rect 6750 3340 8450 3350
rect 0 3330 1300 3340
rect 1400 3330 2100 3340
rect 3150 3330 3450 3340
rect 3650 3330 3950 3340
rect 5350 3330 5600 3340
rect 6750 3330 8450 3340
rect 0 3320 1300 3330
rect 1400 3320 2100 3330
rect 3150 3320 3450 3330
rect 3650 3320 3950 3330
rect 5350 3320 5600 3330
rect 6750 3320 8450 3330
rect 0 3310 1300 3320
rect 1400 3310 2100 3320
rect 3150 3310 3450 3320
rect 3650 3310 3950 3320
rect 5350 3310 5600 3320
rect 6750 3310 8450 3320
rect 0 3300 1300 3310
rect 1400 3300 2100 3310
rect 3150 3300 3450 3310
rect 3650 3300 3950 3310
rect 5350 3300 5600 3310
rect 6750 3300 8450 3310
rect 0 3290 1300 3300
rect 1400 3290 2050 3300
rect 3200 3290 3500 3300
rect 3650 3290 4000 3300
rect 5350 3290 5600 3300
rect 6700 3290 8400 3300
rect 0 3280 1300 3290
rect 1400 3280 2050 3290
rect 3200 3280 3500 3290
rect 3650 3280 4000 3290
rect 5350 3280 5600 3290
rect 6700 3280 8400 3290
rect 0 3270 1300 3280
rect 1400 3270 2050 3280
rect 3200 3270 3500 3280
rect 3650 3270 4000 3280
rect 5350 3270 5600 3280
rect 6700 3270 8400 3280
rect 0 3260 1300 3270
rect 1400 3260 2050 3270
rect 3200 3260 3500 3270
rect 3650 3260 4000 3270
rect 5350 3260 5600 3270
rect 6700 3260 8400 3270
rect 0 3250 1300 3260
rect 1400 3250 2050 3260
rect 3200 3250 3500 3260
rect 3650 3250 4000 3260
rect 5350 3250 5600 3260
rect 6700 3250 8400 3260
rect 0 3240 1300 3250
rect 1400 3240 2050 3250
rect 3200 3240 3550 3250
rect 3650 3240 4050 3250
rect 5350 3240 5650 3250
rect 6700 3240 8400 3250
rect 0 3230 1300 3240
rect 1400 3230 2050 3240
rect 3200 3230 3550 3240
rect 3650 3230 4050 3240
rect 5350 3230 5650 3240
rect 6700 3230 8400 3240
rect 0 3220 1300 3230
rect 1400 3220 2050 3230
rect 3200 3220 3550 3230
rect 3650 3220 4050 3230
rect 5350 3220 5650 3230
rect 6700 3220 8400 3230
rect 0 3210 1300 3220
rect 1400 3210 2050 3220
rect 3200 3210 3550 3220
rect 3650 3210 4050 3220
rect 5350 3210 5650 3220
rect 6700 3210 8400 3220
rect 0 3200 1300 3210
rect 1400 3200 2050 3210
rect 3200 3200 3550 3210
rect 3650 3200 4050 3210
rect 5350 3200 5650 3210
rect 6700 3200 8400 3210
rect 0 3190 1250 3200
rect 1350 3190 2000 3200
rect 3200 3190 4050 3200
rect 5300 3190 5700 3200
rect 6500 3190 6550 3200
rect 6700 3190 8350 3200
rect 0 3180 1250 3190
rect 1350 3180 2000 3190
rect 3200 3180 4050 3190
rect 5300 3180 5700 3190
rect 6500 3180 6550 3190
rect 6700 3180 8350 3190
rect 0 3170 1250 3180
rect 1350 3170 2000 3180
rect 3200 3170 4050 3180
rect 5300 3170 5700 3180
rect 6500 3170 6550 3180
rect 6700 3170 8350 3180
rect 0 3160 1250 3170
rect 1350 3160 2000 3170
rect 3200 3160 4050 3170
rect 5300 3160 5700 3170
rect 6500 3160 6550 3170
rect 6700 3160 8350 3170
rect 0 3150 1250 3160
rect 1350 3150 2000 3160
rect 3200 3150 4050 3160
rect 5300 3150 5700 3160
rect 6500 3150 6550 3160
rect 6700 3150 8350 3160
rect 0 3140 1250 3150
rect 1350 3140 2000 3150
rect 3250 3140 3750 3150
rect 4000 3140 4050 3150
rect 5300 3140 5800 3150
rect 6350 3140 6550 3150
rect 6650 3140 8350 3150
rect 9150 3140 9200 3150
rect 0 3130 1250 3140
rect 1350 3130 2000 3140
rect 3250 3130 3750 3140
rect 4000 3130 4050 3140
rect 5300 3130 5800 3140
rect 6350 3130 6550 3140
rect 6650 3130 8350 3140
rect 9150 3130 9200 3140
rect 0 3120 1250 3130
rect 1350 3120 2000 3130
rect 3250 3120 3750 3130
rect 4000 3120 4050 3130
rect 5300 3120 5800 3130
rect 6350 3120 6550 3130
rect 6650 3120 8350 3130
rect 9150 3120 9200 3130
rect 0 3110 1250 3120
rect 1350 3110 2000 3120
rect 3250 3110 3750 3120
rect 4000 3110 4050 3120
rect 5300 3110 5800 3120
rect 6350 3110 6550 3120
rect 6650 3110 8350 3120
rect 9150 3110 9200 3120
rect 0 3100 1250 3110
rect 1350 3100 2000 3110
rect 3250 3100 3750 3110
rect 4000 3100 4050 3110
rect 5300 3100 5800 3110
rect 6350 3100 6550 3110
rect 6650 3100 8350 3110
rect 9150 3100 9200 3110
rect 0 3090 1200 3100
rect 1350 3090 2000 3100
rect 3200 3090 3750 3100
rect 4050 3090 4100 3100
rect 5300 3090 6550 3100
rect 6650 3090 8300 3100
rect 9100 3090 9200 3100
rect 0 3080 1200 3090
rect 1350 3080 2000 3090
rect 3200 3080 3750 3090
rect 4050 3080 4100 3090
rect 5300 3080 6550 3090
rect 6650 3080 8300 3090
rect 9100 3080 9200 3090
rect 0 3070 1200 3080
rect 1350 3070 2000 3080
rect 3200 3070 3750 3080
rect 4050 3070 4100 3080
rect 5300 3070 6550 3080
rect 6650 3070 8300 3080
rect 9100 3070 9200 3080
rect 0 3060 1200 3070
rect 1350 3060 2000 3070
rect 3200 3060 3750 3070
rect 4050 3060 4100 3070
rect 5300 3060 6550 3070
rect 6650 3060 8300 3070
rect 9100 3060 9200 3070
rect 0 3050 1200 3060
rect 1350 3050 2000 3060
rect 3200 3050 3750 3060
rect 4050 3050 4100 3060
rect 5300 3050 6550 3060
rect 6650 3050 8300 3060
rect 9100 3050 9200 3060
rect 0 3040 1200 3050
rect 1300 3040 2000 3050
rect 3200 3040 3700 3050
rect 5250 3040 6500 3050
rect 6650 3040 8300 3050
rect 0 3030 1200 3040
rect 1300 3030 2000 3040
rect 3200 3030 3700 3040
rect 5250 3030 6500 3040
rect 6650 3030 8300 3040
rect 0 3020 1200 3030
rect 1300 3020 2000 3030
rect 3200 3020 3700 3030
rect 5250 3020 6500 3030
rect 6650 3020 8300 3030
rect 0 3010 1200 3020
rect 1300 3010 2000 3020
rect 3200 3010 3700 3020
rect 5250 3010 6500 3020
rect 6650 3010 8300 3020
rect 0 3000 1200 3010
rect 1300 3000 2000 3010
rect 3200 3000 3700 3010
rect 5250 3000 6500 3010
rect 6650 3000 8300 3010
rect 0 2990 1150 3000
rect 1300 2990 1950 3000
rect 3200 2990 3750 3000
rect 5250 2990 6500 3000
rect 6650 2990 8250 3000
rect 0 2980 1150 2990
rect 1300 2980 1950 2990
rect 3200 2980 3750 2990
rect 5250 2980 6500 2990
rect 6650 2980 8250 2990
rect 0 2970 1150 2980
rect 1300 2970 1950 2980
rect 3200 2970 3750 2980
rect 5250 2970 6500 2980
rect 6650 2970 8250 2980
rect 0 2960 1150 2970
rect 1300 2960 1950 2970
rect 3200 2960 3750 2970
rect 5250 2960 6500 2970
rect 6650 2960 8250 2970
rect 0 2950 1150 2960
rect 1300 2950 1950 2960
rect 3200 2950 3750 2960
rect 5250 2950 6500 2960
rect 6650 2950 8250 2960
rect 0 2940 1150 2950
rect 1300 2940 1950 2950
rect 3200 2940 3800 2950
rect 5200 2940 6500 2950
rect 6600 2940 8250 2950
rect 0 2930 1150 2940
rect 1300 2930 1950 2940
rect 3200 2930 3800 2940
rect 5200 2930 6500 2940
rect 6600 2930 8250 2940
rect 0 2920 1150 2930
rect 1300 2920 1950 2930
rect 3200 2920 3800 2930
rect 5200 2920 6500 2930
rect 6600 2920 8250 2930
rect 0 2910 1150 2920
rect 1300 2910 1950 2920
rect 3200 2910 3800 2920
rect 5200 2910 6500 2920
rect 6600 2910 8250 2920
rect 0 2900 1150 2910
rect 1300 2900 1950 2910
rect 3200 2900 3800 2910
rect 5200 2900 6500 2910
rect 6600 2900 8250 2910
rect 0 2890 1150 2900
rect 1250 2890 1950 2900
rect 3200 2890 3850 2900
rect 4300 2890 4350 2900
rect 5200 2890 6500 2900
rect 6600 2890 7200 2900
rect 7550 2890 8200 2900
rect 0 2880 1150 2890
rect 1250 2880 1950 2890
rect 3200 2880 3850 2890
rect 4300 2880 4350 2890
rect 5200 2880 6500 2890
rect 6600 2880 7200 2890
rect 7550 2880 8200 2890
rect 0 2870 1150 2880
rect 1250 2870 1950 2880
rect 3200 2870 3850 2880
rect 4300 2870 4350 2880
rect 5200 2870 6500 2880
rect 6600 2870 7200 2880
rect 7550 2870 8200 2880
rect 0 2860 1150 2870
rect 1250 2860 1950 2870
rect 3200 2860 3850 2870
rect 4300 2860 4350 2870
rect 5200 2860 6500 2870
rect 6600 2860 7200 2870
rect 7550 2860 8200 2870
rect 0 2850 1150 2860
rect 1250 2850 1950 2860
rect 3200 2850 3850 2860
rect 4300 2850 4350 2860
rect 5200 2850 6500 2860
rect 6600 2850 7200 2860
rect 7550 2850 8200 2860
rect 0 2840 1100 2850
rect 1250 2840 1950 2850
rect 3200 2840 3900 2850
rect 4300 2840 4450 2850
rect 5200 2840 5850 2850
rect 6100 2840 6500 2850
rect 6600 2840 7100 2850
rect 7600 2840 8150 2850
rect 0 2830 1100 2840
rect 1250 2830 1950 2840
rect 3200 2830 3900 2840
rect 4300 2830 4450 2840
rect 5200 2830 5850 2840
rect 6100 2830 6500 2840
rect 6600 2830 7100 2840
rect 7600 2830 8150 2840
rect 0 2820 1100 2830
rect 1250 2820 1950 2830
rect 3200 2820 3900 2830
rect 4300 2820 4450 2830
rect 5200 2820 5850 2830
rect 6100 2820 6500 2830
rect 6600 2820 7100 2830
rect 7600 2820 8150 2830
rect 0 2810 1100 2820
rect 1250 2810 1950 2820
rect 3200 2810 3900 2820
rect 4300 2810 4450 2820
rect 5200 2810 5850 2820
rect 6100 2810 6500 2820
rect 6600 2810 7100 2820
rect 7600 2810 8150 2820
rect 0 2800 1100 2810
rect 1250 2800 1950 2810
rect 3200 2800 3900 2810
rect 4300 2800 4450 2810
rect 5200 2800 5850 2810
rect 6100 2800 6500 2810
rect 6600 2800 7100 2810
rect 7600 2800 8150 2810
rect 0 2790 1100 2800
rect 1200 2790 1950 2800
rect 3200 2790 3900 2800
rect 4300 2790 4500 2800
rect 5200 2790 5550 2800
rect 6150 2790 6500 2800
rect 6550 2790 7000 2800
rect 7700 2790 8100 2800
rect 0 2780 1100 2790
rect 1200 2780 1950 2790
rect 3200 2780 3900 2790
rect 4300 2780 4500 2790
rect 5200 2780 5550 2790
rect 6150 2780 6500 2790
rect 6550 2780 7000 2790
rect 7700 2780 8100 2790
rect 0 2770 1100 2780
rect 1200 2770 1950 2780
rect 3200 2770 3900 2780
rect 4300 2770 4500 2780
rect 5200 2770 5550 2780
rect 6150 2770 6500 2780
rect 6550 2770 7000 2780
rect 7700 2770 8100 2780
rect 0 2760 1100 2770
rect 1200 2760 1950 2770
rect 3200 2760 3900 2770
rect 4300 2760 4500 2770
rect 5200 2760 5550 2770
rect 6150 2760 6500 2770
rect 6550 2760 7000 2770
rect 7700 2760 8100 2770
rect 0 2750 1100 2760
rect 1200 2750 1950 2760
rect 3200 2750 3900 2760
rect 4300 2750 4500 2760
rect 5200 2750 5550 2760
rect 6150 2750 6500 2760
rect 6550 2750 7000 2760
rect 7700 2750 8100 2760
rect 0 2740 1050 2750
rect 1200 2740 1950 2750
rect 3200 2740 3850 2750
rect 4300 2740 4650 2750
rect 5200 2740 5250 2750
rect 5350 2740 5450 2750
rect 6200 2740 6500 2750
rect 6550 2740 6950 2750
rect 7700 2740 8050 2750
rect 0 2730 1050 2740
rect 1200 2730 1950 2740
rect 3200 2730 3850 2740
rect 4300 2730 4650 2740
rect 5200 2730 5250 2740
rect 5350 2730 5450 2740
rect 6200 2730 6500 2740
rect 6550 2730 6950 2740
rect 7700 2730 8050 2740
rect 0 2720 1050 2730
rect 1200 2720 1950 2730
rect 3200 2720 3850 2730
rect 4300 2720 4650 2730
rect 5200 2720 5250 2730
rect 5350 2720 5450 2730
rect 6200 2720 6500 2730
rect 6550 2720 6950 2730
rect 7700 2720 8050 2730
rect 0 2710 1050 2720
rect 1200 2710 1950 2720
rect 3200 2710 3850 2720
rect 4300 2710 4650 2720
rect 5200 2710 5250 2720
rect 5350 2710 5450 2720
rect 6200 2710 6500 2720
rect 6550 2710 6950 2720
rect 7700 2710 8050 2720
rect 0 2700 1050 2710
rect 1200 2700 1950 2710
rect 3200 2700 3850 2710
rect 4300 2700 4650 2710
rect 5200 2700 5250 2710
rect 5350 2700 5450 2710
rect 6200 2700 6500 2710
rect 6550 2700 6950 2710
rect 7700 2700 8050 2710
rect 0 2690 1050 2700
rect 1150 2690 1950 2700
rect 3200 2690 3850 2700
rect 4300 2690 4800 2700
rect 6250 2690 6500 2700
rect 6550 2690 6850 2700
rect 7750 2690 8000 2700
rect 0 2680 1050 2690
rect 1150 2680 1950 2690
rect 3200 2680 3850 2690
rect 4300 2680 4800 2690
rect 6250 2680 6500 2690
rect 6550 2680 6850 2690
rect 7750 2680 8000 2690
rect 0 2670 1050 2680
rect 1150 2670 1950 2680
rect 3200 2670 3850 2680
rect 4300 2670 4800 2680
rect 6250 2670 6500 2680
rect 6550 2670 6850 2680
rect 7750 2670 8000 2680
rect 0 2660 1050 2670
rect 1150 2660 1950 2670
rect 3200 2660 3850 2670
rect 4300 2660 4800 2670
rect 6250 2660 6500 2670
rect 6550 2660 6850 2670
rect 7750 2660 8000 2670
rect 0 2650 1050 2660
rect 1150 2650 1950 2660
rect 3200 2650 3850 2660
rect 4300 2650 4800 2660
rect 6250 2650 6500 2660
rect 6550 2650 6850 2660
rect 7750 2650 8000 2660
rect 0 2640 1000 2650
rect 1100 2640 1900 2650
rect 3150 2640 3850 2650
rect 4300 2640 4800 2650
rect 6300 2640 6850 2650
rect 7800 2640 7950 2650
rect 0 2630 1000 2640
rect 1100 2630 1900 2640
rect 3150 2630 3850 2640
rect 4300 2630 4800 2640
rect 6300 2630 6850 2640
rect 7800 2630 7950 2640
rect 0 2620 1000 2630
rect 1100 2620 1900 2630
rect 3150 2620 3850 2630
rect 4300 2620 4800 2630
rect 6300 2620 6850 2630
rect 7800 2620 7950 2630
rect 0 2610 1000 2620
rect 1100 2610 1900 2620
rect 3150 2610 3850 2620
rect 4300 2610 4800 2620
rect 6300 2610 6850 2620
rect 7800 2610 7950 2620
rect 0 2600 1000 2610
rect 1100 2600 1900 2610
rect 3150 2600 3850 2610
rect 4300 2600 4800 2610
rect 6300 2600 6850 2610
rect 7800 2600 7950 2610
rect 0 2590 1000 2600
rect 1100 2590 1900 2600
rect 2250 2590 2300 2600
rect 3150 2590 3850 2600
rect 4300 2590 4500 2600
rect 6300 2590 6800 2600
rect 7800 2590 7900 2600
rect 0 2580 1000 2590
rect 1100 2580 1900 2590
rect 2250 2580 2300 2590
rect 3150 2580 3850 2590
rect 4300 2580 4500 2590
rect 6300 2580 6800 2590
rect 7800 2580 7900 2590
rect 0 2570 1000 2580
rect 1100 2570 1900 2580
rect 2250 2570 2300 2580
rect 3150 2570 3850 2580
rect 4300 2570 4500 2580
rect 6300 2570 6800 2580
rect 7800 2570 7900 2580
rect 0 2560 1000 2570
rect 1100 2560 1900 2570
rect 2250 2560 2300 2570
rect 3150 2560 3850 2570
rect 4300 2560 4500 2570
rect 6300 2560 6800 2570
rect 7800 2560 7900 2570
rect 0 2550 1000 2560
rect 1100 2550 1900 2560
rect 2250 2550 2300 2560
rect 3150 2550 3850 2560
rect 4300 2550 4500 2560
rect 6300 2550 6800 2560
rect 7800 2550 7900 2560
rect 0 2540 950 2550
rect 1050 2540 1900 2550
rect 3250 2540 3900 2550
rect 4250 2540 4650 2550
rect 6350 2540 6750 2550
rect 0 2530 950 2540
rect 1050 2530 1900 2540
rect 3250 2530 3900 2540
rect 4250 2530 4650 2540
rect 6350 2530 6750 2540
rect 0 2520 950 2530
rect 1050 2520 1900 2530
rect 3250 2520 3900 2530
rect 4250 2520 4650 2530
rect 6350 2520 6750 2530
rect 0 2510 950 2520
rect 1050 2510 1900 2520
rect 3250 2510 3900 2520
rect 4250 2510 4650 2520
rect 6350 2510 6750 2520
rect 0 2500 950 2510
rect 1050 2500 1900 2510
rect 3250 2500 3900 2510
rect 4250 2500 4650 2510
rect 6350 2500 6750 2510
rect 0 2490 950 2500
rect 1050 2490 1850 2500
rect 3300 2490 3950 2500
rect 4150 2490 4600 2500
rect 6350 2490 6700 2500
rect 0 2480 950 2490
rect 1050 2480 1850 2490
rect 3300 2480 3950 2490
rect 4150 2480 4600 2490
rect 6350 2480 6700 2490
rect 0 2470 950 2480
rect 1050 2470 1850 2480
rect 3300 2470 3950 2480
rect 4150 2470 4600 2480
rect 6350 2470 6700 2480
rect 0 2460 950 2470
rect 1050 2460 1850 2470
rect 3300 2460 3950 2470
rect 4150 2460 4600 2470
rect 6350 2460 6700 2470
rect 0 2450 950 2460
rect 1050 2450 1850 2460
rect 3300 2450 3950 2460
rect 4150 2450 4600 2460
rect 6350 2450 6700 2460
rect 0 2440 900 2450
rect 1050 2440 1850 2450
rect 3300 2440 4000 2450
rect 4050 2440 4550 2450
rect 6400 2440 6700 2450
rect 0 2430 900 2440
rect 1050 2430 1850 2440
rect 3300 2430 4000 2440
rect 4050 2430 4550 2440
rect 6400 2430 6700 2440
rect 0 2420 900 2430
rect 1050 2420 1850 2430
rect 3300 2420 4000 2430
rect 4050 2420 4550 2430
rect 6400 2420 6700 2430
rect 0 2410 900 2420
rect 1050 2410 1850 2420
rect 3300 2410 4000 2420
rect 4050 2410 4550 2420
rect 6400 2410 6700 2420
rect 0 2400 900 2410
rect 1050 2400 1850 2410
rect 3300 2400 4000 2410
rect 4050 2400 4550 2410
rect 6400 2400 6700 2410
rect 0 2390 900 2400
rect 1050 2390 1850 2400
rect 3300 2390 4500 2400
rect 6400 2390 6700 2400
rect 0 2380 900 2390
rect 1050 2380 1850 2390
rect 3300 2380 4500 2390
rect 6400 2380 6700 2390
rect 0 2370 900 2380
rect 1050 2370 1850 2380
rect 3300 2370 4500 2380
rect 6400 2370 6700 2380
rect 0 2360 900 2370
rect 1050 2360 1850 2370
rect 3300 2360 4500 2370
rect 6400 2360 6700 2370
rect 0 2350 900 2360
rect 1050 2350 1850 2360
rect 3300 2350 4500 2360
rect 6400 2350 6700 2360
rect 0 2340 850 2350
rect 1000 2340 1850 2350
rect 3350 2340 4450 2350
rect 6450 2340 6700 2350
rect 0 2330 850 2340
rect 1000 2330 1850 2340
rect 3350 2330 4450 2340
rect 6450 2330 6700 2340
rect 0 2320 850 2330
rect 1000 2320 1850 2330
rect 3350 2320 4450 2330
rect 6450 2320 6700 2330
rect 0 2310 850 2320
rect 1000 2310 1850 2320
rect 3350 2310 4450 2320
rect 6450 2310 6700 2320
rect 0 2300 850 2310
rect 1000 2300 1850 2310
rect 3350 2300 4450 2310
rect 6450 2300 6700 2310
rect 0 2290 850 2300
rect 1000 2290 1800 2300
rect 3350 2290 4100 2300
rect 6500 2290 6700 2300
rect 8400 2290 8500 2300
rect 0 2280 850 2290
rect 1000 2280 1800 2290
rect 3350 2280 4100 2290
rect 6500 2280 6700 2290
rect 8400 2280 8500 2290
rect 0 2270 850 2280
rect 1000 2270 1800 2280
rect 3350 2270 4100 2280
rect 6500 2270 6700 2280
rect 8400 2270 8500 2280
rect 0 2260 850 2270
rect 1000 2260 1800 2270
rect 3350 2260 4100 2270
rect 6500 2260 6700 2270
rect 8400 2260 8500 2270
rect 0 2250 850 2260
rect 1000 2250 1800 2260
rect 3350 2250 4100 2260
rect 6500 2250 6700 2260
rect 8400 2250 8500 2260
rect 0 2240 800 2250
rect 1000 2240 1800 2250
rect 3350 2240 4350 2250
rect 6500 2240 6700 2250
rect 8400 2240 8600 2250
rect 9150 2240 9200 2250
rect 0 2230 800 2240
rect 1000 2230 1800 2240
rect 3350 2230 4350 2240
rect 6500 2230 6700 2240
rect 8400 2230 8600 2240
rect 9150 2230 9200 2240
rect 0 2220 800 2230
rect 1000 2220 1800 2230
rect 3350 2220 4350 2230
rect 6500 2220 6700 2230
rect 8400 2220 8600 2230
rect 9150 2220 9200 2230
rect 0 2210 800 2220
rect 1000 2210 1800 2220
rect 3350 2210 4350 2220
rect 6500 2210 6700 2220
rect 8400 2210 8600 2220
rect 9150 2210 9200 2220
rect 0 2200 800 2210
rect 1000 2200 1800 2210
rect 3350 2200 4350 2210
rect 6500 2200 6700 2210
rect 8400 2200 8600 2210
rect 9150 2200 9200 2210
rect 0 2190 800 2200
rect 1000 2190 1800 2200
rect 3350 2190 4350 2200
rect 6550 2190 6700 2200
rect 7100 2190 7250 2200
rect 7550 2190 7600 2200
rect 8400 2190 8800 2200
rect 9050 2190 9200 2200
rect 0 2180 800 2190
rect 1000 2180 1800 2190
rect 3350 2180 4350 2190
rect 6550 2180 6700 2190
rect 7100 2180 7250 2190
rect 7550 2180 7600 2190
rect 8400 2180 8800 2190
rect 9050 2180 9200 2190
rect 0 2170 800 2180
rect 1000 2170 1800 2180
rect 3350 2170 4350 2180
rect 6550 2170 6700 2180
rect 7100 2170 7250 2180
rect 7550 2170 7600 2180
rect 8400 2170 8800 2180
rect 9050 2170 9200 2180
rect 0 2160 800 2170
rect 1000 2160 1800 2170
rect 3350 2160 4350 2170
rect 6550 2160 6700 2170
rect 7100 2160 7250 2170
rect 7550 2160 7600 2170
rect 8400 2160 8800 2170
rect 9050 2160 9200 2170
rect 0 2150 800 2160
rect 1000 2150 1800 2160
rect 3350 2150 4350 2160
rect 6550 2150 6700 2160
rect 7100 2150 7250 2160
rect 7550 2150 7600 2160
rect 8400 2150 8800 2160
rect 9050 2150 9200 2160
rect 0 2140 750 2150
rect 1000 2140 1800 2150
rect 3350 2140 4350 2150
rect 6550 2140 6700 2150
rect 7500 2140 7700 2150
rect 8450 2140 9200 2150
rect 0 2130 750 2140
rect 1000 2130 1800 2140
rect 3350 2130 4350 2140
rect 6550 2130 6700 2140
rect 7500 2130 7700 2140
rect 8450 2130 9200 2140
rect 0 2120 750 2130
rect 1000 2120 1800 2130
rect 3350 2120 4350 2130
rect 6550 2120 6700 2130
rect 7500 2120 7700 2130
rect 8450 2120 9200 2130
rect 0 2110 750 2120
rect 1000 2110 1800 2120
rect 3350 2110 4350 2120
rect 6550 2110 6700 2120
rect 7500 2110 7700 2120
rect 8450 2110 9200 2120
rect 0 2100 750 2110
rect 1000 2100 1800 2110
rect 3350 2100 4350 2110
rect 6550 2100 6700 2110
rect 7500 2100 7700 2110
rect 8450 2100 9200 2110
rect 0 2090 750 2100
rect 950 2090 1800 2100
rect 3350 2090 4350 2100
rect 6550 2090 6750 2100
rect 7350 2090 7800 2100
rect 8550 2090 9100 2100
rect 0 2080 750 2090
rect 950 2080 1800 2090
rect 3350 2080 4350 2090
rect 6550 2080 6750 2090
rect 7350 2080 7800 2090
rect 8550 2080 9100 2090
rect 0 2070 750 2080
rect 950 2070 1800 2080
rect 3350 2070 4350 2080
rect 6550 2070 6750 2080
rect 7350 2070 7800 2080
rect 8550 2070 9100 2080
rect 0 2060 750 2070
rect 950 2060 1800 2070
rect 3350 2060 4350 2070
rect 6550 2060 6750 2070
rect 7350 2060 7800 2070
rect 8550 2060 9100 2070
rect 0 2050 750 2060
rect 950 2050 1800 2060
rect 3350 2050 4350 2060
rect 6550 2050 6750 2060
rect 7350 2050 7800 2060
rect 8550 2050 9100 2060
rect 0 2040 700 2050
rect 950 2040 1800 2050
rect 3350 2040 4350 2050
rect 6550 2040 6750 2050
rect 7350 2040 7750 2050
rect 8650 2040 9050 2050
rect 0 2030 700 2040
rect 950 2030 1800 2040
rect 3350 2030 4350 2040
rect 6550 2030 6750 2040
rect 7350 2030 7750 2040
rect 8650 2030 9050 2040
rect 0 2020 700 2030
rect 950 2020 1800 2030
rect 3350 2020 4350 2030
rect 6550 2020 6750 2030
rect 7350 2020 7750 2030
rect 8650 2020 9050 2030
rect 0 2010 700 2020
rect 950 2010 1800 2020
rect 3350 2010 4350 2020
rect 6550 2010 6750 2020
rect 7350 2010 7750 2020
rect 8650 2010 9050 2020
rect 0 2000 700 2010
rect 950 2000 1800 2010
rect 3350 2000 4350 2010
rect 6550 2000 6750 2010
rect 7350 2000 7750 2010
rect 8650 2000 9050 2010
rect 0 1990 700 2000
rect 950 1990 1800 2000
rect 3350 1990 4350 2000
rect 6550 1990 6750 2000
rect 7400 1990 7700 2000
rect 0 1980 700 1990
rect 950 1980 1800 1990
rect 3350 1980 4350 1990
rect 6550 1980 6750 1990
rect 7400 1980 7700 1990
rect 0 1970 700 1980
rect 950 1970 1800 1980
rect 3350 1970 4350 1980
rect 6550 1970 6750 1980
rect 7400 1970 7700 1980
rect 0 1960 700 1970
rect 950 1960 1800 1970
rect 3350 1960 4350 1970
rect 6550 1960 6750 1970
rect 7400 1960 7700 1970
rect 0 1950 700 1960
rect 950 1950 1800 1960
rect 3350 1950 4350 1960
rect 6550 1950 6750 1960
rect 7400 1950 7700 1960
rect 0 1940 650 1950
rect 950 1940 1800 1950
rect 3350 1940 4350 1950
rect 6600 1940 6750 1950
rect 7400 1940 7700 1950
rect 0 1930 650 1940
rect 950 1930 1800 1940
rect 3350 1930 4350 1940
rect 6600 1930 6750 1940
rect 7400 1930 7700 1940
rect 0 1920 650 1930
rect 950 1920 1800 1930
rect 3350 1920 4350 1930
rect 6600 1920 6750 1930
rect 7400 1920 7700 1930
rect 0 1910 650 1920
rect 950 1910 1800 1920
rect 3350 1910 4350 1920
rect 6600 1910 6750 1920
rect 7400 1910 7700 1920
rect 0 1900 650 1910
rect 950 1900 1800 1910
rect 3350 1900 4350 1910
rect 6600 1900 6750 1910
rect 7400 1900 7700 1910
rect 0 1890 650 1900
rect 950 1890 1800 1900
rect 3350 1890 4250 1900
rect 6600 1890 6750 1900
rect 7400 1890 7700 1900
rect 0 1880 650 1890
rect 950 1880 1800 1890
rect 3350 1880 4250 1890
rect 6600 1880 6750 1890
rect 7400 1880 7700 1890
rect 0 1870 650 1880
rect 950 1870 1800 1880
rect 3350 1870 4250 1880
rect 6600 1870 6750 1880
rect 7400 1870 7700 1880
rect 0 1860 650 1870
rect 950 1860 1800 1870
rect 3350 1860 4250 1870
rect 6600 1860 6750 1870
rect 7400 1860 7700 1870
rect 0 1850 650 1860
rect 950 1850 1800 1860
rect 3350 1850 4250 1860
rect 6600 1850 6750 1860
rect 7400 1850 7700 1860
rect 0 1840 600 1850
rect 900 1840 1800 1850
rect 3350 1840 4050 1850
rect 6600 1840 6750 1850
rect 7400 1840 7750 1850
rect 0 1830 600 1840
rect 900 1830 1800 1840
rect 3350 1830 4050 1840
rect 6600 1830 6750 1840
rect 7400 1830 7750 1840
rect 0 1820 600 1830
rect 900 1820 1800 1830
rect 3350 1820 4050 1830
rect 6600 1820 6750 1830
rect 7400 1820 7750 1830
rect 0 1810 600 1820
rect 900 1810 1800 1820
rect 3350 1810 4050 1820
rect 6600 1810 6750 1820
rect 7400 1810 7750 1820
rect 0 1800 600 1810
rect 900 1800 1800 1810
rect 3350 1800 4050 1810
rect 6600 1800 6750 1810
rect 7400 1800 7750 1810
rect 0 1790 600 1800
rect 900 1790 1800 1800
rect 3350 1790 4050 1800
rect 6650 1790 6750 1800
rect 7400 1790 7750 1800
rect 0 1780 600 1790
rect 900 1780 1800 1790
rect 3350 1780 4050 1790
rect 6650 1780 6750 1790
rect 7400 1780 7750 1790
rect 0 1770 600 1780
rect 900 1770 1800 1780
rect 3350 1770 4050 1780
rect 6650 1770 6750 1780
rect 7400 1770 7750 1780
rect 0 1760 600 1770
rect 900 1760 1800 1770
rect 3350 1760 4050 1770
rect 6650 1760 6750 1770
rect 7400 1760 7750 1770
rect 0 1750 600 1760
rect 900 1750 1800 1760
rect 3350 1750 4050 1760
rect 6650 1750 6750 1760
rect 7400 1750 7750 1760
rect 0 1740 550 1750
rect 900 1740 1850 1750
rect 3350 1740 4000 1750
rect 6650 1740 6750 1750
rect 7400 1740 7750 1750
rect 0 1730 550 1740
rect 900 1730 1850 1740
rect 3350 1730 4000 1740
rect 6650 1730 6750 1740
rect 7400 1730 7750 1740
rect 0 1720 550 1730
rect 900 1720 1850 1730
rect 3350 1720 4000 1730
rect 6650 1720 6750 1730
rect 7400 1720 7750 1730
rect 0 1710 550 1720
rect 900 1710 1850 1720
rect 3350 1710 4000 1720
rect 6650 1710 6750 1720
rect 7400 1710 7750 1720
rect 0 1700 550 1710
rect 900 1700 1850 1710
rect 3350 1700 4000 1710
rect 6650 1700 6750 1710
rect 7400 1700 7750 1710
rect 0 1690 550 1700
rect 900 1690 1850 1700
rect 3300 1690 4050 1700
rect 6650 1690 6750 1700
rect 7400 1690 7750 1700
rect 0 1680 550 1690
rect 900 1680 1850 1690
rect 3300 1680 4050 1690
rect 6650 1680 6750 1690
rect 7400 1680 7750 1690
rect 0 1670 550 1680
rect 900 1670 1850 1680
rect 3300 1670 4050 1680
rect 6650 1670 6750 1680
rect 7400 1670 7750 1680
rect 0 1660 550 1670
rect 900 1660 1850 1670
rect 3300 1660 4050 1670
rect 6650 1660 6750 1670
rect 7400 1660 7750 1670
rect 0 1650 550 1660
rect 900 1650 1850 1660
rect 3300 1650 4050 1660
rect 6650 1650 6750 1660
rect 7400 1650 7750 1660
rect 0 1640 550 1650
rect 900 1640 1900 1650
rect 3300 1640 4050 1650
rect 6200 1640 6250 1650
rect 6700 1640 6750 1650
rect 7400 1640 7750 1650
rect 0 1630 550 1640
rect 900 1630 1900 1640
rect 3300 1630 4050 1640
rect 6200 1630 6250 1640
rect 6700 1630 6750 1640
rect 7400 1630 7750 1640
rect 0 1620 550 1630
rect 900 1620 1900 1630
rect 3300 1620 4050 1630
rect 6200 1620 6250 1630
rect 6700 1620 6750 1630
rect 7400 1620 7750 1630
rect 0 1610 550 1620
rect 900 1610 1900 1620
rect 3300 1610 4050 1620
rect 6200 1610 6250 1620
rect 6700 1610 6750 1620
rect 7400 1610 7750 1620
rect 0 1600 550 1610
rect 900 1600 1900 1610
rect 3300 1600 4050 1610
rect 6200 1600 6250 1610
rect 6700 1600 6750 1610
rect 7400 1600 7750 1610
rect 0 1590 500 1600
rect 850 1590 1900 1600
rect 3250 1590 4050 1600
rect 7400 1590 7750 1600
rect 0 1580 500 1590
rect 850 1580 1900 1590
rect 3250 1580 4050 1590
rect 7400 1580 7750 1590
rect 0 1570 500 1580
rect 850 1570 1900 1580
rect 3250 1570 4050 1580
rect 7400 1570 7750 1580
rect 0 1560 500 1570
rect 850 1560 1900 1570
rect 3250 1560 4050 1570
rect 7400 1560 7750 1570
rect 0 1550 500 1560
rect 850 1550 1900 1560
rect 3250 1550 4050 1560
rect 7400 1550 7750 1560
rect 0 1540 500 1550
rect 850 1540 1950 1550
rect 3200 1540 4100 1550
rect 6250 1540 6300 1550
rect 7400 1540 7750 1550
rect 0 1530 500 1540
rect 850 1530 1950 1540
rect 3200 1530 4100 1540
rect 6250 1530 6300 1540
rect 7400 1530 7750 1540
rect 0 1520 500 1530
rect 850 1520 1950 1530
rect 3200 1520 4100 1530
rect 6250 1520 6300 1530
rect 7400 1520 7750 1530
rect 0 1510 500 1520
rect 850 1510 1950 1520
rect 3200 1510 4100 1520
rect 6250 1510 6300 1520
rect 7400 1510 7750 1520
rect 0 1500 500 1510
rect 850 1500 1950 1510
rect 3200 1500 4100 1510
rect 6250 1500 6300 1510
rect 7400 1500 7750 1510
rect 0 1490 500 1500
rect 1000 1490 1950 1500
rect 3150 1490 4100 1500
rect 6200 1490 6300 1500
rect 7400 1490 7800 1500
rect 0 1480 500 1490
rect 1000 1480 1950 1490
rect 3150 1480 4100 1490
rect 6200 1480 6300 1490
rect 7400 1480 7800 1490
rect 0 1470 500 1480
rect 1000 1470 1950 1480
rect 3150 1470 4100 1480
rect 6200 1470 6300 1480
rect 7400 1470 7800 1480
rect 0 1460 500 1470
rect 1000 1460 1950 1470
rect 3150 1460 4100 1470
rect 6200 1460 6300 1470
rect 7400 1460 7800 1470
rect 0 1450 500 1460
rect 1000 1450 1950 1460
rect 3150 1450 4100 1460
rect 6200 1450 6300 1460
rect 7400 1450 7800 1460
rect 0 1440 450 1450
rect 1050 1440 2000 1450
rect 3100 1440 4100 1450
rect 6200 1440 6300 1450
rect 7450 1440 7800 1450
rect 0 1430 450 1440
rect 1050 1430 2000 1440
rect 3100 1430 4100 1440
rect 6200 1430 6300 1440
rect 7450 1430 7800 1440
rect 0 1420 450 1430
rect 1050 1420 2000 1430
rect 3100 1420 4100 1430
rect 6200 1420 6300 1430
rect 7450 1420 7800 1430
rect 0 1410 450 1420
rect 1050 1410 2000 1420
rect 3100 1410 4100 1420
rect 6200 1410 6300 1420
rect 7450 1410 7800 1420
rect 0 1400 450 1410
rect 1050 1400 2000 1410
rect 3100 1400 4100 1410
rect 6200 1400 6300 1410
rect 7450 1400 7800 1410
rect 0 1390 450 1400
rect 1050 1390 2050 1400
rect 3050 1390 3500 1400
rect 3700 1390 4150 1400
rect 6200 1390 6300 1400
rect 7450 1390 7800 1400
rect 0 1380 450 1390
rect 1050 1380 2050 1390
rect 3050 1380 3500 1390
rect 3700 1380 4150 1390
rect 6200 1380 6300 1390
rect 7450 1380 7800 1390
rect 0 1370 450 1380
rect 1050 1370 2050 1380
rect 3050 1370 3500 1380
rect 3700 1370 4150 1380
rect 6200 1370 6300 1380
rect 7450 1370 7800 1380
rect 0 1360 450 1370
rect 1050 1360 2050 1370
rect 3050 1360 3500 1370
rect 3700 1360 4150 1370
rect 6200 1360 6300 1370
rect 7450 1360 7800 1370
rect 0 1350 450 1360
rect 1050 1350 2050 1360
rect 3050 1350 3500 1360
rect 3700 1350 4150 1360
rect 6200 1350 6300 1360
rect 7450 1350 7800 1360
rect 0 1340 450 1350
rect 1050 1340 2050 1350
rect 3000 1340 3450 1350
rect 3750 1340 4150 1350
rect 6200 1340 6300 1350
rect 7450 1340 7800 1350
rect 0 1330 450 1340
rect 1050 1330 2050 1340
rect 3000 1330 3450 1340
rect 3750 1330 4150 1340
rect 6200 1330 6300 1340
rect 7450 1330 7800 1340
rect 0 1320 450 1330
rect 1050 1320 2050 1330
rect 3000 1320 3450 1330
rect 3750 1320 4150 1330
rect 6200 1320 6300 1330
rect 7450 1320 7800 1330
rect 0 1310 450 1320
rect 1050 1310 2050 1320
rect 3000 1310 3450 1320
rect 3750 1310 4150 1320
rect 6200 1310 6300 1320
rect 7450 1310 7800 1320
rect 0 1300 450 1310
rect 1050 1300 2050 1310
rect 3000 1300 3450 1310
rect 3750 1300 4150 1310
rect 6200 1300 6300 1310
rect 7450 1300 7800 1310
rect 0 1290 400 1300
rect 1050 1290 2050 1300
rect 2900 1290 3450 1300
rect 3800 1290 4150 1300
rect 6250 1290 6300 1300
rect 7450 1290 7800 1300
rect 0 1280 400 1290
rect 1050 1280 2050 1290
rect 2900 1280 3450 1290
rect 3800 1280 4150 1290
rect 6250 1280 6300 1290
rect 7450 1280 7800 1290
rect 0 1270 400 1280
rect 1050 1270 2050 1280
rect 2900 1270 3450 1280
rect 3800 1270 4150 1280
rect 6250 1270 6300 1280
rect 7450 1270 7800 1280
rect 0 1260 400 1270
rect 1050 1260 2050 1270
rect 2900 1260 3450 1270
rect 3800 1260 4150 1270
rect 6250 1260 6300 1270
rect 7450 1260 7800 1270
rect 0 1250 400 1260
rect 1050 1250 2050 1260
rect 2900 1250 3450 1260
rect 3800 1250 4150 1260
rect 6250 1250 6300 1260
rect 7450 1250 7800 1260
rect 0 1240 400 1250
rect 1000 1240 2000 1250
rect 2800 1240 3450 1250
rect 3900 1240 4150 1250
rect 6250 1240 6300 1250
rect 7450 1240 7850 1250
rect 0 1230 400 1240
rect 1000 1230 2000 1240
rect 2800 1230 3450 1240
rect 3900 1230 4150 1240
rect 6250 1230 6300 1240
rect 7450 1230 7850 1240
rect 0 1220 400 1230
rect 1000 1220 2000 1230
rect 2800 1220 3450 1230
rect 3900 1220 4150 1230
rect 6250 1220 6300 1230
rect 7450 1220 7850 1230
rect 0 1210 400 1220
rect 1000 1210 2000 1220
rect 2800 1210 3450 1220
rect 3900 1210 4150 1220
rect 6250 1210 6300 1220
rect 7450 1210 7850 1220
rect 0 1200 400 1210
rect 1000 1200 2000 1210
rect 2800 1200 3450 1210
rect 3900 1200 4150 1210
rect 6250 1200 6300 1210
rect 7450 1200 7850 1210
rect 0 1190 400 1200
rect 1000 1190 2000 1200
rect 2850 1190 3500 1200
rect 3950 1190 4150 1200
rect 6250 1190 6350 1200
rect 7450 1190 7850 1200
rect 0 1180 400 1190
rect 1000 1180 2000 1190
rect 2850 1180 3500 1190
rect 3950 1180 4150 1190
rect 6250 1180 6350 1190
rect 7450 1180 7850 1190
rect 0 1170 400 1180
rect 1000 1170 2000 1180
rect 2850 1170 3500 1180
rect 3950 1170 4150 1180
rect 6250 1170 6350 1180
rect 7450 1170 7850 1180
rect 0 1160 400 1170
rect 1000 1160 2000 1170
rect 2850 1160 3500 1170
rect 3950 1160 4150 1170
rect 6250 1160 6350 1170
rect 7450 1160 7850 1170
rect 0 1150 400 1160
rect 1000 1150 2000 1160
rect 2850 1150 3500 1160
rect 3950 1150 4150 1160
rect 6250 1150 6350 1160
rect 7450 1150 7850 1160
rect 0 1140 350 1150
rect 650 1140 700 1150
rect 1000 1140 1500 1150
rect 1650 1140 2000 1150
rect 2900 1140 3550 1150
rect 4000 1140 4150 1150
rect 6300 1140 6400 1150
rect 7450 1140 7850 1150
rect 0 1130 350 1140
rect 650 1130 700 1140
rect 1000 1130 1500 1140
rect 1650 1130 2000 1140
rect 2900 1130 3550 1140
rect 4000 1130 4150 1140
rect 6300 1130 6400 1140
rect 7450 1130 7850 1140
rect 0 1120 350 1130
rect 650 1120 700 1130
rect 1000 1120 1500 1130
rect 1650 1120 2000 1130
rect 2900 1120 3550 1130
rect 4000 1120 4150 1130
rect 6300 1120 6400 1130
rect 7450 1120 7850 1130
rect 0 1110 350 1120
rect 650 1110 700 1120
rect 1000 1110 1500 1120
rect 1650 1110 2000 1120
rect 2900 1110 3550 1120
rect 4000 1110 4150 1120
rect 6300 1110 6400 1120
rect 7450 1110 7850 1120
rect 0 1100 350 1110
rect 650 1100 700 1110
rect 1000 1100 1500 1110
rect 1650 1100 2000 1110
rect 2900 1100 3550 1110
rect 4000 1100 4150 1110
rect 6300 1100 6400 1110
rect 7450 1100 7850 1110
rect 0 1090 350 1100
rect 650 1090 700 1100
rect 1000 1090 1450 1100
rect 1700 1090 1950 1100
rect 2900 1090 3600 1100
rect 4100 1090 4150 1100
rect 6300 1090 6400 1100
rect 7450 1090 7850 1100
rect 0 1080 350 1090
rect 650 1080 700 1090
rect 1000 1080 1450 1090
rect 1700 1080 1950 1090
rect 2900 1080 3600 1090
rect 4100 1080 4150 1090
rect 6300 1080 6400 1090
rect 7450 1080 7850 1090
rect 0 1070 350 1080
rect 650 1070 700 1080
rect 1000 1070 1450 1080
rect 1700 1070 1950 1080
rect 2900 1070 3600 1080
rect 4100 1070 4150 1080
rect 6300 1070 6400 1080
rect 7450 1070 7850 1080
rect 0 1060 350 1070
rect 650 1060 700 1070
rect 1000 1060 1450 1070
rect 1700 1060 1950 1070
rect 2900 1060 3600 1070
rect 4100 1060 4150 1070
rect 6300 1060 6400 1070
rect 7450 1060 7850 1070
rect 0 1050 350 1060
rect 650 1050 700 1060
rect 1000 1050 1450 1060
rect 1700 1050 1950 1060
rect 2900 1050 3600 1060
rect 4100 1050 4150 1060
rect 6300 1050 6400 1060
rect 7450 1050 7850 1060
rect 0 1040 300 1050
rect 1000 1040 1400 1050
rect 1700 1040 1950 1050
rect 2900 1040 3650 1050
rect 6300 1040 6350 1050
rect 7450 1040 7900 1050
rect 0 1030 300 1040
rect 1000 1030 1400 1040
rect 1700 1030 1950 1040
rect 2900 1030 3650 1040
rect 6300 1030 6350 1040
rect 7450 1030 7900 1040
rect 0 1020 300 1030
rect 1000 1020 1400 1030
rect 1700 1020 1950 1030
rect 2900 1020 3650 1030
rect 6300 1020 6350 1030
rect 7450 1020 7900 1030
rect 0 1010 300 1020
rect 1000 1010 1400 1020
rect 1700 1010 1950 1020
rect 2900 1010 3650 1020
rect 6300 1010 6350 1020
rect 7450 1010 7900 1020
rect 0 1000 300 1010
rect 1000 1000 1400 1010
rect 1700 1000 1950 1010
rect 2900 1000 3650 1010
rect 6300 1000 6350 1010
rect 7450 1000 7900 1010
rect 0 990 300 1000
rect 950 990 1350 1000
rect 1650 990 1950 1000
rect 2900 990 3700 1000
rect 7450 990 7900 1000
rect 0 980 300 990
rect 950 980 1350 990
rect 1650 980 1950 990
rect 2900 980 3700 990
rect 7450 980 7900 990
rect 0 970 300 980
rect 950 970 1350 980
rect 1650 970 1950 980
rect 2900 970 3700 980
rect 7450 970 7900 980
rect 0 960 300 970
rect 950 960 1350 970
rect 1650 960 1950 970
rect 2900 960 3700 970
rect 7450 960 7900 970
rect 0 950 300 960
rect 950 950 1350 960
rect 1650 950 1950 960
rect 2900 950 3700 960
rect 7450 950 7900 960
rect 0 940 250 950
rect 950 940 1250 950
rect 1600 940 1950 950
rect 2850 940 3750 950
rect 7450 940 7900 950
rect 0 930 250 940
rect 950 930 1250 940
rect 1600 930 1950 940
rect 2850 930 3750 940
rect 7450 930 7900 940
rect 0 920 250 930
rect 950 920 1250 930
rect 1600 920 1950 930
rect 2850 920 3750 930
rect 7450 920 7900 930
rect 0 910 250 920
rect 950 910 1250 920
rect 1600 910 1950 920
rect 2850 910 3750 920
rect 7450 910 7900 920
rect 0 900 250 910
rect 950 900 1250 910
rect 1600 900 1950 910
rect 2850 900 3750 910
rect 7450 900 7900 910
rect 0 890 250 900
rect 950 890 1200 900
rect 1550 890 1950 900
rect 2800 890 3800 900
rect 4900 890 5100 900
rect 5150 890 5200 900
rect 6300 890 6350 900
rect 7450 890 7900 900
rect 0 880 250 890
rect 950 880 1200 890
rect 1550 880 1950 890
rect 2800 880 3800 890
rect 4900 880 5100 890
rect 5150 880 5200 890
rect 6300 880 6350 890
rect 7450 880 7900 890
rect 0 870 250 880
rect 950 870 1200 880
rect 1550 870 1950 880
rect 2800 870 3800 880
rect 4900 870 5100 880
rect 5150 870 5200 880
rect 6300 870 6350 880
rect 7450 870 7900 880
rect 0 860 250 870
rect 950 860 1200 870
rect 1550 860 1950 870
rect 2800 860 3800 870
rect 4900 860 5100 870
rect 5150 860 5200 870
rect 6300 860 6350 870
rect 7450 860 7900 870
rect 0 850 250 860
rect 950 850 1200 860
rect 1550 850 1950 860
rect 2800 850 3800 860
rect 4900 850 5100 860
rect 5150 850 5200 860
rect 6300 850 6350 860
rect 7450 850 7900 860
rect 0 840 200 850
rect 950 840 1150 850
rect 1500 840 2000 850
rect 2700 840 3800 850
rect 4950 840 5200 850
rect 6350 840 6400 850
rect 7450 840 7900 850
rect 0 830 200 840
rect 950 830 1150 840
rect 1500 830 2000 840
rect 2700 830 3800 840
rect 4950 830 5200 840
rect 6350 830 6400 840
rect 7450 830 7900 840
rect 0 820 200 830
rect 950 820 1150 830
rect 1500 820 2000 830
rect 2700 820 3800 830
rect 4950 820 5200 830
rect 6350 820 6400 830
rect 7450 820 7900 830
rect 0 810 200 820
rect 950 810 1150 820
rect 1500 810 2000 820
rect 2700 810 3800 820
rect 4950 810 5200 820
rect 6350 810 6400 820
rect 7450 810 7900 820
rect 0 800 200 810
rect 950 800 1150 810
rect 1500 800 2000 810
rect 2700 800 3800 810
rect 4950 800 5200 810
rect 6350 800 6400 810
rect 7450 800 7900 810
rect 0 790 150 800
rect 950 790 1050 800
rect 1500 790 2000 800
rect 2650 790 3400 800
rect 4950 790 5200 800
rect 6350 790 6400 800
rect 7450 790 7950 800
rect 0 780 150 790
rect 950 780 1050 790
rect 1500 780 2000 790
rect 2650 780 3400 790
rect 4950 780 5200 790
rect 6350 780 6400 790
rect 7450 780 7950 790
rect 0 770 150 780
rect 950 770 1050 780
rect 1500 770 2000 780
rect 2650 770 3400 780
rect 4950 770 5200 780
rect 6350 770 6400 780
rect 7450 770 7950 780
rect 0 760 150 770
rect 950 760 1050 770
rect 1500 760 2000 770
rect 2650 760 3400 770
rect 4950 760 5200 770
rect 6350 760 6400 770
rect 7450 760 7950 770
rect 0 750 150 760
rect 950 750 1050 760
rect 1500 750 2000 760
rect 2650 750 3400 760
rect 4950 750 5200 760
rect 6350 750 6400 760
rect 7450 750 7950 760
rect 0 740 100 750
rect 900 740 1000 750
rect 1450 740 2050 750
rect 2550 740 3300 750
rect 4950 740 5150 750
rect 5200 740 5400 750
rect 6350 740 6400 750
rect 7450 740 7950 750
rect 0 730 100 740
rect 900 730 1000 740
rect 1450 730 2050 740
rect 2550 730 3300 740
rect 4950 730 5150 740
rect 5200 730 5400 740
rect 6350 730 6400 740
rect 7450 730 7950 740
rect 0 720 100 730
rect 900 720 1000 730
rect 1450 720 2050 730
rect 2550 720 3300 730
rect 4950 720 5150 730
rect 5200 720 5400 730
rect 6350 720 6400 730
rect 7450 720 7950 730
rect 0 710 100 720
rect 900 710 1000 720
rect 1450 710 2050 720
rect 2550 710 3300 720
rect 4950 710 5150 720
rect 5200 710 5400 720
rect 6350 710 6400 720
rect 7450 710 7950 720
rect 0 700 100 710
rect 900 700 1000 710
rect 1450 700 2050 710
rect 2550 700 3300 710
rect 4950 700 5150 710
rect 5200 700 5400 710
rect 6350 700 6400 710
rect 7450 700 7950 710
rect 1400 690 2050 700
rect 2450 690 3200 700
rect 5000 690 5150 700
rect 5200 690 5400 700
rect 6350 690 6450 700
rect 7450 690 7950 700
rect 1400 680 2050 690
rect 2450 680 3200 690
rect 5000 680 5150 690
rect 5200 680 5400 690
rect 6350 680 6450 690
rect 7450 680 7950 690
rect 1400 670 2050 680
rect 2450 670 3200 680
rect 5000 670 5150 680
rect 5200 670 5400 680
rect 6350 670 6450 680
rect 7450 670 7950 680
rect 1400 660 2050 670
rect 2450 660 3200 670
rect 5000 660 5150 670
rect 5200 660 5400 670
rect 6350 660 6450 670
rect 7450 660 7950 670
rect 1400 650 2050 660
rect 2450 650 3200 660
rect 5000 650 5150 660
rect 5200 650 5400 660
rect 6350 650 6450 660
rect 7450 650 7950 660
rect 1450 640 2050 650
rect 2350 640 3050 650
rect 5000 640 5400 650
rect 5450 640 5500 650
rect 6350 640 6500 650
rect 7450 640 8000 650
rect 1450 630 2050 640
rect 2350 630 3050 640
rect 5000 630 5400 640
rect 5450 630 5500 640
rect 6350 630 6500 640
rect 7450 630 8000 640
rect 1450 620 2050 630
rect 2350 620 3050 630
rect 5000 620 5400 630
rect 5450 620 5500 630
rect 6350 620 6500 630
rect 7450 620 8000 630
rect 1450 610 2050 620
rect 2350 610 3050 620
rect 5000 610 5400 620
rect 5450 610 5500 620
rect 6350 610 6500 620
rect 7450 610 8000 620
rect 1450 600 2050 610
rect 2350 600 3050 610
rect 5000 600 5400 610
rect 5450 600 5500 610
rect 6350 600 6500 610
rect 7450 600 8000 610
rect 1500 590 2100 600
rect 2300 590 2950 600
rect 5000 590 5550 600
rect 6350 590 6500 600
rect 7450 590 8000 600
rect 1500 580 2100 590
rect 2300 580 2950 590
rect 5000 580 5550 590
rect 6350 580 6500 590
rect 7450 580 8000 590
rect 1500 570 2100 580
rect 2300 570 2950 580
rect 5000 570 5550 580
rect 6350 570 6500 580
rect 7450 570 8000 580
rect 1500 560 2100 570
rect 2300 560 2950 570
rect 5000 560 5550 570
rect 6350 560 6500 570
rect 7450 560 8000 570
rect 1500 550 2100 560
rect 2300 550 2950 560
rect 5000 550 5550 560
rect 6350 550 6500 560
rect 7450 550 8000 560
rect 1550 540 2150 550
rect 2200 540 2800 550
rect 5000 540 5400 550
rect 5500 540 5600 550
rect 6350 540 6550 550
rect 7450 540 8050 550
rect 1550 530 2150 540
rect 2200 530 2800 540
rect 5000 530 5400 540
rect 5500 530 5600 540
rect 6350 530 6550 540
rect 7450 530 8050 540
rect 1550 520 2150 530
rect 2200 520 2800 530
rect 5000 520 5400 530
rect 5500 520 5600 530
rect 6350 520 6550 530
rect 7450 520 8050 530
rect 1550 510 2150 520
rect 2200 510 2800 520
rect 5000 510 5400 520
rect 5500 510 5600 520
rect 6350 510 6550 520
rect 7450 510 8050 520
rect 1550 500 2150 510
rect 2200 500 2800 510
rect 5000 500 5400 510
rect 5500 500 5600 510
rect 6350 500 6550 510
rect 7450 500 8050 510
rect 1750 490 1800 500
rect 2350 490 2550 500
rect 5000 490 5400 500
rect 5450 490 5650 500
rect 6350 490 6550 500
rect 7450 490 8100 500
rect 1750 480 1800 490
rect 2350 480 2550 490
rect 5000 480 5400 490
rect 5450 480 5650 490
rect 6350 480 6550 490
rect 7450 480 8100 490
rect 1750 470 1800 480
rect 2350 470 2550 480
rect 5000 470 5400 480
rect 5450 470 5650 480
rect 6350 470 6550 480
rect 7450 470 8100 480
rect 1750 460 1800 470
rect 2350 460 2550 470
rect 5000 460 5400 470
rect 5450 460 5650 470
rect 6350 460 6550 470
rect 7450 460 8100 470
rect 1750 450 1800 460
rect 2350 450 2550 460
rect 5000 450 5400 460
rect 5450 450 5650 460
rect 6350 450 6550 460
rect 7450 450 8100 460
rect 700 440 750 450
rect 5000 440 5700 450
rect 6350 440 6600 450
rect 7450 440 8200 450
rect 700 430 750 440
rect 5000 430 5700 440
rect 6350 430 6600 440
rect 7450 430 8200 440
rect 700 420 750 430
rect 5000 420 5700 430
rect 6350 420 6600 430
rect 7450 420 8200 430
rect 700 410 750 420
rect 5000 410 5700 420
rect 6350 410 6600 420
rect 7450 410 8200 420
rect 700 400 750 410
rect 5000 400 5700 410
rect 6350 400 6600 410
rect 7450 400 8200 410
rect 5000 390 5200 400
rect 5250 390 5300 400
rect 5400 390 5750 400
rect 6350 390 6600 400
rect 7450 390 8250 400
rect 5000 380 5200 390
rect 5250 380 5300 390
rect 5400 380 5750 390
rect 6350 380 6600 390
rect 7450 380 8250 390
rect 5000 370 5200 380
rect 5250 370 5300 380
rect 5400 370 5750 380
rect 6350 370 6600 380
rect 7450 370 8250 380
rect 5000 360 5200 370
rect 5250 360 5300 370
rect 5400 360 5750 370
rect 6350 360 6600 370
rect 7450 360 8250 370
rect 5000 350 5200 360
rect 5250 350 5300 360
rect 5400 350 5750 360
rect 6350 350 6600 360
rect 7450 350 8250 360
rect 5050 340 5700 350
rect 6350 340 6650 350
rect 7450 340 8300 350
rect 5050 330 5700 340
rect 6350 330 6650 340
rect 7450 330 8300 340
rect 5050 320 5700 330
rect 6350 320 6650 330
rect 7450 320 8300 330
rect 5050 310 5700 320
rect 6350 310 6650 320
rect 7450 310 8300 320
rect 5050 300 5700 310
rect 6350 300 6650 310
rect 7450 300 8300 310
rect 5050 290 5700 300
rect 6350 290 6700 300
rect 7450 290 8350 300
rect 5050 280 5700 290
rect 6350 280 6700 290
rect 7450 280 8350 290
rect 5050 270 5700 280
rect 6350 270 6700 280
rect 7450 270 8350 280
rect 5050 260 5700 270
rect 6350 260 6700 270
rect 7450 260 8350 270
rect 5050 250 5700 260
rect 6350 250 6700 260
rect 7450 250 8350 260
rect 5050 240 5950 250
rect 6400 240 6750 250
rect 7400 240 8400 250
rect 5050 230 5950 240
rect 6400 230 6750 240
rect 7400 230 8400 240
rect 5050 220 5950 230
rect 6400 220 6750 230
rect 7400 220 8400 230
rect 5050 210 5950 220
rect 6400 210 6750 220
rect 7400 210 8400 220
rect 5050 200 5950 210
rect 6400 200 6750 210
rect 7400 200 8400 210
rect 5050 190 5350 200
rect 5700 190 5950 200
rect 6400 190 6800 200
rect 7400 190 8450 200
rect 5050 180 5350 190
rect 5700 180 5950 190
rect 6400 180 6800 190
rect 7400 180 8450 190
rect 5050 170 5350 180
rect 5700 170 5950 180
rect 6400 170 6800 180
rect 7400 170 8450 180
rect 5050 160 5350 170
rect 5700 160 5950 170
rect 6400 160 6800 170
rect 7400 160 8450 170
rect 5050 150 5350 160
rect 5700 150 5950 160
rect 6400 150 6800 160
rect 7400 150 8450 160
rect 5100 140 5350 150
rect 6450 140 6800 150
rect 7400 140 8500 150
rect 5100 130 5350 140
rect 6450 130 6800 140
rect 7400 130 8500 140
rect 5100 120 5350 130
rect 6450 120 6800 130
rect 7400 120 8500 130
rect 5100 110 5350 120
rect 6450 110 6800 120
rect 7400 110 8500 120
rect 5100 100 5350 110
rect 6450 100 6800 110
rect 7400 100 8500 110
rect 400 90 500 100
rect 5100 90 5350 100
rect 6450 90 6800 100
rect 7400 90 8550 100
rect 400 80 500 90
rect 5100 80 5350 90
rect 6450 80 6800 90
rect 7400 80 8550 90
rect 400 70 500 80
rect 5100 70 5350 80
rect 6450 70 6800 80
rect 7400 70 8550 80
rect 400 60 500 70
rect 5100 60 5350 70
rect 6450 60 6800 70
rect 7400 60 8550 70
rect 400 50 500 60
rect 5100 50 5350 60
rect 6450 50 6800 60
rect 7400 50 8550 60
rect 350 40 600 50
rect 5100 40 5350 50
rect 5700 40 5800 50
rect 6500 40 6850 50
rect 7400 40 8550 50
rect 9250 40 9350 50
rect 350 30 600 40
rect 5100 30 5350 40
rect 5700 30 5800 40
rect 6500 30 6850 40
rect 7400 30 8550 40
rect 9250 30 9350 40
rect 350 20 600 30
rect 5100 20 5350 30
rect 5700 20 5800 30
rect 6500 20 6850 30
rect 7400 20 8550 30
rect 9250 20 9350 30
rect 350 10 600 20
rect 5100 10 5350 20
rect 5700 10 5800 20
rect 6500 10 6850 20
rect 7400 10 8550 20
rect 9250 10 9350 20
rect 350 0 600 10
rect 5100 0 5350 10
rect 5700 0 5800 10
rect 6500 0 6850 10
rect 7400 0 8550 10
rect 9250 0 9350 10
<< metal1 >>
rect 2200 7490 2250 7500
rect 3600 7490 3650 7500
rect 9800 7490 9990 7500
rect 2200 7480 2250 7490
rect 3600 7480 3650 7490
rect 9800 7480 9990 7490
rect 2200 7470 2250 7480
rect 3600 7470 3650 7480
rect 9800 7470 9990 7480
rect 2200 7460 2250 7470
rect 3600 7460 3650 7470
rect 9800 7460 9990 7470
rect 2200 7450 2250 7460
rect 3600 7450 3650 7460
rect 9800 7450 9990 7460
rect 2150 7440 2200 7450
rect 9750 7440 9950 7450
rect 2150 7430 2200 7440
rect 9750 7430 9950 7440
rect 2150 7420 2200 7430
rect 9750 7420 9950 7430
rect 2150 7410 2200 7420
rect 9750 7410 9950 7420
rect 2150 7400 2200 7410
rect 9750 7400 9950 7410
rect 2100 7390 2150 7400
rect 9650 7390 9950 7400
rect 2100 7380 2150 7390
rect 9650 7380 9950 7390
rect 2100 7370 2150 7380
rect 9650 7370 9950 7380
rect 2100 7360 2150 7370
rect 9650 7360 9950 7370
rect 2100 7350 2150 7360
rect 9650 7350 9950 7360
rect 3300 7340 3350 7350
rect 9750 7340 9800 7350
rect 9900 7340 9950 7350
rect 3300 7330 3350 7340
rect 9750 7330 9800 7340
rect 9900 7330 9950 7340
rect 3300 7320 3350 7330
rect 9750 7320 9800 7330
rect 9900 7320 9950 7330
rect 3300 7310 3350 7320
rect 9750 7310 9800 7320
rect 9900 7310 9950 7320
rect 3300 7300 3350 7310
rect 9750 7300 9800 7310
rect 9900 7300 9950 7310
rect 2050 7290 2100 7300
rect 2500 7290 2550 7300
rect 3300 7290 3350 7300
rect 2050 7280 2100 7290
rect 2500 7280 2550 7290
rect 3300 7280 3350 7290
rect 2050 7270 2100 7280
rect 2500 7270 2550 7280
rect 3300 7270 3350 7280
rect 2050 7260 2100 7270
rect 2500 7260 2550 7270
rect 3300 7260 3350 7270
rect 2050 7250 2100 7260
rect 2500 7250 2550 7260
rect 3300 7250 3350 7260
rect 2000 7240 2050 7250
rect 2400 7240 2450 7250
rect 2500 7240 2550 7250
rect 3300 7240 3350 7250
rect 9900 7240 9950 7250
rect 2000 7230 2050 7240
rect 2400 7230 2450 7240
rect 2500 7230 2550 7240
rect 3300 7230 3350 7240
rect 9900 7230 9950 7240
rect 2000 7220 2050 7230
rect 2400 7220 2450 7230
rect 2500 7220 2550 7230
rect 3300 7220 3350 7230
rect 9900 7220 9950 7230
rect 2000 7210 2050 7220
rect 2400 7210 2450 7220
rect 2500 7210 2550 7220
rect 3300 7210 3350 7220
rect 9900 7210 9950 7220
rect 2000 7200 2050 7210
rect 2400 7200 2450 7210
rect 2500 7200 2550 7210
rect 3300 7200 3350 7210
rect 9900 7200 9950 7210
rect 2000 7190 2050 7200
rect 2100 7190 2300 7200
rect 3300 7190 3350 7200
rect 9850 7190 9950 7200
rect 2000 7180 2050 7190
rect 2100 7180 2300 7190
rect 3300 7180 3350 7190
rect 9850 7180 9950 7190
rect 2000 7170 2050 7180
rect 2100 7170 2300 7180
rect 3300 7170 3350 7180
rect 9850 7170 9950 7180
rect 2000 7160 2050 7170
rect 2100 7160 2300 7170
rect 3300 7160 3350 7170
rect 9850 7160 9950 7170
rect 2000 7150 2050 7160
rect 2100 7150 2300 7160
rect 3300 7150 3350 7160
rect 9850 7150 9950 7160
rect 1950 7140 2250 7150
rect 3300 7140 3350 7150
rect 9850 7140 9990 7150
rect 1950 7130 2250 7140
rect 3300 7130 3350 7140
rect 9850 7130 9990 7140
rect 1950 7120 2250 7130
rect 3300 7120 3350 7130
rect 9850 7120 9990 7130
rect 1950 7110 2250 7120
rect 3300 7110 3350 7120
rect 9850 7110 9990 7120
rect 1950 7100 2250 7110
rect 3300 7100 3350 7110
rect 9850 7100 9990 7110
rect 2100 7090 2150 7100
rect 2250 7090 2400 7100
rect 3400 7090 3450 7100
rect 9800 7090 9850 7100
rect 9950 7090 9990 7100
rect 2100 7080 2150 7090
rect 2250 7080 2400 7090
rect 3400 7080 3450 7090
rect 9800 7080 9850 7090
rect 9950 7080 9990 7090
rect 2100 7070 2150 7080
rect 2250 7070 2400 7080
rect 3400 7070 3450 7080
rect 9800 7070 9850 7080
rect 9950 7070 9990 7080
rect 2100 7060 2150 7070
rect 2250 7060 2400 7070
rect 3400 7060 3450 7070
rect 9800 7060 9850 7070
rect 9950 7060 9990 7070
rect 2100 7050 2150 7060
rect 2250 7050 2400 7060
rect 3400 7050 3450 7060
rect 9800 7050 9850 7060
rect 9950 7050 9990 7060
rect 2200 7040 2250 7050
rect 2400 7040 2850 7050
rect 2900 7040 3000 7050
rect 3100 7040 3250 7050
rect 3450 7040 3500 7050
rect 9700 7040 9850 7050
rect 9900 7040 9990 7050
rect 2200 7030 2250 7040
rect 2400 7030 2850 7040
rect 2900 7030 3000 7040
rect 3100 7030 3250 7040
rect 3450 7030 3500 7040
rect 9700 7030 9850 7040
rect 9900 7030 9990 7040
rect 2200 7020 2250 7030
rect 2400 7020 2850 7030
rect 2900 7020 3000 7030
rect 3100 7020 3250 7030
rect 3450 7020 3500 7030
rect 9700 7020 9850 7030
rect 9900 7020 9990 7030
rect 2200 7010 2250 7020
rect 2400 7010 2850 7020
rect 2900 7010 3000 7020
rect 3100 7010 3250 7020
rect 3450 7010 3500 7020
rect 9700 7010 9850 7020
rect 9900 7010 9990 7020
rect 2200 7000 2250 7010
rect 2400 7000 2850 7010
rect 2900 7000 3000 7010
rect 3100 7000 3250 7010
rect 3450 7000 3500 7010
rect 9700 7000 9850 7010
rect 9900 7000 9990 7010
rect 2000 6990 2050 7000
rect 2150 6990 2250 7000
rect 3350 6990 3400 7000
rect 3500 6990 3550 7000
rect 9650 6990 9900 7000
rect 2000 6980 2050 6990
rect 2150 6980 2250 6990
rect 3350 6980 3400 6990
rect 3500 6980 3550 6990
rect 9650 6980 9900 6990
rect 2000 6970 2050 6980
rect 2150 6970 2250 6980
rect 3350 6970 3400 6980
rect 3500 6970 3550 6980
rect 9650 6970 9900 6980
rect 2000 6960 2050 6970
rect 2150 6960 2250 6970
rect 3350 6960 3400 6970
rect 3500 6960 3550 6970
rect 9650 6960 9900 6970
rect 2000 6950 2050 6960
rect 2150 6950 2250 6960
rect 3350 6950 3400 6960
rect 3500 6950 3550 6960
rect 9650 6950 9900 6960
rect 1950 6940 2000 6950
rect 2200 6940 2300 6950
rect 3500 6940 3650 6950
rect 9700 6940 9850 6950
rect 1950 6930 2000 6940
rect 2200 6930 2300 6940
rect 3500 6930 3650 6940
rect 9700 6930 9850 6940
rect 1950 6920 2000 6930
rect 2200 6920 2300 6930
rect 3500 6920 3650 6930
rect 9700 6920 9850 6930
rect 1950 6910 2000 6920
rect 2200 6910 2300 6920
rect 3500 6910 3650 6920
rect 9700 6910 9850 6920
rect 1950 6900 2000 6910
rect 2200 6900 2300 6910
rect 3500 6900 3650 6910
rect 9700 6900 9850 6910
rect 2250 6890 2350 6900
rect 3600 6890 3750 6900
rect 9700 6890 9850 6900
rect 2250 6880 2350 6890
rect 3600 6880 3750 6890
rect 9700 6880 9850 6890
rect 2250 6870 2350 6880
rect 3600 6870 3750 6880
rect 9700 6870 9850 6880
rect 2250 6860 2350 6870
rect 3600 6860 3750 6870
rect 9700 6860 9850 6870
rect 2250 6850 2350 6860
rect 3600 6850 3750 6860
rect 9700 6850 9850 6860
rect 1900 6840 2000 6850
rect 2300 6840 2450 6850
rect 3650 6840 3800 6850
rect 9700 6840 9990 6850
rect 1900 6830 2000 6840
rect 2300 6830 2450 6840
rect 3650 6830 3800 6840
rect 9700 6830 9990 6840
rect 1900 6820 2000 6830
rect 2300 6820 2450 6830
rect 3650 6820 3800 6830
rect 9700 6820 9990 6830
rect 1900 6810 2000 6820
rect 2300 6810 2450 6820
rect 3650 6810 3800 6820
rect 9700 6810 9990 6820
rect 1900 6800 2000 6810
rect 2300 6800 2450 6810
rect 3650 6800 3800 6810
rect 9700 6800 9990 6810
rect 1900 6790 1950 6800
rect 2000 6790 2050 6800
rect 2250 6790 2300 6800
rect 2450 6790 2650 6800
rect 3750 6790 3850 6800
rect 9700 6790 9850 6800
rect 9900 6790 9990 6800
rect 1900 6780 1950 6790
rect 2000 6780 2050 6790
rect 2250 6780 2300 6790
rect 2450 6780 2650 6790
rect 3750 6780 3850 6790
rect 9700 6780 9850 6790
rect 9900 6780 9990 6790
rect 1900 6770 1950 6780
rect 2000 6770 2050 6780
rect 2250 6770 2300 6780
rect 2450 6770 2650 6780
rect 3750 6770 3850 6780
rect 9700 6770 9850 6780
rect 9900 6770 9990 6780
rect 1900 6760 1950 6770
rect 2000 6760 2050 6770
rect 2250 6760 2300 6770
rect 2450 6760 2650 6770
rect 3750 6760 3850 6770
rect 9700 6760 9850 6770
rect 9900 6760 9990 6770
rect 1900 6750 1950 6760
rect 2000 6750 2050 6760
rect 2250 6750 2300 6760
rect 2450 6750 2650 6760
rect 3750 6750 3850 6760
rect 9700 6750 9850 6760
rect 9900 6750 9990 6760
rect 1900 6740 2000 6750
rect 2200 6740 2250 6750
rect 2550 6740 2600 6750
rect 2800 6740 3050 6750
rect 3800 6740 3850 6750
rect 9700 6740 9850 6750
rect 9950 6740 9990 6750
rect 1900 6730 2000 6740
rect 2200 6730 2250 6740
rect 2550 6730 2600 6740
rect 2800 6730 3050 6740
rect 3800 6730 3850 6740
rect 9700 6730 9850 6740
rect 9950 6730 9990 6740
rect 1900 6720 2000 6730
rect 2200 6720 2250 6730
rect 2550 6720 2600 6730
rect 2800 6720 3050 6730
rect 3800 6720 3850 6730
rect 9700 6720 9850 6730
rect 9950 6720 9990 6730
rect 1900 6710 2000 6720
rect 2200 6710 2250 6720
rect 2550 6710 2600 6720
rect 2800 6710 3050 6720
rect 3800 6710 3850 6720
rect 9700 6710 9850 6720
rect 9950 6710 9990 6720
rect 1900 6700 2000 6710
rect 2200 6700 2250 6710
rect 2550 6700 2600 6710
rect 2800 6700 3050 6710
rect 3800 6700 3850 6710
rect 9700 6700 9850 6710
rect 9950 6700 9990 6710
rect 1900 6690 1950 6700
rect 2600 6690 2650 6700
rect 3200 6690 3350 6700
rect 3850 6690 3900 6700
rect 9700 6690 9850 6700
rect 1900 6680 1950 6690
rect 2600 6680 2650 6690
rect 3200 6680 3350 6690
rect 3850 6680 3900 6690
rect 9700 6680 9850 6690
rect 1900 6670 1950 6680
rect 2600 6670 2650 6680
rect 3200 6670 3350 6680
rect 3850 6670 3900 6680
rect 9700 6670 9850 6680
rect 1900 6660 1950 6670
rect 2600 6660 2650 6670
rect 3200 6660 3350 6670
rect 3850 6660 3900 6670
rect 9700 6660 9850 6670
rect 1900 6650 1950 6660
rect 2600 6650 2650 6660
rect 3200 6650 3350 6660
rect 3850 6650 3900 6660
rect 9700 6650 9850 6660
rect 1850 6640 1900 6650
rect 2100 6640 2200 6650
rect 3450 6640 3550 6650
rect 1850 6630 1900 6640
rect 2100 6630 2200 6640
rect 3450 6630 3550 6640
rect 1850 6620 1900 6630
rect 2100 6620 2200 6630
rect 3450 6620 3550 6630
rect 1850 6610 1900 6620
rect 2100 6610 2200 6620
rect 3450 6610 3550 6620
rect 1850 6600 1900 6610
rect 2100 6600 2200 6610
rect 3450 6600 3550 6610
rect 1800 6590 1850 6600
rect 2000 6590 2050 6600
rect 2650 6590 2700 6600
rect 3600 6590 3650 6600
rect 1800 6580 1850 6590
rect 2000 6580 2050 6590
rect 2650 6580 2700 6590
rect 3600 6580 3650 6590
rect 1800 6570 1850 6580
rect 2000 6570 2050 6580
rect 2650 6570 2700 6580
rect 3600 6570 3650 6580
rect 1800 6560 1850 6570
rect 2000 6560 2050 6570
rect 2650 6560 2700 6570
rect 3600 6560 3650 6570
rect 1800 6550 1850 6560
rect 2000 6550 2050 6560
rect 2650 6550 2700 6560
rect 3600 6550 3650 6560
rect 1500 6540 1650 6550
rect 1850 6540 1900 6550
rect 2000 6540 2050 6550
rect 2600 6540 2650 6550
rect 3700 6540 3750 6550
rect 1500 6530 1650 6540
rect 1850 6530 1900 6540
rect 2000 6530 2050 6540
rect 2600 6530 2650 6540
rect 3700 6530 3750 6540
rect 1500 6520 1650 6530
rect 1850 6520 1900 6530
rect 2000 6520 2050 6530
rect 2600 6520 2650 6530
rect 3700 6520 3750 6530
rect 1500 6510 1650 6520
rect 1850 6510 1900 6520
rect 2000 6510 2050 6520
rect 2600 6510 2650 6520
rect 3700 6510 3750 6520
rect 1500 6500 1650 6510
rect 1850 6500 1900 6510
rect 2000 6500 2050 6510
rect 2600 6500 2650 6510
rect 3700 6500 3750 6510
rect 1400 6490 1450 6500
rect 1550 6490 1650 6500
rect 1900 6490 2100 6500
rect 3800 6490 3850 6500
rect 9950 6490 9990 6500
rect 1400 6480 1450 6490
rect 1550 6480 1650 6490
rect 1900 6480 2100 6490
rect 3800 6480 3850 6490
rect 9950 6480 9990 6490
rect 1400 6470 1450 6480
rect 1550 6470 1650 6480
rect 1900 6470 2100 6480
rect 3800 6470 3850 6480
rect 9950 6470 9990 6480
rect 1400 6460 1450 6470
rect 1550 6460 1650 6470
rect 1900 6460 2100 6470
rect 3800 6460 3850 6470
rect 9950 6460 9990 6470
rect 1400 6450 1450 6460
rect 1550 6450 1650 6460
rect 1900 6450 2100 6460
rect 3800 6450 3850 6460
rect 9950 6450 9990 6460
rect 1450 6440 1500 6450
rect 1550 6440 1600 6450
rect 2400 6440 2500 6450
rect 2550 6440 2600 6450
rect 3900 6440 3950 6450
rect 6400 6440 6550 6450
rect 9750 6440 9850 6450
rect 9900 6440 9950 6450
rect 1450 6430 1500 6440
rect 1550 6430 1600 6440
rect 2400 6430 2500 6440
rect 2550 6430 2600 6440
rect 3900 6430 3950 6440
rect 6400 6430 6550 6440
rect 9750 6430 9850 6440
rect 9900 6430 9950 6440
rect 1450 6420 1500 6430
rect 1550 6420 1600 6430
rect 2400 6420 2500 6430
rect 2550 6420 2600 6430
rect 3900 6420 3950 6430
rect 6400 6420 6550 6430
rect 9750 6420 9850 6430
rect 9900 6420 9950 6430
rect 1450 6410 1500 6420
rect 1550 6410 1600 6420
rect 2400 6410 2500 6420
rect 2550 6410 2600 6420
rect 3900 6410 3950 6420
rect 6400 6410 6550 6420
rect 9750 6410 9850 6420
rect 9900 6410 9950 6420
rect 1450 6400 1500 6410
rect 1550 6400 1600 6410
rect 2400 6400 2500 6410
rect 2550 6400 2600 6410
rect 3900 6400 3950 6410
rect 6400 6400 6550 6410
rect 9750 6400 9850 6410
rect 9900 6400 9950 6410
rect 1450 6390 1500 6400
rect 1550 6390 1600 6400
rect 2450 6390 2500 6400
rect 6450 6390 6550 6400
rect 9700 6390 9850 6400
rect 9900 6390 9950 6400
rect 1450 6380 1500 6390
rect 1550 6380 1600 6390
rect 2450 6380 2500 6390
rect 6450 6380 6550 6390
rect 9700 6380 9850 6390
rect 9900 6380 9950 6390
rect 1450 6370 1500 6380
rect 1550 6370 1600 6380
rect 2450 6370 2500 6380
rect 6450 6370 6550 6380
rect 9700 6370 9850 6380
rect 9900 6370 9950 6380
rect 1450 6360 1500 6370
rect 1550 6360 1600 6370
rect 2450 6360 2500 6370
rect 6450 6360 6550 6370
rect 9700 6360 9850 6370
rect 9900 6360 9950 6370
rect 1450 6350 1500 6360
rect 1550 6350 1600 6360
rect 2450 6350 2500 6360
rect 6450 6350 6550 6360
rect 9700 6350 9850 6360
rect 9900 6350 9950 6360
rect 1450 6340 1500 6350
rect 1700 6340 1800 6350
rect 4050 6340 4100 6350
rect 9650 6340 9950 6350
rect 1450 6330 1500 6340
rect 1700 6330 1800 6340
rect 4050 6330 4100 6340
rect 9650 6330 9950 6340
rect 1450 6320 1500 6330
rect 1700 6320 1800 6330
rect 4050 6320 4100 6330
rect 9650 6320 9950 6330
rect 1450 6310 1500 6320
rect 1700 6310 1800 6320
rect 4050 6310 4100 6320
rect 9650 6310 9950 6320
rect 1450 6300 1500 6310
rect 1700 6300 1800 6310
rect 4050 6300 4100 6310
rect 9650 6300 9950 6310
rect 1650 6290 1800 6300
rect 4100 6290 4150 6300
rect 5400 6290 5500 6300
rect 6650 6290 6750 6300
rect 1650 6280 1800 6290
rect 4100 6280 4150 6290
rect 5400 6280 5500 6290
rect 6650 6280 6750 6290
rect 1650 6270 1800 6280
rect 4100 6270 4150 6280
rect 5400 6270 5500 6280
rect 6650 6270 6750 6280
rect 1650 6260 1800 6270
rect 4100 6260 4150 6270
rect 5400 6260 5500 6270
rect 6650 6260 6750 6270
rect 1650 6250 1800 6260
rect 4100 6250 4150 6260
rect 5400 6250 5500 6260
rect 6650 6250 6750 6260
rect 1550 6240 1600 6250
rect 1650 6240 1750 6250
rect 2450 6240 2500 6250
rect 4150 6240 4200 6250
rect 5350 6240 5450 6250
rect 6700 6240 6750 6250
rect 9750 6240 9800 6250
rect 1550 6230 1600 6240
rect 1650 6230 1750 6240
rect 2450 6230 2500 6240
rect 4150 6230 4200 6240
rect 5350 6230 5450 6240
rect 6700 6230 6750 6240
rect 9750 6230 9800 6240
rect 1550 6220 1600 6230
rect 1650 6220 1750 6230
rect 2450 6220 2500 6230
rect 4150 6220 4200 6230
rect 5350 6220 5450 6230
rect 6700 6220 6750 6230
rect 9750 6220 9800 6230
rect 1550 6210 1600 6220
rect 1650 6210 1750 6220
rect 2450 6210 2500 6220
rect 4150 6210 4200 6220
rect 5350 6210 5450 6220
rect 6700 6210 6750 6220
rect 9750 6210 9800 6220
rect 1550 6200 1600 6210
rect 1650 6200 1750 6210
rect 2450 6200 2500 6210
rect 4150 6200 4200 6210
rect 5350 6200 5450 6210
rect 6700 6200 6750 6210
rect 9750 6200 9800 6210
rect 1550 6190 1600 6200
rect 4200 6190 4250 6200
rect 5350 6190 5400 6200
rect 9400 6190 9500 6200
rect 9550 6190 9600 6200
rect 9700 6190 9800 6200
rect 1550 6180 1600 6190
rect 4200 6180 4250 6190
rect 5350 6180 5400 6190
rect 9400 6180 9500 6190
rect 9550 6180 9600 6190
rect 9700 6180 9800 6190
rect 1550 6170 1600 6180
rect 4200 6170 4250 6180
rect 5350 6170 5400 6180
rect 9400 6170 9500 6180
rect 9550 6170 9600 6180
rect 9700 6170 9800 6180
rect 1550 6160 1600 6170
rect 4200 6160 4250 6170
rect 5350 6160 5400 6170
rect 9400 6160 9500 6170
rect 9550 6160 9600 6170
rect 9700 6160 9800 6170
rect 1550 6150 1600 6160
rect 4200 6150 4250 6160
rect 5350 6150 5400 6160
rect 9400 6150 9500 6160
rect 9550 6150 9600 6160
rect 9700 6150 9800 6160
rect 2450 6140 2500 6150
rect 3850 6140 3900 6150
rect 3950 6140 4000 6150
rect 5300 6140 5400 6150
rect 9250 6140 9350 6150
rect 9600 6140 9700 6150
rect 2450 6130 2500 6140
rect 3850 6130 3900 6140
rect 3950 6130 4000 6140
rect 5300 6130 5400 6140
rect 9250 6130 9350 6140
rect 9600 6130 9700 6140
rect 2450 6120 2500 6130
rect 3850 6120 3900 6130
rect 3950 6120 4000 6130
rect 5300 6120 5400 6130
rect 9250 6120 9350 6130
rect 9600 6120 9700 6130
rect 2450 6110 2500 6120
rect 3850 6110 3900 6120
rect 3950 6110 4000 6120
rect 5300 6110 5400 6120
rect 9250 6110 9350 6120
rect 9600 6110 9700 6120
rect 2450 6100 2500 6110
rect 3850 6100 3900 6110
rect 3950 6100 4000 6110
rect 5300 6100 5400 6110
rect 9250 6100 9350 6110
rect 9600 6100 9700 6110
rect 1350 6090 1450 6100
rect 1550 6090 1600 6100
rect 3750 6090 3800 6100
rect 4000 6090 4050 6100
rect 4250 6090 4300 6100
rect 9500 6090 9550 6100
rect 9600 6090 9750 6100
rect 9800 6090 9850 6100
rect 1350 6080 1450 6090
rect 1550 6080 1600 6090
rect 3750 6080 3800 6090
rect 4000 6080 4050 6090
rect 4250 6080 4300 6090
rect 9500 6080 9550 6090
rect 9600 6080 9750 6090
rect 9800 6080 9850 6090
rect 1350 6070 1450 6080
rect 1550 6070 1600 6080
rect 3750 6070 3800 6080
rect 4000 6070 4050 6080
rect 4250 6070 4300 6080
rect 9500 6070 9550 6080
rect 9600 6070 9750 6080
rect 9800 6070 9850 6080
rect 1350 6060 1450 6070
rect 1550 6060 1600 6070
rect 3750 6060 3800 6070
rect 4000 6060 4050 6070
rect 4250 6060 4300 6070
rect 9500 6060 9550 6070
rect 9600 6060 9750 6070
rect 9800 6060 9850 6070
rect 1350 6050 1450 6060
rect 1550 6050 1600 6060
rect 3750 6050 3800 6060
rect 4000 6050 4050 6060
rect 4250 6050 4300 6060
rect 9500 6050 9550 6060
rect 9600 6050 9750 6060
rect 9800 6050 9850 6060
rect 1300 6040 1350 6050
rect 2500 6040 2550 6050
rect 3150 6040 3300 6050
rect 4050 6040 4100 6050
rect 5250 6040 5350 6050
rect 9500 6040 9550 6050
rect 9650 6040 9750 6050
rect 9800 6040 9850 6050
rect 1300 6030 1350 6040
rect 2500 6030 2550 6040
rect 3150 6030 3300 6040
rect 4050 6030 4100 6040
rect 5250 6030 5350 6040
rect 9500 6030 9550 6040
rect 9650 6030 9750 6040
rect 9800 6030 9850 6040
rect 1300 6020 1350 6030
rect 2500 6020 2550 6030
rect 3150 6020 3300 6030
rect 4050 6020 4100 6030
rect 5250 6020 5350 6030
rect 9500 6020 9550 6030
rect 9650 6020 9750 6030
rect 9800 6020 9850 6030
rect 1300 6010 1350 6020
rect 2500 6010 2550 6020
rect 3150 6010 3300 6020
rect 4050 6010 4100 6020
rect 5250 6010 5350 6020
rect 9500 6010 9550 6020
rect 9650 6010 9750 6020
rect 9800 6010 9850 6020
rect 1300 6000 1350 6010
rect 2500 6000 2550 6010
rect 3150 6000 3300 6010
rect 4050 6000 4100 6010
rect 5250 6000 5350 6010
rect 9500 6000 9550 6010
rect 9650 6000 9750 6010
rect 9800 6000 9850 6010
rect 1200 5990 1350 6000
rect 1600 5990 1650 6000
rect 2550 5990 2600 6000
rect 3100 5990 3150 6000
rect 3250 5990 3300 6000
rect 3700 5990 3750 6000
rect 4150 5990 4200 6000
rect 5200 5990 5250 6000
rect 5300 5990 5350 6000
rect 9500 5990 9550 6000
rect 9650 5990 9750 6000
rect 1200 5980 1350 5990
rect 1600 5980 1650 5990
rect 2550 5980 2600 5990
rect 3100 5980 3150 5990
rect 3250 5980 3300 5990
rect 3700 5980 3750 5990
rect 4150 5980 4200 5990
rect 5200 5980 5250 5990
rect 5300 5980 5350 5990
rect 9500 5980 9550 5990
rect 9650 5980 9750 5990
rect 1200 5970 1350 5980
rect 1600 5970 1650 5980
rect 2550 5970 2600 5980
rect 3100 5970 3150 5980
rect 3250 5970 3300 5980
rect 3700 5970 3750 5980
rect 4150 5970 4200 5980
rect 5200 5970 5250 5980
rect 5300 5970 5350 5980
rect 9500 5970 9550 5980
rect 9650 5970 9750 5980
rect 1200 5960 1350 5970
rect 1600 5960 1650 5970
rect 2550 5960 2600 5970
rect 3100 5960 3150 5970
rect 3250 5960 3300 5970
rect 3700 5960 3750 5970
rect 4150 5960 4200 5970
rect 5200 5960 5250 5970
rect 5300 5960 5350 5970
rect 9500 5960 9550 5970
rect 9650 5960 9750 5970
rect 1200 5950 1350 5960
rect 1600 5950 1650 5960
rect 2550 5950 2600 5960
rect 3100 5950 3150 5960
rect 3250 5950 3300 5960
rect 3700 5950 3750 5960
rect 4150 5950 4200 5960
rect 5200 5950 5250 5960
rect 5300 5950 5350 5960
rect 9500 5950 9550 5960
rect 9650 5950 9750 5960
rect 1050 5940 1200 5950
rect 1650 5940 1700 5950
rect 2600 5940 2650 5950
rect 3050 5940 3100 5950
rect 3250 5940 3300 5950
rect 3700 5940 3750 5950
rect 6850 5940 6950 5950
rect 9700 5940 9750 5950
rect 1050 5930 1200 5940
rect 1650 5930 1700 5940
rect 2600 5930 2650 5940
rect 3050 5930 3100 5940
rect 3250 5930 3300 5940
rect 3700 5930 3750 5940
rect 6850 5930 6950 5940
rect 9700 5930 9750 5940
rect 1050 5920 1200 5930
rect 1650 5920 1700 5930
rect 2600 5920 2650 5930
rect 3050 5920 3100 5930
rect 3250 5920 3300 5930
rect 3700 5920 3750 5930
rect 6850 5920 6950 5930
rect 9700 5920 9750 5930
rect 1050 5910 1200 5920
rect 1650 5910 1700 5920
rect 2600 5910 2650 5920
rect 3050 5910 3100 5920
rect 3250 5910 3300 5920
rect 3700 5910 3750 5920
rect 6850 5910 6950 5920
rect 9700 5910 9750 5920
rect 1050 5900 1200 5910
rect 1650 5900 1700 5910
rect 2600 5900 2650 5910
rect 3050 5900 3100 5910
rect 3250 5900 3300 5910
rect 3700 5900 3750 5910
rect 6850 5900 6950 5910
rect 9700 5900 9750 5910
rect 1000 5890 1050 5900
rect 1700 5890 1750 5900
rect 2650 5890 2700 5900
rect 2900 5890 3000 5900
rect 3700 5890 3750 5900
rect 5150 5890 5200 5900
rect 6850 5890 6950 5900
rect 8500 5890 8600 5900
rect 9350 5890 9450 5900
rect 9850 5890 9900 5900
rect 1000 5880 1050 5890
rect 1700 5880 1750 5890
rect 2650 5880 2700 5890
rect 2900 5880 3000 5890
rect 3700 5880 3750 5890
rect 5150 5880 5200 5890
rect 6850 5880 6950 5890
rect 8500 5880 8600 5890
rect 9350 5880 9450 5890
rect 9850 5880 9900 5890
rect 1000 5870 1050 5880
rect 1700 5870 1750 5880
rect 2650 5870 2700 5880
rect 2900 5870 3000 5880
rect 3700 5870 3750 5880
rect 5150 5870 5200 5880
rect 6850 5870 6950 5880
rect 8500 5870 8600 5880
rect 9350 5870 9450 5880
rect 9850 5870 9900 5880
rect 1000 5860 1050 5870
rect 1700 5860 1750 5870
rect 2650 5860 2700 5870
rect 2900 5860 3000 5870
rect 3700 5860 3750 5870
rect 5150 5860 5200 5870
rect 6850 5860 6950 5870
rect 8500 5860 8600 5870
rect 9350 5860 9450 5870
rect 9850 5860 9900 5870
rect 1000 5850 1050 5860
rect 1700 5850 1750 5860
rect 2650 5850 2700 5860
rect 2900 5850 3000 5860
rect 3700 5850 3750 5860
rect 5150 5850 5200 5860
rect 6850 5850 6950 5860
rect 8500 5850 8600 5860
rect 9350 5850 9450 5860
rect 9850 5850 9900 5860
rect 1800 5840 1850 5850
rect 2700 5840 2850 5850
rect 5250 5840 5300 5850
rect 6850 5840 6950 5850
rect 8400 5840 8600 5850
rect 9300 5840 9350 5850
rect 1800 5830 1850 5840
rect 2700 5830 2850 5840
rect 5250 5830 5300 5840
rect 6850 5830 6950 5840
rect 8400 5830 8600 5840
rect 9300 5830 9350 5840
rect 1800 5820 1850 5830
rect 2700 5820 2850 5830
rect 5250 5820 5300 5830
rect 6850 5820 6950 5830
rect 8400 5820 8600 5830
rect 9300 5820 9350 5830
rect 1800 5810 1850 5820
rect 2700 5810 2850 5820
rect 5250 5810 5300 5820
rect 6850 5810 6950 5820
rect 8400 5810 8600 5820
rect 9300 5810 9350 5820
rect 1800 5800 1850 5810
rect 2700 5800 2850 5810
rect 5250 5800 5300 5810
rect 6850 5800 6950 5810
rect 8400 5800 8600 5810
rect 9300 5800 9350 5810
rect 900 5790 950 5800
rect 1800 5790 1850 5800
rect 2700 5790 2800 5800
rect 3700 5790 3750 5800
rect 5100 5790 5150 5800
rect 5250 5790 5300 5800
rect 6850 5790 6950 5800
rect 8300 5790 8350 5800
rect 8450 5790 8650 5800
rect 9100 5790 9250 5800
rect 900 5780 950 5790
rect 1800 5780 1850 5790
rect 2700 5780 2800 5790
rect 3700 5780 3750 5790
rect 5100 5780 5150 5790
rect 5250 5780 5300 5790
rect 6850 5780 6950 5790
rect 8300 5780 8350 5790
rect 8450 5780 8650 5790
rect 9100 5780 9250 5790
rect 900 5770 950 5780
rect 1800 5770 1850 5780
rect 2700 5770 2800 5780
rect 3700 5770 3750 5780
rect 5100 5770 5150 5780
rect 5250 5770 5300 5780
rect 6850 5770 6950 5780
rect 8300 5770 8350 5780
rect 8450 5770 8650 5780
rect 9100 5770 9250 5780
rect 900 5760 950 5770
rect 1800 5760 1850 5770
rect 2700 5760 2800 5770
rect 3700 5760 3750 5770
rect 5100 5760 5150 5770
rect 5250 5760 5300 5770
rect 6850 5760 6950 5770
rect 8300 5760 8350 5770
rect 8450 5760 8650 5770
rect 9100 5760 9250 5770
rect 900 5750 950 5760
rect 1800 5750 1850 5760
rect 2700 5750 2800 5760
rect 3700 5750 3750 5760
rect 5100 5750 5150 5760
rect 5250 5750 5300 5760
rect 6850 5750 6950 5760
rect 8300 5750 8350 5760
rect 8450 5750 8650 5760
rect 9100 5750 9250 5760
rect 850 5740 900 5750
rect 1100 5740 1250 5750
rect 1800 5740 1850 5750
rect 2600 5740 2750 5750
rect 3300 5740 3350 5750
rect 3700 5740 3750 5750
rect 3850 5740 3900 5750
rect 5100 5740 5150 5750
rect 8500 5740 8650 5750
rect 8750 5740 8850 5750
rect 8950 5740 9050 5750
rect 9900 5740 9950 5750
rect 850 5730 900 5740
rect 1100 5730 1250 5740
rect 1800 5730 1850 5740
rect 2600 5730 2750 5740
rect 3300 5730 3350 5740
rect 3700 5730 3750 5740
rect 3850 5730 3900 5740
rect 5100 5730 5150 5740
rect 8500 5730 8650 5740
rect 8750 5730 8850 5740
rect 8950 5730 9050 5740
rect 9900 5730 9950 5740
rect 850 5720 900 5730
rect 1100 5720 1250 5730
rect 1800 5720 1850 5730
rect 2600 5720 2750 5730
rect 3300 5720 3350 5730
rect 3700 5720 3750 5730
rect 3850 5720 3900 5730
rect 5100 5720 5150 5730
rect 8500 5720 8650 5730
rect 8750 5720 8850 5730
rect 8950 5720 9050 5730
rect 9900 5720 9950 5730
rect 850 5710 900 5720
rect 1100 5710 1250 5720
rect 1800 5710 1850 5720
rect 2600 5710 2750 5720
rect 3300 5710 3350 5720
rect 3700 5710 3750 5720
rect 3850 5710 3900 5720
rect 5100 5710 5150 5720
rect 8500 5710 8650 5720
rect 8750 5710 8850 5720
rect 8950 5710 9050 5720
rect 9900 5710 9950 5720
rect 850 5700 900 5710
rect 1100 5700 1250 5710
rect 1800 5700 1850 5710
rect 2600 5700 2750 5710
rect 3300 5700 3350 5710
rect 3700 5700 3750 5710
rect 3850 5700 3900 5710
rect 5100 5700 5150 5710
rect 8500 5700 8650 5710
rect 8750 5700 8850 5710
rect 8950 5700 9050 5710
rect 9900 5700 9950 5710
rect 1050 5690 1100 5700
rect 1150 5690 1250 5700
rect 2550 5690 2650 5700
rect 3300 5690 3350 5700
rect 3650 5690 3700 5700
rect 7950 5690 8000 5700
rect 8550 5690 8700 5700
rect 8750 5690 8800 5700
rect 8950 5690 9000 5700
rect 1050 5680 1100 5690
rect 1150 5680 1250 5690
rect 2550 5680 2650 5690
rect 3300 5680 3350 5690
rect 3650 5680 3700 5690
rect 7950 5680 8000 5690
rect 8550 5680 8700 5690
rect 8750 5680 8800 5690
rect 8950 5680 9000 5690
rect 1050 5670 1100 5680
rect 1150 5670 1250 5680
rect 2550 5670 2650 5680
rect 3300 5670 3350 5680
rect 3650 5670 3700 5680
rect 7950 5670 8000 5680
rect 8550 5670 8700 5680
rect 8750 5670 8800 5680
rect 8950 5670 9000 5680
rect 1050 5660 1100 5670
rect 1150 5660 1250 5670
rect 2550 5660 2650 5670
rect 3300 5660 3350 5670
rect 3650 5660 3700 5670
rect 7950 5660 8000 5670
rect 8550 5660 8700 5670
rect 8750 5660 8800 5670
rect 8950 5660 9000 5670
rect 1050 5650 1100 5660
rect 1150 5650 1250 5660
rect 2550 5650 2650 5660
rect 3300 5650 3350 5660
rect 3650 5650 3700 5660
rect 7950 5650 8000 5660
rect 8550 5650 8700 5660
rect 8750 5650 8800 5660
rect 8950 5650 9000 5660
rect 800 5640 850 5650
rect 1850 5640 1900 5650
rect 2550 5640 2600 5650
rect 3400 5640 3450 5650
rect 3650 5640 3700 5650
rect 6900 5640 6950 5650
rect 8900 5640 9000 5650
rect 9050 5640 9100 5650
rect 800 5630 850 5640
rect 1850 5630 1900 5640
rect 2550 5630 2600 5640
rect 3400 5630 3450 5640
rect 3650 5630 3700 5640
rect 6900 5630 6950 5640
rect 8900 5630 9000 5640
rect 9050 5630 9100 5640
rect 800 5620 850 5630
rect 1850 5620 1900 5630
rect 2550 5620 2600 5630
rect 3400 5620 3450 5630
rect 3650 5620 3700 5630
rect 6900 5620 6950 5630
rect 8900 5620 9000 5630
rect 9050 5620 9100 5630
rect 800 5610 850 5620
rect 1850 5610 1900 5620
rect 2550 5610 2600 5620
rect 3400 5610 3450 5620
rect 3650 5610 3700 5620
rect 6900 5610 6950 5620
rect 8900 5610 9000 5620
rect 9050 5610 9100 5620
rect 800 5600 850 5610
rect 1850 5600 1900 5610
rect 2550 5600 2600 5610
rect 3400 5600 3450 5610
rect 3650 5600 3700 5610
rect 6900 5600 6950 5610
rect 8900 5600 9000 5610
rect 9050 5600 9100 5610
rect 700 5590 750 5600
rect 1850 5590 1900 5600
rect 2500 5590 2600 5600
rect 3300 5590 3350 5600
rect 3400 5590 3450 5600
rect 3600 5590 3650 5600
rect 5200 5590 5250 5600
rect 5650 5590 5800 5600
rect 8400 5590 8500 5600
rect 8750 5590 8850 5600
rect 9100 5590 9150 5600
rect 9950 5590 9990 5600
rect 700 5580 750 5590
rect 1850 5580 1900 5590
rect 2500 5580 2600 5590
rect 3300 5580 3350 5590
rect 3400 5580 3450 5590
rect 3600 5580 3650 5590
rect 5200 5580 5250 5590
rect 5650 5580 5800 5590
rect 8400 5580 8500 5590
rect 8750 5580 8850 5590
rect 9100 5580 9150 5590
rect 9950 5580 9990 5590
rect 700 5570 750 5580
rect 1850 5570 1900 5580
rect 2500 5570 2600 5580
rect 3300 5570 3350 5580
rect 3400 5570 3450 5580
rect 3600 5570 3650 5580
rect 5200 5570 5250 5580
rect 5650 5570 5800 5580
rect 8400 5570 8500 5580
rect 8750 5570 8850 5580
rect 9100 5570 9150 5580
rect 9950 5570 9990 5580
rect 700 5560 750 5570
rect 1850 5560 1900 5570
rect 2500 5560 2600 5570
rect 3300 5560 3350 5570
rect 3400 5560 3450 5570
rect 3600 5560 3650 5570
rect 5200 5560 5250 5570
rect 5650 5560 5800 5570
rect 8400 5560 8500 5570
rect 8750 5560 8850 5570
rect 9100 5560 9150 5570
rect 9950 5560 9990 5570
rect 700 5550 750 5560
rect 1850 5550 1900 5560
rect 2500 5550 2600 5560
rect 3300 5550 3350 5560
rect 3400 5550 3450 5560
rect 3600 5550 3650 5560
rect 5200 5550 5250 5560
rect 5650 5550 5800 5560
rect 8400 5550 8500 5560
rect 8750 5550 8850 5560
rect 9100 5550 9150 5560
rect 9950 5550 9990 5560
rect 650 5540 700 5550
rect 900 5540 1000 5550
rect 1850 5540 1900 5550
rect 2450 5540 2550 5550
rect 3300 5540 3350 5550
rect 3500 5540 3550 5550
rect 3600 5540 3650 5550
rect 5200 5540 5250 5550
rect 5750 5540 5900 5550
rect 6250 5540 6500 5550
rect 7400 5540 7450 5550
rect 8250 5540 8350 5550
rect 8600 5540 8700 5550
rect 650 5530 700 5540
rect 900 5530 1000 5540
rect 1850 5530 1900 5540
rect 2450 5530 2550 5540
rect 3300 5530 3350 5540
rect 3500 5530 3550 5540
rect 3600 5530 3650 5540
rect 5200 5530 5250 5540
rect 5750 5530 5900 5540
rect 6250 5530 6500 5540
rect 7400 5530 7450 5540
rect 8250 5530 8350 5540
rect 8600 5530 8700 5540
rect 650 5520 700 5530
rect 900 5520 1000 5530
rect 1850 5520 1900 5530
rect 2450 5520 2550 5530
rect 3300 5520 3350 5530
rect 3500 5520 3550 5530
rect 3600 5520 3650 5530
rect 5200 5520 5250 5530
rect 5750 5520 5900 5530
rect 6250 5520 6500 5530
rect 7400 5520 7450 5530
rect 8250 5520 8350 5530
rect 8600 5520 8700 5530
rect 650 5510 700 5520
rect 900 5510 1000 5520
rect 1850 5510 1900 5520
rect 2450 5510 2550 5520
rect 3300 5510 3350 5520
rect 3500 5510 3550 5520
rect 3600 5510 3650 5520
rect 5200 5510 5250 5520
rect 5750 5510 5900 5520
rect 6250 5510 6500 5520
rect 7400 5510 7450 5520
rect 8250 5510 8350 5520
rect 8600 5510 8700 5520
rect 650 5500 700 5510
rect 900 5500 1000 5510
rect 1850 5500 1900 5510
rect 2450 5500 2550 5510
rect 3300 5500 3350 5510
rect 3500 5500 3550 5510
rect 3600 5500 3650 5510
rect 5200 5500 5250 5510
rect 5750 5500 5900 5510
rect 6250 5500 6500 5510
rect 7400 5500 7450 5510
rect 8250 5500 8350 5510
rect 8600 5500 8700 5510
rect 600 5490 650 5500
rect 900 5490 1000 5500
rect 1900 5490 1950 5500
rect 2450 5490 2550 5500
rect 3300 5490 3350 5500
rect 5700 5490 5900 5500
rect 6200 5490 6250 5500
rect 6350 5490 6450 5500
rect 8000 5490 8050 5500
rect 8100 5490 8200 5500
rect 8400 5490 8500 5500
rect 600 5480 650 5490
rect 900 5480 1000 5490
rect 1900 5480 1950 5490
rect 2450 5480 2550 5490
rect 3300 5480 3350 5490
rect 5700 5480 5900 5490
rect 6200 5480 6250 5490
rect 6350 5480 6450 5490
rect 8000 5480 8050 5490
rect 8100 5480 8200 5490
rect 8400 5480 8500 5490
rect 600 5470 650 5480
rect 900 5470 1000 5480
rect 1900 5470 1950 5480
rect 2450 5470 2550 5480
rect 3300 5470 3350 5480
rect 5700 5470 5900 5480
rect 6200 5470 6250 5480
rect 6350 5470 6450 5480
rect 8000 5470 8050 5480
rect 8100 5470 8200 5480
rect 8400 5470 8500 5480
rect 600 5460 650 5470
rect 900 5460 1000 5470
rect 1900 5460 1950 5470
rect 2450 5460 2550 5470
rect 3300 5460 3350 5470
rect 5700 5460 5900 5470
rect 6200 5460 6250 5470
rect 6350 5460 6450 5470
rect 8000 5460 8050 5470
rect 8100 5460 8200 5470
rect 8400 5460 8500 5470
rect 600 5450 650 5460
rect 900 5450 1000 5460
rect 1900 5450 1950 5460
rect 2450 5450 2550 5460
rect 3300 5450 3350 5460
rect 5700 5450 5900 5460
rect 6200 5450 6250 5460
rect 6350 5450 6450 5460
rect 8000 5450 8050 5460
rect 8100 5450 8200 5460
rect 8400 5450 8500 5460
rect 600 5440 650 5450
rect 1900 5440 1950 5450
rect 2400 5440 2450 5450
rect 2550 5440 2600 5450
rect 2900 5440 2950 5450
rect 3250 5440 3300 5450
rect 5500 5440 5600 5450
rect 5650 5440 5750 5450
rect 5800 5440 5900 5450
rect 6200 5440 6250 5450
rect 6400 5440 6500 5450
rect 7400 5440 7450 5450
rect 8000 5440 8150 5450
rect 8250 5440 8350 5450
rect 9400 5440 9450 5450
rect 9600 5440 9650 5450
rect 600 5430 650 5440
rect 1900 5430 1950 5440
rect 2400 5430 2450 5440
rect 2550 5430 2600 5440
rect 2900 5430 2950 5440
rect 3250 5430 3300 5440
rect 5500 5430 5600 5440
rect 5650 5430 5750 5440
rect 5800 5430 5900 5440
rect 6200 5430 6250 5440
rect 6400 5430 6500 5440
rect 7400 5430 7450 5440
rect 8000 5430 8150 5440
rect 8250 5430 8350 5440
rect 9400 5430 9450 5440
rect 9600 5430 9650 5440
rect 600 5420 650 5430
rect 1900 5420 1950 5430
rect 2400 5420 2450 5430
rect 2550 5420 2600 5430
rect 2900 5420 2950 5430
rect 3250 5420 3300 5430
rect 5500 5420 5600 5430
rect 5650 5420 5750 5430
rect 5800 5420 5900 5430
rect 6200 5420 6250 5430
rect 6400 5420 6500 5430
rect 7400 5420 7450 5430
rect 8000 5420 8150 5430
rect 8250 5420 8350 5430
rect 9400 5420 9450 5430
rect 9600 5420 9650 5430
rect 600 5410 650 5420
rect 1900 5410 1950 5420
rect 2400 5410 2450 5420
rect 2550 5410 2600 5420
rect 2900 5410 2950 5420
rect 3250 5410 3300 5420
rect 5500 5410 5600 5420
rect 5650 5410 5750 5420
rect 5800 5410 5900 5420
rect 6200 5410 6250 5420
rect 6400 5410 6500 5420
rect 7400 5410 7450 5420
rect 8000 5410 8150 5420
rect 8250 5410 8350 5420
rect 9400 5410 9450 5420
rect 9600 5410 9650 5420
rect 600 5400 650 5410
rect 1900 5400 1950 5410
rect 2400 5400 2450 5410
rect 2550 5400 2600 5410
rect 2900 5400 2950 5410
rect 3250 5400 3300 5410
rect 5500 5400 5600 5410
rect 5650 5400 5750 5410
rect 5800 5400 5900 5410
rect 6200 5400 6250 5410
rect 6400 5400 6500 5410
rect 7400 5400 7450 5410
rect 8000 5400 8150 5410
rect 8250 5400 8350 5410
rect 9400 5400 9450 5410
rect 9600 5400 9650 5410
rect 1900 5390 1950 5400
rect 2400 5390 2500 5400
rect 2550 5390 2600 5400
rect 2900 5390 3200 5400
rect 3500 5390 3550 5400
rect 5100 5390 5150 5400
rect 5600 5390 5750 5400
rect 5800 5390 5850 5400
rect 6200 5390 6250 5400
rect 6550 5390 6650 5400
rect 7450 5390 7500 5400
rect 7800 5390 7850 5400
rect 8000 5390 8100 5400
rect 8150 5390 8200 5400
rect 8950 5390 9000 5400
rect 9050 5390 9100 5400
rect 9600 5390 9650 5400
rect 1900 5380 1950 5390
rect 2400 5380 2500 5390
rect 2550 5380 2600 5390
rect 2900 5380 3200 5390
rect 3500 5380 3550 5390
rect 5100 5380 5150 5390
rect 5600 5380 5750 5390
rect 5800 5380 5850 5390
rect 6200 5380 6250 5390
rect 6550 5380 6650 5390
rect 7450 5380 7500 5390
rect 7800 5380 7850 5390
rect 8000 5380 8100 5390
rect 8150 5380 8200 5390
rect 8950 5380 9000 5390
rect 9050 5380 9100 5390
rect 9600 5380 9650 5390
rect 1900 5370 1950 5380
rect 2400 5370 2500 5380
rect 2550 5370 2600 5380
rect 2900 5370 3200 5380
rect 3500 5370 3550 5380
rect 5100 5370 5150 5380
rect 5600 5370 5750 5380
rect 5800 5370 5850 5380
rect 6200 5370 6250 5380
rect 6550 5370 6650 5380
rect 7450 5370 7500 5380
rect 7800 5370 7850 5380
rect 8000 5370 8100 5380
rect 8150 5370 8200 5380
rect 8950 5370 9000 5380
rect 9050 5370 9100 5380
rect 9600 5370 9650 5380
rect 1900 5360 1950 5370
rect 2400 5360 2500 5370
rect 2550 5360 2600 5370
rect 2900 5360 3200 5370
rect 3500 5360 3550 5370
rect 5100 5360 5150 5370
rect 5600 5360 5750 5370
rect 5800 5360 5850 5370
rect 6200 5360 6250 5370
rect 6550 5360 6650 5370
rect 7450 5360 7500 5370
rect 7800 5360 7850 5370
rect 8000 5360 8100 5370
rect 8150 5360 8200 5370
rect 8950 5360 9000 5370
rect 9050 5360 9100 5370
rect 9600 5360 9650 5370
rect 1900 5350 1950 5360
rect 2400 5350 2500 5360
rect 2550 5350 2600 5360
rect 2900 5350 3200 5360
rect 3500 5350 3550 5360
rect 5100 5350 5150 5360
rect 5600 5350 5750 5360
rect 5800 5350 5850 5360
rect 6200 5350 6250 5360
rect 6550 5350 6650 5360
rect 7450 5350 7500 5360
rect 7800 5350 7850 5360
rect 8000 5350 8100 5360
rect 8150 5350 8200 5360
rect 8950 5350 9000 5360
rect 9050 5350 9100 5360
rect 9600 5350 9650 5360
rect 1900 5340 2000 5350
rect 2400 5340 2450 5350
rect 2550 5340 2600 5350
rect 2750 5340 3050 5350
rect 5150 5340 5200 5350
rect 6200 5340 6500 5350
rect 7400 5340 7500 5350
rect 7600 5340 7750 5350
rect 7800 5340 7900 5350
rect 8850 5340 8950 5350
rect 9000 5340 9100 5350
rect 9150 5340 9250 5350
rect 9900 5340 9990 5350
rect 1900 5330 2000 5340
rect 2400 5330 2450 5340
rect 2550 5330 2600 5340
rect 2750 5330 3050 5340
rect 5150 5330 5200 5340
rect 6200 5330 6500 5340
rect 7400 5330 7500 5340
rect 7600 5330 7750 5340
rect 7800 5330 7900 5340
rect 8850 5330 8950 5340
rect 9000 5330 9100 5340
rect 9150 5330 9250 5340
rect 9900 5330 9990 5340
rect 1900 5320 2000 5330
rect 2400 5320 2450 5330
rect 2550 5320 2600 5330
rect 2750 5320 3050 5330
rect 5150 5320 5200 5330
rect 6200 5320 6500 5330
rect 7400 5320 7500 5330
rect 7600 5320 7750 5330
rect 7800 5320 7900 5330
rect 8850 5320 8950 5330
rect 9000 5320 9100 5330
rect 9150 5320 9250 5330
rect 9900 5320 9990 5330
rect 1900 5310 2000 5320
rect 2400 5310 2450 5320
rect 2550 5310 2600 5320
rect 2750 5310 3050 5320
rect 5150 5310 5200 5320
rect 6200 5310 6500 5320
rect 7400 5310 7500 5320
rect 7600 5310 7750 5320
rect 7800 5310 7900 5320
rect 8850 5310 8950 5320
rect 9000 5310 9100 5320
rect 9150 5310 9250 5320
rect 9900 5310 9990 5320
rect 1900 5300 2000 5310
rect 2400 5300 2450 5310
rect 2550 5300 2600 5310
rect 2750 5300 3050 5310
rect 5150 5300 5200 5310
rect 6200 5300 6500 5310
rect 7400 5300 7500 5310
rect 7600 5300 7750 5310
rect 7800 5300 7900 5310
rect 8850 5300 8950 5310
rect 9000 5300 9100 5310
rect 9150 5300 9250 5310
rect 9900 5300 9990 5310
rect 1950 5290 2000 5300
rect 2900 5290 3000 5300
rect 3450 5290 3500 5300
rect 7350 5290 7700 5300
rect 7850 5290 7900 5300
rect 8600 5290 8650 5300
rect 8700 5290 8750 5300
rect 8800 5290 8950 5300
rect 9200 5290 9250 5300
rect 9700 5290 9750 5300
rect 1950 5280 2000 5290
rect 2900 5280 3000 5290
rect 3450 5280 3500 5290
rect 7350 5280 7700 5290
rect 7850 5280 7900 5290
rect 8600 5280 8650 5290
rect 8700 5280 8750 5290
rect 8800 5280 8950 5290
rect 9200 5280 9250 5290
rect 9700 5280 9750 5290
rect 1950 5270 2000 5280
rect 2900 5270 3000 5280
rect 3450 5270 3500 5280
rect 7350 5270 7700 5280
rect 7850 5270 7900 5280
rect 8600 5270 8650 5280
rect 8700 5270 8750 5280
rect 8800 5270 8950 5280
rect 9200 5270 9250 5280
rect 9700 5270 9750 5280
rect 1950 5260 2000 5270
rect 2900 5260 3000 5270
rect 3450 5260 3500 5270
rect 7350 5260 7700 5270
rect 7850 5260 7900 5270
rect 8600 5260 8650 5270
rect 8700 5260 8750 5270
rect 8800 5260 8950 5270
rect 9200 5260 9250 5270
rect 9700 5260 9750 5270
rect 1950 5250 2000 5260
rect 2900 5250 3000 5260
rect 3450 5250 3500 5260
rect 7350 5250 7700 5260
rect 7850 5250 7900 5260
rect 8600 5250 8650 5260
rect 8700 5250 8750 5260
rect 8800 5250 8950 5260
rect 9200 5250 9250 5260
rect 9700 5250 9750 5260
rect 650 5240 700 5250
rect 1950 5240 2000 5250
rect 2900 5240 3000 5250
rect 7350 5240 7450 5250
rect 7550 5240 7650 5250
rect 7850 5240 7900 5250
rect 8500 5240 8750 5250
rect 9200 5240 9250 5250
rect 9500 5240 9700 5250
rect 650 5230 700 5240
rect 1950 5230 2000 5240
rect 2900 5230 3000 5240
rect 7350 5230 7450 5240
rect 7550 5230 7650 5240
rect 7850 5230 7900 5240
rect 8500 5230 8750 5240
rect 9200 5230 9250 5240
rect 9500 5230 9700 5240
rect 650 5220 700 5230
rect 1950 5220 2000 5230
rect 2900 5220 3000 5230
rect 7350 5220 7450 5230
rect 7550 5220 7650 5230
rect 7850 5220 7900 5230
rect 8500 5220 8750 5230
rect 9200 5220 9250 5230
rect 9500 5220 9700 5230
rect 650 5210 700 5220
rect 1950 5210 2000 5220
rect 2900 5210 3000 5220
rect 7350 5210 7450 5220
rect 7550 5210 7650 5220
rect 7850 5210 7900 5220
rect 8500 5210 8750 5220
rect 9200 5210 9250 5220
rect 9500 5210 9700 5220
rect 650 5200 700 5210
rect 1950 5200 2000 5210
rect 2900 5200 3000 5210
rect 7350 5200 7450 5210
rect 7550 5200 7650 5210
rect 7850 5200 7900 5210
rect 8500 5200 8750 5210
rect 9200 5200 9250 5210
rect 9500 5200 9700 5210
rect 700 5190 750 5200
rect 1800 5190 1850 5200
rect 1950 5190 2000 5200
rect 3000 5190 3050 5200
rect 3400 5190 3450 5200
rect 7350 5190 7450 5200
rect 7550 5190 7650 5200
rect 7850 5190 7950 5200
rect 8300 5190 8600 5200
rect 9200 5190 9350 5200
rect 9650 5190 9700 5200
rect 700 5180 750 5190
rect 1800 5180 1850 5190
rect 1950 5180 2000 5190
rect 3000 5180 3050 5190
rect 3400 5180 3450 5190
rect 7350 5180 7450 5190
rect 7550 5180 7650 5190
rect 7850 5180 7950 5190
rect 8300 5180 8600 5190
rect 9200 5180 9350 5190
rect 9650 5180 9700 5190
rect 700 5170 750 5180
rect 1800 5170 1850 5180
rect 1950 5170 2000 5180
rect 3000 5170 3050 5180
rect 3400 5170 3450 5180
rect 7350 5170 7450 5180
rect 7550 5170 7650 5180
rect 7850 5170 7950 5180
rect 8300 5170 8600 5180
rect 9200 5170 9350 5180
rect 9650 5170 9700 5180
rect 700 5160 750 5170
rect 1800 5160 1850 5170
rect 1950 5160 2000 5170
rect 3000 5160 3050 5170
rect 3400 5160 3450 5170
rect 7350 5160 7450 5170
rect 7550 5160 7650 5170
rect 7850 5160 7950 5170
rect 8300 5160 8600 5170
rect 9200 5160 9350 5170
rect 9650 5160 9700 5170
rect 700 5150 750 5160
rect 1800 5150 1850 5160
rect 1950 5150 2000 5160
rect 3000 5150 3050 5160
rect 3400 5150 3450 5160
rect 7350 5150 7450 5160
rect 7550 5150 7650 5160
rect 7850 5150 7950 5160
rect 8300 5150 8600 5160
rect 9200 5150 9350 5160
rect 9650 5150 9700 5160
rect 600 5140 750 5150
rect 1800 5140 1900 5150
rect 1950 5140 2050 5150
rect 3000 5140 3050 5150
rect 7350 5140 7450 5150
rect 7850 5140 7950 5150
rect 8200 5140 8400 5150
rect 9100 5140 9250 5150
rect 9650 5140 9700 5150
rect 9950 5140 9990 5150
rect 600 5130 750 5140
rect 1800 5130 1900 5140
rect 1950 5130 2050 5140
rect 3000 5130 3050 5140
rect 7350 5130 7450 5140
rect 7850 5130 7950 5140
rect 8200 5130 8400 5140
rect 9100 5130 9250 5140
rect 9650 5130 9700 5140
rect 9950 5130 9990 5140
rect 600 5120 750 5130
rect 1800 5120 1900 5130
rect 1950 5120 2050 5130
rect 3000 5120 3050 5130
rect 7350 5120 7450 5130
rect 7850 5120 7950 5130
rect 8200 5120 8400 5130
rect 9100 5120 9250 5130
rect 9650 5120 9700 5130
rect 9950 5120 9990 5130
rect 600 5110 750 5120
rect 1800 5110 1900 5120
rect 1950 5110 2050 5120
rect 3000 5110 3050 5120
rect 7350 5110 7450 5120
rect 7850 5110 7950 5120
rect 8200 5110 8400 5120
rect 9100 5110 9250 5120
rect 9650 5110 9700 5120
rect 9950 5110 9990 5120
rect 600 5100 750 5110
rect 1800 5100 1900 5110
rect 1950 5100 2050 5110
rect 3000 5100 3050 5110
rect 7350 5100 7450 5110
rect 7850 5100 7950 5110
rect 8200 5100 8400 5110
rect 9100 5100 9250 5110
rect 9650 5100 9700 5110
rect 9950 5100 9990 5110
rect 600 5090 750 5100
rect 1750 5090 1900 5100
rect 1950 5090 2050 5100
rect 2850 5090 3050 5100
rect 3350 5090 3400 5100
rect 7350 5090 7450 5100
rect 7850 5090 7950 5100
rect 8050 5090 8150 5100
rect 8600 5090 8650 5100
rect 8900 5090 9050 5100
rect 9650 5090 9750 5100
rect 9850 5090 9900 5100
rect 600 5080 750 5090
rect 1750 5080 1900 5090
rect 1950 5080 2050 5090
rect 2850 5080 3050 5090
rect 3350 5080 3400 5090
rect 7350 5080 7450 5090
rect 7850 5080 7950 5090
rect 8050 5080 8150 5090
rect 8600 5080 8650 5090
rect 8900 5080 9050 5090
rect 9650 5080 9750 5090
rect 9850 5080 9900 5090
rect 600 5070 750 5080
rect 1750 5070 1900 5080
rect 1950 5070 2050 5080
rect 2850 5070 3050 5080
rect 3350 5070 3400 5080
rect 7350 5070 7450 5080
rect 7850 5070 7950 5080
rect 8050 5070 8150 5080
rect 8600 5070 8650 5080
rect 8900 5070 9050 5080
rect 9650 5070 9750 5080
rect 9850 5070 9900 5080
rect 600 5060 750 5070
rect 1750 5060 1900 5070
rect 1950 5060 2050 5070
rect 2850 5060 3050 5070
rect 3350 5060 3400 5070
rect 7350 5060 7450 5070
rect 7850 5060 7950 5070
rect 8050 5060 8150 5070
rect 8600 5060 8650 5070
rect 8900 5060 9050 5070
rect 9650 5060 9750 5070
rect 9850 5060 9900 5070
rect 600 5050 750 5060
rect 1750 5050 1900 5060
rect 1950 5050 2050 5060
rect 2850 5050 3050 5060
rect 3350 5050 3400 5060
rect 7350 5050 7450 5060
rect 7850 5050 7950 5060
rect 8050 5050 8150 5060
rect 8600 5050 8650 5060
rect 8900 5050 9050 5060
rect 9650 5050 9750 5060
rect 9850 5050 9900 5060
rect 450 5040 600 5050
rect 1750 5040 1900 5050
rect 2000 5040 2100 5050
rect 2900 5040 3050 5050
rect 7350 5040 7450 5050
rect 7850 5040 7950 5050
rect 8550 5040 8600 5050
rect 8700 5040 8850 5050
rect 9200 5040 9250 5050
rect 9650 5040 9700 5050
rect 450 5030 600 5040
rect 1750 5030 1900 5040
rect 2000 5030 2100 5040
rect 2900 5030 3050 5040
rect 7350 5030 7450 5040
rect 7850 5030 7950 5040
rect 8550 5030 8600 5040
rect 8700 5030 8850 5040
rect 9200 5030 9250 5040
rect 9650 5030 9700 5040
rect 450 5020 600 5030
rect 1750 5020 1900 5030
rect 2000 5020 2100 5030
rect 2900 5020 3050 5030
rect 7350 5020 7450 5030
rect 7850 5020 7950 5030
rect 8550 5020 8600 5030
rect 8700 5020 8850 5030
rect 9200 5020 9250 5030
rect 9650 5020 9700 5030
rect 450 5010 600 5020
rect 1750 5010 1900 5020
rect 2000 5010 2100 5020
rect 2900 5010 3050 5020
rect 7350 5010 7450 5020
rect 7850 5010 7950 5020
rect 8550 5010 8600 5020
rect 8700 5010 8850 5020
rect 9200 5010 9250 5020
rect 9650 5010 9700 5020
rect 450 5000 600 5010
rect 1750 5000 1900 5010
rect 2000 5000 2100 5010
rect 2900 5000 3050 5010
rect 7350 5000 7450 5010
rect 7850 5000 7950 5010
rect 8550 5000 8600 5010
rect 8700 5000 8850 5010
rect 9200 5000 9250 5010
rect 9650 5000 9700 5010
rect 450 4990 550 5000
rect 1800 4990 1850 5000
rect 2050 4990 2100 5000
rect 2800 4990 3000 5000
rect 3300 4990 3350 5000
rect 7350 4990 7400 5000
rect 7750 4990 7850 5000
rect 8550 4990 8650 5000
rect 9350 4990 9400 5000
rect 9500 4990 9600 5000
rect 450 4980 550 4990
rect 1800 4980 1850 4990
rect 2050 4980 2100 4990
rect 2800 4980 3000 4990
rect 3300 4980 3350 4990
rect 7350 4980 7400 4990
rect 7750 4980 7850 4990
rect 8550 4980 8650 4990
rect 9350 4980 9400 4990
rect 9500 4980 9600 4990
rect 450 4970 550 4980
rect 1800 4970 1850 4980
rect 2050 4970 2100 4980
rect 2800 4970 3000 4980
rect 3300 4970 3350 4980
rect 7350 4970 7400 4980
rect 7750 4970 7850 4980
rect 8550 4970 8650 4980
rect 9350 4970 9400 4980
rect 9500 4970 9600 4980
rect 450 4960 550 4970
rect 1800 4960 1850 4970
rect 2050 4960 2100 4970
rect 2800 4960 3000 4970
rect 3300 4960 3350 4970
rect 7350 4960 7400 4970
rect 7750 4960 7850 4970
rect 8550 4960 8650 4970
rect 9350 4960 9400 4970
rect 9500 4960 9600 4970
rect 450 4950 550 4960
rect 1800 4950 1850 4960
rect 2050 4950 2100 4960
rect 2800 4950 3000 4960
rect 3300 4950 3350 4960
rect 7350 4950 7400 4960
rect 7750 4950 7850 4960
rect 8550 4950 8650 4960
rect 9350 4950 9400 4960
rect 9500 4950 9600 4960
rect 450 4940 700 4950
rect 2100 4940 2200 4950
rect 2700 4940 2900 4950
rect 4200 4940 4350 4950
rect 7350 4940 7400 4950
rect 7650 4940 7700 4950
rect 8350 4940 8450 4950
rect 9350 4940 9450 4950
rect 450 4930 700 4940
rect 2100 4930 2200 4940
rect 2700 4930 2900 4940
rect 4200 4930 4350 4940
rect 7350 4930 7400 4940
rect 7650 4930 7700 4940
rect 8350 4930 8450 4940
rect 9350 4930 9450 4940
rect 450 4920 700 4930
rect 2100 4920 2200 4930
rect 2700 4920 2900 4930
rect 4200 4920 4350 4930
rect 7350 4920 7400 4930
rect 7650 4920 7700 4930
rect 8350 4920 8450 4930
rect 9350 4920 9450 4930
rect 450 4910 700 4920
rect 2100 4910 2200 4920
rect 2700 4910 2900 4920
rect 4200 4910 4350 4920
rect 7350 4910 7400 4920
rect 7650 4910 7700 4920
rect 8350 4910 8450 4920
rect 9350 4910 9450 4920
rect 450 4900 700 4910
rect 2100 4900 2200 4910
rect 2700 4900 2900 4910
rect 4200 4900 4350 4910
rect 7350 4900 7400 4910
rect 7650 4900 7700 4910
rect 8350 4900 8450 4910
rect 9350 4900 9450 4910
rect 150 4890 750 4900
rect 1050 4890 1100 4900
rect 2150 4890 2350 4900
rect 2700 4890 2850 4900
rect 3100 4890 3200 4900
rect 3250 4890 3300 4900
rect 4100 4890 4200 4900
rect 4450 4890 4550 4900
rect 4600 4890 4700 4900
rect 5600 4890 5650 4900
rect 6150 4890 6400 4900
rect 7350 4890 7400 4900
rect 8150 4890 8200 4900
rect 8400 4890 8450 4900
rect 9750 4890 9800 4900
rect 150 4880 750 4890
rect 1050 4880 1100 4890
rect 2150 4880 2350 4890
rect 2700 4880 2850 4890
rect 3100 4880 3200 4890
rect 3250 4880 3300 4890
rect 4100 4880 4200 4890
rect 4450 4880 4550 4890
rect 4600 4880 4700 4890
rect 5600 4880 5650 4890
rect 6150 4880 6400 4890
rect 7350 4880 7400 4890
rect 8150 4880 8200 4890
rect 8400 4880 8450 4890
rect 9750 4880 9800 4890
rect 150 4870 750 4880
rect 1050 4870 1100 4880
rect 2150 4870 2350 4880
rect 2700 4870 2850 4880
rect 3100 4870 3200 4880
rect 3250 4870 3300 4880
rect 4100 4870 4200 4880
rect 4450 4870 4550 4880
rect 4600 4870 4700 4880
rect 5600 4870 5650 4880
rect 6150 4870 6400 4880
rect 7350 4870 7400 4880
rect 8150 4870 8200 4880
rect 8400 4870 8450 4880
rect 9750 4870 9800 4880
rect 150 4860 750 4870
rect 1050 4860 1100 4870
rect 2150 4860 2350 4870
rect 2700 4860 2850 4870
rect 3100 4860 3200 4870
rect 3250 4860 3300 4870
rect 4100 4860 4200 4870
rect 4450 4860 4550 4870
rect 4600 4860 4700 4870
rect 5600 4860 5650 4870
rect 6150 4860 6400 4870
rect 7350 4860 7400 4870
rect 8150 4860 8200 4870
rect 8400 4860 8450 4870
rect 9750 4860 9800 4870
rect 150 4850 750 4860
rect 1050 4850 1100 4860
rect 2150 4850 2350 4860
rect 2700 4850 2850 4860
rect 3100 4850 3200 4860
rect 3250 4850 3300 4860
rect 4100 4850 4200 4860
rect 4450 4850 4550 4860
rect 4600 4850 4700 4860
rect 5600 4850 5650 4860
rect 6150 4850 6400 4860
rect 7350 4850 7400 4860
rect 8150 4850 8200 4860
rect 8400 4850 8450 4860
rect 9750 4850 9800 4860
rect 250 4840 850 4850
rect 1000 4840 1100 4850
rect 2300 4840 2350 4850
rect 2750 4840 2850 4850
rect 3050 4840 3350 4850
rect 3850 4840 3950 4850
rect 4000 4840 4050 4850
rect 4850 4840 4900 4850
rect 5550 4840 5650 4850
rect 6000 4840 6300 4850
rect 6400 4840 6450 4850
rect 7650 4840 7700 4850
rect 8400 4840 8450 4850
rect 8800 4840 9000 4850
rect 9750 4840 9800 4850
rect 250 4830 850 4840
rect 1000 4830 1100 4840
rect 2300 4830 2350 4840
rect 2750 4830 2850 4840
rect 3050 4830 3350 4840
rect 3850 4830 3950 4840
rect 4000 4830 4050 4840
rect 4850 4830 4900 4840
rect 5550 4830 5650 4840
rect 6000 4830 6300 4840
rect 6400 4830 6450 4840
rect 7650 4830 7700 4840
rect 8400 4830 8450 4840
rect 8800 4830 9000 4840
rect 9750 4830 9800 4840
rect 250 4820 850 4830
rect 1000 4820 1100 4830
rect 2300 4820 2350 4830
rect 2750 4820 2850 4830
rect 3050 4820 3350 4830
rect 3850 4820 3950 4830
rect 4000 4820 4050 4830
rect 4850 4820 4900 4830
rect 5550 4820 5650 4830
rect 6000 4820 6300 4830
rect 6400 4820 6450 4830
rect 7650 4820 7700 4830
rect 8400 4820 8450 4830
rect 8800 4820 9000 4830
rect 9750 4820 9800 4830
rect 250 4810 850 4820
rect 1000 4810 1100 4820
rect 2300 4810 2350 4820
rect 2750 4810 2850 4820
rect 3050 4810 3350 4820
rect 3850 4810 3950 4820
rect 4000 4810 4050 4820
rect 4850 4810 4900 4820
rect 5550 4810 5650 4820
rect 6000 4810 6300 4820
rect 6400 4810 6450 4820
rect 7650 4810 7700 4820
rect 8400 4810 8450 4820
rect 8800 4810 9000 4820
rect 9750 4810 9800 4820
rect 250 4800 850 4810
rect 1000 4800 1100 4810
rect 2300 4800 2350 4810
rect 2750 4800 2850 4810
rect 3050 4800 3350 4810
rect 3850 4800 3950 4810
rect 4000 4800 4050 4810
rect 4850 4800 4900 4810
rect 5550 4800 5650 4810
rect 6000 4800 6300 4810
rect 6400 4800 6450 4810
rect 7650 4800 7700 4810
rect 8400 4800 8450 4810
rect 8800 4800 9000 4810
rect 9750 4800 9800 4810
rect 200 4790 400 4800
rect 500 4790 950 4800
rect 1050 4790 1150 4800
rect 2350 4790 2400 4800
rect 2850 4790 3150 4800
rect 3200 4790 3250 4800
rect 3800 4790 3950 4800
rect 4950 4790 5000 4800
rect 5500 4790 5600 4800
rect 6450 4790 6500 4800
rect 7650 4790 7700 4800
rect 7800 4790 7850 4800
rect 8400 4790 8450 4800
rect 8550 4790 8650 4800
rect 8700 4790 8800 4800
rect 9600 4790 9750 4800
rect 9850 4790 9900 4800
rect 200 4780 400 4790
rect 500 4780 950 4790
rect 1050 4780 1150 4790
rect 2350 4780 2400 4790
rect 2850 4780 3150 4790
rect 3200 4780 3250 4790
rect 3800 4780 3950 4790
rect 4950 4780 5000 4790
rect 5500 4780 5600 4790
rect 6450 4780 6500 4790
rect 7650 4780 7700 4790
rect 7800 4780 7850 4790
rect 8400 4780 8450 4790
rect 8550 4780 8650 4790
rect 8700 4780 8800 4790
rect 9600 4780 9750 4790
rect 9850 4780 9900 4790
rect 200 4770 400 4780
rect 500 4770 950 4780
rect 1050 4770 1150 4780
rect 2350 4770 2400 4780
rect 2850 4770 3150 4780
rect 3200 4770 3250 4780
rect 3800 4770 3950 4780
rect 4950 4770 5000 4780
rect 5500 4770 5600 4780
rect 6450 4770 6500 4780
rect 7650 4770 7700 4780
rect 7800 4770 7850 4780
rect 8400 4770 8450 4780
rect 8550 4770 8650 4780
rect 8700 4770 8800 4780
rect 9600 4770 9750 4780
rect 9850 4770 9900 4780
rect 200 4760 400 4770
rect 500 4760 950 4770
rect 1050 4760 1150 4770
rect 2350 4760 2400 4770
rect 2850 4760 3150 4770
rect 3200 4760 3250 4770
rect 3800 4760 3950 4770
rect 4950 4760 5000 4770
rect 5500 4760 5600 4770
rect 6450 4760 6500 4770
rect 7650 4760 7700 4770
rect 7800 4760 7850 4770
rect 8400 4760 8450 4770
rect 8550 4760 8650 4770
rect 8700 4760 8800 4770
rect 9600 4760 9750 4770
rect 9850 4760 9900 4770
rect 200 4750 400 4760
rect 500 4750 950 4760
rect 1050 4750 1150 4760
rect 2350 4750 2400 4760
rect 2850 4750 3150 4760
rect 3200 4750 3250 4760
rect 3800 4750 3950 4760
rect 4950 4750 5000 4760
rect 5500 4750 5600 4760
rect 6450 4750 6500 4760
rect 7650 4750 7700 4760
rect 7800 4750 7850 4760
rect 8400 4750 8450 4760
rect 8550 4750 8650 4760
rect 8700 4750 8800 4760
rect 9600 4750 9750 4760
rect 9850 4750 9900 4760
rect 200 4740 450 4750
rect 550 4740 1150 4750
rect 2400 4740 2450 4750
rect 2900 4740 2950 4750
rect 3000 4740 3250 4750
rect 3800 4740 3850 4750
rect 5500 4740 5600 4750
rect 6450 4740 6550 4750
rect 7400 4740 7450 4750
rect 7600 4740 7700 4750
rect 8400 4740 8450 4750
rect 8500 4740 8600 4750
rect 9350 4740 9500 4750
rect 200 4730 450 4740
rect 550 4730 1150 4740
rect 2400 4730 2450 4740
rect 2900 4730 2950 4740
rect 3000 4730 3250 4740
rect 3800 4730 3850 4740
rect 5500 4730 5600 4740
rect 6450 4730 6550 4740
rect 7400 4730 7450 4740
rect 7600 4730 7700 4740
rect 8400 4730 8450 4740
rect 8500 4730 8600 4740
rect 9350 4730 9500 4740
rect 200 4720 450 4730
rect 550 4720 1150 4730
rect 2400 4720 2450 4730
rect 2900 4720 2950 4730
rect 3000 4720 3250 4730
rect 3800 4720 3850 4730
rect 5500 4720 5600 4730
rect 6450 4720 6550 4730
rect 7400 4720 7450 4730
rect 7600 4720 7700 4730
rect 8400 4720 8450 4730
rect 8500 4720 8600 4730
rect 9350 4720 9500 4730
rect 200 4710 450 4720
rect 550 4710 1150 4720
rect 2400 4710 2450 4720
rect 2900 4710 2950 4720
rect 3000 4710 3250 4720
rect 3800 4710 3850 4720
rect 5500 4710 5600 4720
rect 6450 4710 6550 4720
rect 7400 4710 7450 4720
rect 7600 4710 7700 4720
rect 8400 4710 8450 4720
rect 8500 4710 8600 4720
rect 9350 4710 9500 4720
rect 200 4700 450 4710
rect 550 4700 1150 4710
rect 2400 4700 2450 4710
rect 2900 4700 2950 4710
rect 3000 4700 3250 4710
rect 3800 4700 3850 4710
rect 5500 4700 5600 4710
rect 6450 4700 6550 4710
rect 7400 4700 7450 4710
rect 7600 4700 7700 4710
rect 8400 4700 8450 4710
rect 8500 4700 8600 4710
rect 9350 4700 9500 4710
rect 150 4690 550 4700
rect 750 4690 1200 4700
rect 2450 4690 2550 4700
rect 2750 4690 2800 4700
rect 2850 4690 2950 4700
rect 3000 4690 3150 4700
rect 3200 4690 3250 4700
rect 3500 4690 3550 4700
rect 5050 4690 5100 4700
rect 5500 4690 5600 4700
rect 6450 4690 6550 4700
rect 7400 4690 7500 4700
rect 8350 4690 8400 4700
rect 8450 4690 8500 4700
rect 9300 4690 9350 4700
rect 150 4680 550 4690
rect 750 4680 1200 4690
rect 2450 4680 2550 4690
rect 2750 4680 2800 4690
rect 2850 4680 2950 4690
rect 3000 4680 3150 4690
rect 3200 4680 3250 4690
rect 3500 4680 3550 4690
rect 5050 4680 5100 4690
rect 5500 4680 5600 4690
rect 6450 4680 6550 4690
rect 7400 4680 7500 4690
rect 8350 4680 8400 4690
rect 8450 4680 8500 4690
rect 9300 4680 9350 4690
rect 150 4670 550 4680
rect 750 4670 1200 4680
rect 2450 4670 2550 4680
rect 2750 4670 2800 4680
rect 2850 4670 2950 4680
rect 3000 4670 3150 4680
rect 3200 4670 3250 4680
rect 3500 4670 3550 4680
rect 5050 4670 5100 4680
rect 5500 4670 5600 4680
rect 6450 4670 6550 4680
rect 7400 4670 7500 4680
rect 8350 4670 8400 4680
rect 8450 4670 8500 4680
rect 9300 4670 9350 4680
rect 150 4660 550 4670
rect 750 4660 1200 4670
rect 2450 4660 2550 4670
rect 2750 4660 2800 4670
rect 2850 4660 2950 4670
rect 3000 4660 3150 4670
rect 3200 4660 3250 4670
rect 3500 4660 3550 4670
rect 5050 4660 5100 4670
rect 5500 4660 5600 4670
rect 6450 4660 6550 4670
rect 7400 4660 7500 4670
rect 8350 4660 8400 4670
rect 8450 4660 8500 4670
rect 9300 4660 9350 4670
rect 150 4650 550 4660
rect 750 4650 1200 4660
rect 2450 4650 2550 4660
rect 2750 4650 2800 4660
rect 2850 4650 2950 4660
rect 3000 4650 3150 4660
rect 3200 4650 3250 4660
rect 3500 4650 3550 4660
rect 5050 4650 5100 4660
rect 5500 4650 5600 4660
rect 6450 4650 6550 4660
rect 7400 4650 7500 4660
rect 8350 4650 8400 4660
rect 8450 4650 8500 4660
rect 9300 4650 9350 4660
rect 50 4640 650 4650
rect 850 4640 1200 4650
rect 2550 4640 3250 4650
rect 5100 4640 5150 4650
rect 5550 4640 5750 4650
rect 6400 4640 6550 4650
rect 7400 4640 7450 4650
rect 8100 4640 8150 4650
rect 8400 4640 8450 4650
rect 8750 4640 8800 4650
rect 50 4630 650 4640
rect 850 4630 1200 4640
rect 2550 4630 3250 4640
rect 5100 4630 5150 4640
rect 5550 4630 5750 4640
rect 6400 4630 6550 4640
rect 7400 4630 7450 4640
rect 8100 4630 8150 4640
rect 8400 4630 8450 4640
rect 8750 4630 8800 4640
rect 50 4620 650 4630
rect 850 4620 1200 4630
rect 2550 4620 3250 4630
rect 5100 4620 5150 4630
rect 5550 4620 5750 4630
rect 6400 4620 6550 4630
rect 7400 4620 7450 4630
rect 8100 4620 8150 4630
rect 8400 4620 8450 4630
rect 8750 4620 8800 4630
rect 50 4610 650 4620
rect 850 4610 1200 4620
rect 2550 4610 3250 4620
rect 5100 4610 5150 4620
rect 5550 4610 5750 4620
rect 6400 4610 6550 4620
rect 7400 4610 7450 4620
rect 8100 4610 8150 4620
rect 8400 4610 8450 4620
rect 8750 4610 8800 4620
rect 50 4600 650 4610
rect 850 4600 1200 4610
rect 2550 4600 3250 4610
rect 5100 4600 5150 4610
rect 5550 4600 5750 4610
rect 6400 4600 6550 4610
rect 7400 4600 7450 4610
rect 8100 4600 8150 4610
rect 8400 4600 8450 4610
rect 8750 4600 8800 4610
rect 0 4590 700 4600
rect 900 4590 1250 4600
rect 3000 4590 3050 4600
rect 3100 4590 3250 4600
rect 6250 4590 6350 4600
rect 6450 4590 6500 4600
rect 7400 4590 7450 4600
rect 7850 4590 7900 4600
rect 7950 4590 8000 4600
rect 8400 4590 8450 4600
rect 8800 4590 8950 4600
rect 9250 4590 9300 4600
rect 0 4580 700 4590
rect 900 4580 1250 4590
rect 3000 4580 3050 4590
rect 3100 4580 3250 4590
rect 6250 4580 6350 4590
rect 6450 4580 6500 4590
rect 7400 4580 7450 4590
rect 7850 4580 7900 4590
rect 7950 4580 8000 4590
rect 8400 4580 8450 4590
rect 8800 4580 8950 4590
rect 9250 4580 9300 4590
rect 0 4570 700 4580
rect 900 4570 1250 4580
rect 3000 4570 3050 4580
rect 3100 4570 3250 4580
rect 6250 4570 6350 4580
rect 6450 4570 6500 4580
rect 7400 4570 7450 4580
rect 7850 4570 7900 4580
rect 7950 4570 8000 4580
rect 8400 4570 8450 4580
rect 8800 4570 8950 4580
rect 9250 4570 9300 4580
rect 0 4560 700 4570
rect 900 4560 1250 4570
rect 3000 4560 3050 4570
rect 3100 4560 3250 4570
rect 6250 4560 6350 4570
rect 6450 4560 6500 4570
rect 7400 4560 7450 4570
rect 7850 4560 7900 4570
rect 7950 4560 8000 4570
rect 8400 4560 8450 4570
rect 8800 4560 8950 4570
rect 9250 4560 9300 4570
rect 0 4550 700 4560
rect 900 4550 1250 4560
rect 3000 4550 3050 4560
rect 3100 4550 3250 4560
rect 6250 4550 6350 4560
rect 6450 4550 6500 4560
rect 7400 4550 7450 4560
rect 7850 4550 7900 4560
rect 7950 4550 8000 4560
rect 8400 4550 8450 4560
rect 8800 4550 8950 4560
rect 9250 4550 9300 4560
rect 0 4540 750 4550
rect 950 4540 1200 4550
rect 2950 4540 3000 4550
rect 3050 4540 3100 4550
rect 3150 4540 3200 4550
rect 3450 4540 3500 4550
rect 3850 4540 3950 4550
rect 5200 4540 5250 4550
rect 5700 4540 5800 4550
rect 6300 4540 6350 4550
rect 6400 4540 6500 4550
rect 7550 4540 7600 4550
rect 8400 4540 8450 4550
rect 8600 4540 8700 4550
rect 9250 4540 9300 4550
rect 0 4530 750 4540
rect 950 4530 1200 4540
rect 2950 4530 3000 4540
rect 3050 4530 3100 4540
rect 3150 4530 3200 4540
rect 3450 4530 3500 4540
rect 3850 4530 3950 4540
rect 5200 4530 5250 4540
rect 5700 4530 5800 4540
rect 6300 4530 6350 4540
rect 6400 4530 6500 4540
rect 7550 4530 7600 4540
rect 8400 4530 8450 4540
rect 8600 4530 8700 4540
rect 9250 4530 9300 4540
rect 0 4520 750 4530
rect 950 4520 1200 4530
rect 2950 4520 3000 4530
rect 3050 4520 3100 4530
rect 3150 4520 3200 4530
rect 3450 4520 3500 4530
rect 3850 4520 3950 4530
rect 5200 4520 5250 4530
rect 5700 4520 5800 4530
rect 6300 4520 6350 4530
rect 6400 4520 6500 4530
rect 7550 4520 7600 4530
rect 8400 4520 8450 4530
rect 8600 4520 8700 4530
rect 9250 4520 9300 4530
rect 0 4510 750 4520
rect 950 4510 1200 4520
rect 2950 4510 3000 4520
rect 3050 4510 3100 4520
rect 3150 4510 3200 4520
rect 3450 4510 3500 4520
rect 3850 4510 3950 4520
rect 5200 4510 5250 4520
rect 5700 4510 5800 4520
rect 6300 4510 6350 4520
rect 6400 4510 6500 4520
rect 7550 4510 7600 4520
rect 8400 4510 8450 4520
rect 8600 4510 8700 4520
rect 9250 4510 9300 4520
rect 0 4500 750 4510
rect 950 4500 1200 4510
rect 2950 4500 3000 4510
rect 3050 4500 3100 4510
rect 3150 4500 3200 4510
rect 3450 4500 3500 4510
rect 3850 4500 3950 4510
rect 5200 4500 5250 4510
rect 5700 4500 5800 4510
rect 6300 4500 6350 4510
rect 6400 4500 6500 4510
rect 7550 4500 7600 4510
rect 8400 4500 8450 4510
rect 8600 4500 8700 4510
rect 9250 4500 9300 4510
rect 0 4490 650 4500
rect 1000 4490 1200 4500
rect 2800 4490 2900 4500
rect 3150 4490 3250 4500
rect 3850 4490 3950 4500
rect 6250 4490 6300 4500
rect 6350 4490 6400 4500
rect 7450 4490 7550 4500
rect 7700 4490 7750 4500
rect 8400 4490 8450 4500
rect 8850 4490 8900 4500
rect 0 4480 650 4490
rect 1000 4480 1200 4490
rect 2800 4480 2900 4490
rect 3150 4480 3250 4490
rect 3850 4480 3950 4490
rect 6250 4480 6300 4490
rect 6350 4480 6400 4490
rect 7450 4480 7550 4490
rect 7700 4480 7750 4490
rect 8400 4480 8450 4490
rect 8850 4480 8900 4490
rect 0 4470 650 4480
rect 1000 4470 1200 4480
rect 2800 4470 2900 4480
rect 3150 4470 3250 4480
rect 3850 4470 3950 4480
rect 6250 4470 6300 4480
rect 6350 4470 6400 4480
rect 7450 4470 7550 4480
rect 7700 4470 7750 4480
rect 8400 4470 8450 4480
rect 8850 4470 8900 4480
rect 0 4460 650 4470
rect 1000 4460 1200 4470
rect 2800 4460 2900 4470
rect 3150 4460 3250 4470
rect 3850 4460 3950 4470
rect 6250 4460 6300 4470
rect 6350 4460 6400 4470
rect 7450 4460 7550 4470
rect 7700 4460 7750 4470
rect 8400 4460 8450 4470
rect 8850 4460 8900 4470
rect 0 4450 650 4460
rect 1000 4450 1200 4460
rect 2800 4450 2900 4460
rect 3150 4450 3250 4460
rect 3850 4450 3950 4460
rect 6250 4450 6300 4460
rect 6350 4450 6400 4460
rect 7450 4450 7550 4460
rect 7700 4450 7750 4460
rect 8400 4450 8450 4460
rect 8850 4450 8900 4460
rect 0 4440 450 4450
rect 1050 4440 1150 4450
rect 2800 4440 2900 4450
rect 3150 4440 3200 4450
rect 3400 4440 3450 4450
rect 3850 4440 3950 4450
rect 4250 4440 4300 4450
rect 4700 4440 4750 4450
rect 5250 4440 5300 4450
rect 6200 4440 6350 4450
rect 8250 4440 8350 4450
rect 8650 4440 8750 4450
rect 8800 4440 8850 4450
rect 0 4430 450 4440
rect 1050 4430 1150 4440
rect 2800 4430 2900 4440
rect 3150 4430 3200 4440
rect 3400 4430 3450 4440
rect 3850 4430 3950 4440
rect 4250 4430 4300 4440
rect 4700 4430 4750 4440
rect 5250 4430 5300 4440
rect 6200 4430 6350 4440
rect 8250 4430 8350 4440
rect 8650 4430 8750 4440
rect 8800 4430 8850 4440
rect 0 4420 450 4430
rect 1050 4420 1150 4430
rect 2800 4420 2900 4430
rect 3150 4420 3200 4430
rect 3400 4420 3450 4430
rect 3850 4420 3950 4430
rect 4250 4420 4300 4430
rect 4700 4420 4750 4430
rect 5250 4420 5300 4430
rect 6200 4420 6350 4430
rect 8250 4420 8350 4430
rect 8650 4420 8750 4430
rect 8800 4420 8850 4430
rect 0 4410 450 4420
rect 1050 4410 1150 4420
rect 2800 4410 2900 4420
rect 3150 4410 3200 4420
rect 3400 4410 3450 4420
rect 3850 4410 3950 4420
rect 4250 4410 4300 4420
rect 4700 4410 4750 4420
rect 5250 4410 5300 4420
rect 6200 4410 6350 4420
rect 8250 4410 8350 4420
rect 8650 4410 8750 4420
rect 8800 4410 8850 4420
rect 0 4400 450 4410
rect 1050 4400 1150 4410
rect 2800 4400 2900 4410
rect 3150 4400 3200 4410
rect 3400 4400 3450 4410
rect 3850 4400 3950 4410
rect 4250 4400 4300 4410
rect 4700 4400 4750 4410
rect 5250 4400 5300 4410
rect 6200 4400 6350 4410
rect 8250 4400 8350 4410
rect 8650 4400 8750 4410
rect 8800 4400 8850 4410
rect 0 4390 250 4400
rect 2800 4390 2950 4400
rect 3100 4390 3200 4400
rect 3800 4390 3950 4400
rect 4250 4390 4350 4400
rect 4850 4390 4950 4400
rect 7750 4390 7800 4400
rect 8000 4390 8200 4400
rect 8450 4390 8550 4400
rect 8800 4390 8850 4400
rect 9200 4390 9250 4400
rect 0 4380 250 4390
rect 2800 4380 2950 4390
rect 3100 4380 3200 4390
rect 3800 4380 3950 4390
rect 4250 4380 4350 4390
rect 4850 4380 4950 4390
rect 7750 4380 7800 4390
rect 8000 4380 8200 4390
rect 8450 4380 8550 4390
rect 8800 4380 8850 4390
rect 9200 4380 9250 4390
rect 0 4370 250 4380
rect 2800 4370 2950 4380
rect 3100 4370 3200 4380
rect 3800 4370 3950 4380
rect 4250 4370 4350 4380
rect 4850 4370 4950 4380
rect 7750 4370 7800 4380
rect 8000 4370 8200 4380
rect 8450 4370 8550 4380
rect 8800 4370 8850 4380
rect 9200 4370 9250 4380
rect 0 4360 250 4370
rect 2800 4360 2950 4370
rect 3100 4360 3200 4370
rect 3800 4360 3950 4370
rect 4250 4360 4350 4370
rect 4850 4360 4950 4370
rect 7750 4360 7800 4370
rect 8000 4360 8200 4370
rect 8450 4360 8550 4370
rect 8800 4360 8850 4370
rect 9200 4360 9250 4370
rect 0 4350 250 4360
rect 2800 4350 2950 4360
rect 3100 4350 3200 4360
rect 3800 4350 3950 4360
rect 4250 4350 4350 4360
rect 4850 4350 4950 4360
rect 7750 4350 7800 4360
rect 8000 4350 8200 4360
rect 8450 4350 8550 4360
rect 8800 4350 8850 4360
rect 9200 4350 9250 4360
rect 0 4340 250 4350
rect 2800 4340 2900 4350
rect 3050 4340 3150 4350
rect 3300 4340 3400 4350
rect 4150 4340 4200 4350
rect 4250 4340 4350 4350
rect 4500 4340 4550 4350
rect 7400 4340 7450 4350
rect 7800 4340 7900 4350
rect 8150 4340 8200 4350
rect 8750 4340 8850 4350
rect 9200 4340 9250 4350
rect 0 4330 250 4340
rect 2800 4330 2900 4340
rect 3050 4330 3150 4340
rect 3300 4330 3400 4340
rect 4150 4330 4200 4340
rect 4250 4330 4350 4340
rect 4500 4330 4550 4340
rect 7400 4330 7450 4340
rect 7800 4330 7900 4340
rect 8150 4330 8200 4340
rect 8750 4330 8850 4340
rect 9200 4330 9250 4340
rect 0 4320 250 4330
rect 2800 4320 2900 4330
rect 3050 4320 3150 4330
rect 3300 4320 3400 4330
rect 4150 4320 4200 4330
rect 4250 4320 4350 4330
rect 4500 4320 4550 4330
rect 7400 4320 7450 4330
rect 7800 4320 7900 4330
rect 8150 4320 8200 4330
rect 8750 4320 8850 4330
rect 9200 4320 9250 4330
rect 0 4310 250 4320
rect 2800 4310 2900 4320
rect 3050 4310 3150 4320
rect 3300 4310 3400 4320
rect 4150 4310 4200 4320
rect 4250 4310 4350 4320
rect 4500 4310 4550 4320
rect 7400 4310 7450 4320
rect 7800 4310 7900 4320
rect 8150 4310 8200 4320
rect 8750 4310 8850 4320
rect 9200 4310 9250 4320
rect 0 4300 250 4310
rect 2800 4300 2900 4310
rect 3050 4300 3150 4310
rect 3300 4300 3400 4310
rect 4150 4300 4200 4310
rect 4250 4300 4350 4310
rect 4500 4300 4550 4310
rect 7400 4300 7450 4310
rect 7800 4300 7900 4310
rect 8150 4300 8200 4310
rect 8750 4300 8850 4310
rect 9200 4300 9250 4310
rect 0 4290 100 4300
rect 2800 4290 2900 4300
rect 3250 4290 3300 4300
rect 4100 4290 4150 4300
rect 4450 4290 4500 4300
rect 4950 4290 5000 4300
rect 5300 4290 5350 4300
rect 7300 4290 7450 4300
rect 8150 4290 8200 4300
rect 9200 4290 9250 4300
rect 9350 4290 9400 4300
rect 0 4280 100 4290
rect 2800 4280 2900 4290
rect 3250 4280 3300 4290
rect 4100 4280 4150 4290
rect 4450 4280 4500 4290
rect 4950 4280 5000 4290
rect 5300 4280 5350 4290
rect 7300 4280 7450 4290
rect 8150 4280 8200 4290
rect 9200 4280 9250 4290
rect 9350 4280 9400 4290
rect 0 4270 100 4280
rect 2800 4270 2900 4280
rect 3250 4270 3300 4280
rect 4100 4270 4150 4280
rect 4450 4270 4500 4280
rect 4950 4270 5000 4280
rect 5300 4270 5350 4280
rect 7300 4270 7450 4280
rect 8150 4270 8200 4280
rect 9200 4270 9250 4280
rect 9350 4270 9400 4280
rect 0 4260 100 4270
rect 2800 4260 2900 4270
rect 3250 4260 3300 4270
rect 4100 4260 4150 4270
rect 4450 4260 4500 4270
rect 4950 4260 5000 4270
rect 5300 4260 5350 4270
rect 7300 4260 7450 4270
rect 8150 4260 8200 4270
rect 9200 4260 9250 4270
rect 9350 4260 9400 4270
rect 0 4250 100 4260
rect 2800 4250 2900 4260
rect 3250 4250 3300 4260
rect 4100 4250 4150 4260
rect 4450 4250 4500 4260
rect 4950 4250 5000 4260
rect 5300 4250 5350 4260
rect 7300 4250 7450 4260
rect 8150 4250 8200 4260
rect 9200 4250 9250 4260
rect 9350 4250 9400 4260
rect 0 4240 150 4250
rect 2750 4240 2900 4250
rect 2950 4240 3000 4250
rect 3250 4240 3300 4250
rect 4400 4240 4450 4250
rect 5000 4240 5050 4250
rect 8150 4240 8200 4250
rect 8400 4240 8450 4250
rect 8500 4240 8550 4250
rect 0 4230 150 4240
rect 2750 4230 2900 4240
rect 2950 4230 3000 4240
rect 3250 4230 3300 4240
rect 4400 4230 4450 4240
rect 5000 4230 5050 4240
rect 8150 4230 8200 4240
rect 8400 4230 8450 4240
rect 8500 4230 8550 4240
rect 0 4220 150 4230
rect 2750 4220 2900 4230
rect 2950 4220 3000 4230
rect 3250 4220 3300 4230
rect 4400 4220 4450 4230
rect 5000 4220 5050 4230
rect 8150 4220 8200 4230
rect 8400 4220 8450 4230
rect 8500 4220 8550 4230
rect 0 4210 150 4220
rect 2750 4210 2900 4220
rect 2950 4210 3000 4220
rect 3250 4210 3300 4220
rect 4400 4210 4450 4220
rect 5000 4210 5050 4220
rect 8150 4210 8200 4220
rect 8400 4210 8450 4220
rect 8500 4210 8550 4220
rect 0 4200 150 4210
rect 2750 4200 2900 4210
rect 2950 4200 3000 4210
rect 3250 4200 3300 4210
rect 4400 4200 4450 4210
rect 5000 4200 5050 4210
rect 8150 4200 8200 4210
rect 8400 4200 8450 4210
rect 8500 4200 8550 4210
rect 0 4190 150 4200
rect 2550 4190 2850 4200
rect 2950 4190 3000 4200
rect 3250 4190 3300 4200
rect 4050 4190 4100 4200
rect 5350 4190 5400 4200
rect 8750 4190 8800 4200
rect 0 4180 150 4190
rect 2550 4180 2850 4190
rect 2950 4180 3000 4190
rect 3250 4180 3300 4190
rect 4050 4180 4100 4190
rect 5350 4180 5400 4190
rect 8750 4180 8800 4190
rect 0 4170 150 4180
rect 2550 4170 2850 4180
rect 2950 4170 3000 4180
rect 3250 4170 3300 4180
rect 4050 4170 4100 4180
rect 5350 4170 5400 4180
rect 8750 4170 8800 4180
rect 0 4160 150 4170
rect 2550 4160 2850 4170
rect 2950 4160 3000 4170
rect 3250 4160 3300 4170
rect 4050 4160 4100 4170
rect 5350 4160 5400 4170
rect 8750 4160 8800 4170
rect 0 4150 150 4160
rect 2550 4150 2850 4160
rect 2950 4150 3000 4160
rect 3250 4150 3300 4160
rect 4050 4150 4100 4160
rect 5350 4150 5400 4160
rect 8750 4150 8800 4160
rect 50 4140 150 4150
rect 2600 4140 2850 4150
rect 3300 4140 3350 4150
rect 5100 4140 5150 4150
rect 5550 4140 5600 4150
rect 7250 4140 7350 4150
rect 7500 4140 7550 4150
rect 8750 4140 8800 4150
rect 50 4130 150 4140
rect 2600 4130 2850 4140
rect 3300 4130 3350 4140
rect 5100 4130 5150 4140
rect 5550 4130 5600 4140
rect 7250 4130 7350 4140
rect 7500 4130 7550 4140
rect 8750 4130 8800 4140
rect 50 4120 150 4130
rect 2600 4120 2850 4130
rect 3300 4120 3350 4130
rect 5100 4120 5150 4130
rect 5550 4120 5600 4130
rect 7250 4120 7350 4130
rect 7500 4120 7550 4130
rect 8750 4120 8800 4130
rect 50 4110 150 4120
rect 2600 4110 2850 4120
rect 3300 4110 3350 4120
rect 5100 4110 5150 4120
rect 5550 4110 5600 4120
rect 7250 4110 7350 4120
rect 7500 4110 7550 4120
rect 8750 4110 8800 4120
rect 50 4100 150 4110
rect 2600 4100 2850 4110
rect 3300 4100 3350 4110
rect 5100 4100 5150 4110
rect 5550 4100 5600 4110
rect 7250 4100 7350 4110
rect 7500 4100 7550 4110
rect 8750 4100 8800 4110
rect 100 4090 150 4100
rect 2600 4090 2850 4100
rect 2900 4090 2950 4100
rect 4000 4090 4050 4100
rect 4650 4090 4800 4100
rect 5100 4090 5150 4100
rect 5600 4090 5650 4100
rect 7250 4090 7300 4100
rect 7450 4090 7600 4100
rect 7650 4090 7700 4100
rect 8550 4090 8700 4100
rect 100 4080 150 4090
rect 2600 4080 2850 4090
rect 2900 4080 2950 4090
rect 4000 4080 4050 4090
rect 4650 4080 4800 4090
rect 5100 4080 5150 4090
rect 5600 4080 5650 4090
rect 7250 4080 7300 4090
rect 7450 4080 7600 4090
rect 7650 4080 7700 4090
rect 8550 4080 8700 4090
rect 100 4070 150 4080
rect 2600 4070 2850 4080
rect 2900 4070 2950 4080
rect 4000 4070 4050 4080
rect 4650 4070 4800 4080
rect 5100 4070 5150 4080
rect 5600 4070 5650 4080
rect 7250 4070 7300 4080
rect 7450 4070 7600 4080
rect 7650 4070 7700 4080
rect 8550 4070 8700 4080
rect 100 4060 150 4070
rect 2600 4060 2850 4070
rect 2900 4060 2950 4070
rect 4000 4060 4050 4070
rect 4650 4060 4800 4070
rect 5100 4060 5150 4070
rect 5600 4060 5650 4070
rect 7250 4060 7300 4070
rect 7450 4060 7600 4070
rect 7650 4060 7700 4070
rect 8550 4060 8700 4070
rect 100 4050 150 4060
rect 2600 4050 2850 4060
rect 2900 4050 2950 4060
rect 4000 4050 4050 4060
rect 4650 4050 4800 4060
rect 5100 4050 5150 4060
rect 5600 4050 5650 4060
rect 7250 4050 7300 4060
rect 7450 4050 7600 4060
rect 7650 4050 7700 4060
rect 8550 4050 8700 4060
rect 2600 4040 2750 4050
rect 2800 4040 2950 4050
rect 4650 4040 4700 4050
rect 5150 4040 5200 4050
rect 5350 4040 5400 4050
rect 5650 4040 5700 4050
rect 7600 4040 7850 4050
rect 8300 4040 8350 4050
rect 8700 4040 8750 4050
rect 2600 4030 2750 4040
rect 2800 4030 2950 4040
rect 4650 4030 4700 4040
rect 5150 4030 5200 4040
rect 5350 4030 5400 4040
rect 5650 4030 5700 4040
rect 7600 4030 7850 4040
rect 8300 4030 8350 4040
rect 8700 4030 8750 4040
rect 2600 4020 2750 4030
rect 2800 4020 2950 4030
rect 4650 4020 4700 4030
rect 5150 4020 5200 4030
rect 5350 4020 5400 4030
rect 5650 4020 5700 4030
rect 7600 4020 7850 4030
rect 8300 4020 8350 4030
rect 8700 4020 8750 4030
rect 2600 4010 2750 4020
rect 2800 4010 2950 4020
rect 4650 4010 4700 4020
rect 5150 4010 5200 4020
rect 5350 4010 5400 4020
rect 5650 4010 5700 4020
rect 7600 4010 7850 4020
rect 8300 4010 8350 4020
rect 8700 4010 8750 4020
rect 2600 4000 2750 4010
rect 2800 4000 2950 4010
rect 4650 4000 4700 4010
rect 5150 4000 5200 4010
rect 5350 4000 5400 4010
rect 5650 4000 5700 4010
rect 7600 4000 7850 4010
rect 8300 4000 8350 4010
rect 8700 4000 8750 4010
rect 2600 3990 2900 4000
rect 3000 3990 3050 4000
rect 3900 3990 3950 4000
rect 5350 3990 5400 4000
rect 5500 3990 5550 4000
rect 5750 3990 5800 4000
rect 7750 3990 7850 4000
rect 7900 3990 7950 4000
rect 8100 3990 8200 4000
rect 2600 3980 2900 3990
rect 3000 3980 3050 3990
rect 3900 3980 3950 3990
rect 5350 3980 5400 3990
rect 5500 3980 5550 3990
rect 5750 3980 5800 3990
rect 7750 3980 7850 3990
rect 7900 3980 7950 3990
rect 8100 3980 8200 3990
rect 2600 3970 2900 3980
rect 3000 3970 3050 3980
rect 3900 3970 3950 3980
rect 5350 3970 5400 3980
rect 5500 3970 5550 3980
rect 5750 3970 5800 3980
rect 7750 3970 7850 3980
rect 7900 3970 7950 3980
rect 8100 3970 8200 3980
rect 2600 3960 2900 3970
rect 3000 3960 3050 3970
rect 3900 3960 3950 3970
rect 5350 3960 5400 3970
rect 5500 3960 5550 3970
rect 5750 3960 5800 3970
rect 7750 3960 7850 3970
rect 7900 3960 7950 3970
rect 8100 3960 8200 3970
rect 2600 3950 2900 3960
rect 3000 3950 3050 3960
rect 3900 3950 3950 3960
rect 5350 3950 5400 3960
rect 5500 3950 5550 3960
rect 5750 3950 5800 3960
rect 7750 3950 7850 3960
rect 7900 3950 7950 3960
rect 8100 3950 8200 3960
rect 2600 3940 2850 3950
rect 3850 3940 3900 3950
rect 5200 3940 5250 3950
rect 5400 3940 5500 3950
rect 5900 3940 6300 3950
rect 7850 3940 7950 3950
rect 2600 3930 2850 3940
rect 3850 3930 3900 3940
rect 5200 3930 5250 3940
rect 5400 3930 5500 3940
rect 5900 3930 6300 3940
rect 7850 3930 7950 3940
rect 2600 3920 2850 3930
rect 3850 3920 3900 3930
rect 5200 3920 5250 3930
rect 5400 3920 5500 3930
rect 5900 3920 6300 3930
rect 7850 3920 7950 3930
rect 2600 3910 2850 3920
rect 3850 3910 3900 3920
rect 5200 3910 5250 3920
rect 5400 3910 5500 3920
rect 5900 3910 6300 3920
rect 7850 3910 7950 3920
rect 2600 3900 2850 3910
rect 3850 3900 3900 3910
rect 5200 3900 5250 3910
rect 5400 3900 5500 3910
rect 5900 3900 6300 3910
rect 7850 3900 7950 3910
rect 2550 3890 2850 3900
rect 3300 3890 3350 3900
rect 4150 3890 4250 3900
rect 5250 3890 5300 3900
rect 6000 3890 6300 3900
rect 7150 3890 7200 3900
rect 7950 3890 8000 3900
rect 8150 3890 8200 3900
rect 2550 3880 2850 3890
rect 3300 3880 3350 3890
rect 4150 3880 4250 3890
rect 5250 3880 5300 3890
rect 6000 3880 6300 3890
rect 7150 3880 7200 3890
rect 7950 3880 8000 3890
rect 8150 3880 8200 3890
rect 2550 3870 2850 3880
rect 3300 3870 3350 3880
rect 4150 3870 4250 3880
rect 5250 3870 5300 3880
rect 6000 3870 6300 3880
rect 7150 3870 7200 3880
rect 7950 3870 8000 3880
rect 8150 3870 8200 3880
rect 2550 3860 2850 3870
rect 3300 3860 3350 3870
rect 4150 3860 4250 3870
rect 5250 3860 5300 3870
rect 6000 3860 6300 3870
rect 7150 3860 7200 3870
rect 7950 3860 8000 3870
rect 8150 3860 8200 3870
rect 2550 3850 2850 3860
rect 3300 3850 3350 3860
rect 4150 3850 4250 3860
rect 5250 3850 5300 3860
rect 6000 3850 6300 3860
rect 7150 3850 7200 3860
rect 7950 3850 8000 3860
rect 8150 3850 8200 3860
rect 2400 3840 2450 3850
rect 2550 3840 2850 3850
rect 4100 3840 4150 3850
rect 4200 3840 4250 3850
rect 5250 3840 5300 3850
rect 5950 3840 6300 3850
rect 8000 3840 8200 3850
rect 9650 3840 9700 3850
rect 2400 3830 2450 3840
rect 2550 3830 2850 3840
rect 4100 3830 4150 3840
rect 4200 3830 4250 3840
rect 5250 3830 5300 3840
rect 5950 3830 6300 3840
rect 8000 3830 8200 3840
rect 9650 3830 9700 3840
rect 2400 3820 2450 3830
rect 2550 3820 2850 3830
rect 4100 3820 4150 3830
rect 4200 3820 4250 3830
rect 5250 3820 5300 3830
rect 5950 3820 6300 3830
rect 8000 3820 8200 3830
rect 9650 3820 9700 3830
rect 2400 3810 2450 3820
rect 2550 3810 2850 3820
rect 4100 3810 4150 3820
rect 4200 3810 4250 3820
rect 5250 3810 5300 3820
rect 5950 3810 6300 3820
rect 8000 3810 8200 3820
rect 9650 3810 9700 3820
rect 2400 3800 2450 3810
rect 2550 3800 2850 3810
rect 4100 3800 4150 3810
rect 4200 3800 4250 3810
rect 5250 3800 5300 3810
rect 5950 3800 6300 3810
rect 8000 3800 8200 3810
rect 9650 3800 9700 3810
rect 2550 3790 2900 3800
rect 3300 3790 3350 3800
rect 4050 3790 4100 3800
rect 6000 3790 6300 3800
rect 2550 3780 2900 3790
rect 3300 3780 3350 3790
rect 4050 3780 4100 3790
rect 6000 3780 6300 3790
rect 2550 3770 2900 3780
rect 3300 3770 3350 3780
rect 4050 3770 4100 3780
rect 6000 3770 6300 3780
rect 2550 3760 2900 3770
rect 3300 3760 3350 3770
rect 4050 3760 4100 3770
rect 6000 3760 6300 3770
rect 2550 3750 2900 3760
rect 3300 3750 3350 3760
rect 4050 3750 4100 3760
rect 6000 3750 6300 3760
rect 1600 3740 1700 3750
rect 2700 3740 2850 3750
rect 3300 3740 3350 3750
rect 5300 3740 5350 3750
rect 6050 3740 6400 3750
rect 7050 3740 7100 3750
rect 1600 3730 1700 3740
rect 2700 3730 2850 3740
rect 3300 3730 3350 3740
rect 5300 3730 5350 3740
rect 6050 3730 6400 3740
rect 7050 3730 7100 3740
rect 1600 3720 1700 3730
rect 2700 3720 2850 3730
rect 3300 3720 3350 3730
rect 5300 3720 5350 3730
rect 6050 3720 6400 3730
rect 7050 3720 7100 3730
rect 1600 3710 1700 3720
rect 2700 3710 2850 3720
rect 3300 3710 3350 3720
rect 5300 3710 5350 3720
rect 6050 3710 6400 3720
rect 7050 3710 7100 3720
rect 1600 3700 1700 3710
rect 2700 3700 2850 3710
rect 3300 3700 3350 3710
rect 5300 3700 5350 3710
rect 6050 3700 6400 3710
rect 7050 3700 7100 3710
rect 0 3690 50 3700
rect 1600 3690 1700 3700
rect 2850 3690 3050 3700
rect 3850 3690 3900 3700
rect 5300 3690 5350 3700
rect 6050 3690 6450 3700
rect 8150 3690 8200 3700
rect 0 3680 50 3690
rect 1600 3680 1700 3690
rect 2850 3680 3050 3690
rect 3850 3680 3900 3690
rect 5300 3680 5350 3690
rect 6050 3680 6450 3690
rect 8150 3680 8200 3690
rect 0 3670 50 3680
rect 1600 3670 1700 3680
rect 2850 3670 3050 3680
rect 3850 3670 3900 3680
rect 5300 3670 5350 3680
rect 6050 3670 6450 3680
rect 8150 3670 8200 3680
rect 0 3660 50 3670
rect 1600 3660 1700 3670
rect 2850 3660 3050 3670
rect 3850 3660 3900 3670
rect 5300 3660 5350 3670
rect 6050 3660 6450 3670
rect 8150 3660 8200 3670
rect 0 3650 50 3660
rect 1600 3650 1700 3660
rect 2850 3650 3050 3660
rect 3850 3650 3900 3660
rect 5300 3650 5350 3660
rect 6050 3650 6450 3660
rect 8150 3650 8200 3660
rect 3050 3640 3150 3650
rect 3350 3640 3400 3650
rect 6150 3640 6400 3650
rect 8400 3640 8500 3650
rect 3050 3630 3150 3640
rect 3350 3630 3400 3640
rect 6150 3630 6400 3640
rect 8400 3630 8500 3640
rect 3050 3620 3150 3630
rect 3350 3620 3400 3630
rect 6150 3620 6400 3630
rect 8400 3620 8500 3630
rect 3050 3610 3150 3620
rect 3350 3610 3400 3620
rect 6150 3610 6400 3620
rect 8400 3610 8500 3620
rect 3050 3600 3150 3610
rect 3350 3600 3400 3610
rect 6150 3600 6400 3610
rect 8400 3600 8500 3610
rect 3200 3590 3250 3600
rect 3400 3590 3450 3600
rect 6150 3590 6350 3600
rect 6950 3590 7000 3600
rect 3200 3580 3250 3590
rect 3400 3580 3450 3590
rect 6150 3580 6350 3590
rect 6950 3580 7000 3590
rect 3200 3570 3250 3580
rect 3400 3570 3450 3580
rect 6150 3570 6350 3580
rect 6950 3570 7000 3580
rect 3200 3560 3250 3570
rect 3400 3560 3450 3570
rect 6150 3560 6350 3570
rect 6950 3560 7000 3570
rect 3200 3550 3250 3560
rect 3400 3550 3450 3560
rect 6150 3550 6350 3560
rect 6950 3550 7000 3560
rect 1400 3540 1500 3550
rect 2400 3540 2500 3550
rect 2600 3540 2750 3550
rect 5350 3540 5400 3550
rect 6150 3540 6350 3550
rect 6900 3540 6950 3550
rect 1400 3530 1500 3540
rect 2400 3530 2500 3540
rect 2600 3530 2750 3540
rect 5350 3530 5400 3540
rect 6150 3530 6350 3540
rect 6900 3530 6950 3540
rect 1400 3520 1500 3530
rect 2400 3520 2500 3530
rect 2600 3520 2750 3530
rect 5350 3520 5400 3530
rect 6150 3520 6350 3530
rect 6900 3520 6950 3530
rect 1400 3510 1500 3520
rect 2400 3510 2500 3520
rect 2600 3510 2750 3520
rect 5350 3510 5400 3520
rect 6150 3510 6350 3520
rect 6900 3510 6950 3520
rect 1400 3500 1500 3510
rect 2400 3500 2500 3510
rect 2600 3500 2750 3510
rect 5350 3500 5400 3510
rect 6150 3500 6350 3510
rect 6900 3500 6950 3510
rect 1400 3490 1450 3500
rect 2250 3490 2300 3500
rect 2850 3490 2900 3500
rect 3300 3490 3350 3500
rect 3900 3490 3950 3500
rect 5350 3490 5400 3500
rect 6150 3490 6300 3500
rect 6850 3490 6900 3500
rect 8350 3490 8400 3500
rect 1400 3480 1450 3490
rect 2250 3480 2300 3490
rect 2850 3480 2900 3490
rect 3300 3480 3350 3490
rect 3900 3480 3950 3490
rect 5350 3480 5400 3490
rect 6150 3480 6300 3490
rect 6850 3480 6900 3490
rect 8350 3480 8400 3490
rect 1400 3470 1450 3480
rect 2250 3470 2300 3480
rect 2850 3470 2900 3480
rect 3300 3470 3350 3480
rect 3900 3470 3950 3480
rect 5350 3470 5400 3480
rect 6150 3470 6300 3480
rect 6850 3470 6900 3480
rect 8350 3470 8400 3480
rect 1400 3460 1450 3470
rect 2250 3460 2300 3470
rect 2850 3460 2900 3470
rect 3300 3460 3350 3470
rect 3900 3460 3950 3470
rect 5350 3460 5400 3470
rect 6150 3460 6300 3470
rect 6850 3460 6900 3470
rect 8350 3460 8400 3470
rect 1400 3450 1450 3460
rect 2250 3450 2300 3460
rect 2850 3450 2900 3460
rect 3300 3450 3350 3460
rect 3900 3450 3950 3460
rect 5350 3450 5400 3460
rect 6150 3450 6300 3460
rect 6850 3450 6900 3460
rect 8350 3450 8400 3460
rect 1350 3440 1450 3450
rect 3000 3440 3050 3450
rect 3350 3440 3450 3450
rect 3900 3440 3950 3450
rect 4500 3440 4600 3450
rect 5850 3440 6050 3450
rect 6100 3440 6200 3450
rect 6800 3440 6850 3450
rect 8400 3440 8500 3450
rect 1350 3430 1450 3440
rect 3000 3430 3050 3440
rect 3350 3430 3450 3440
rect 3900 3430 3950 3440
rect 4500 3430 4600 3440
rect 5850 3430 6050 3440
rect 6100 3430 6200 3440
rect 6800 3430 6850 3440
rect 8400 3430 8500 3440
rect 1350 3420 1450 3430
rect 3000 3420 3050 3430
rect 3350 3420 3450 3430
rect 3900 3420 3950 3430
rect 4500 3420 4600 3430
rect 5850 3420 6050 3430
rect 6100 3420 6200 3430
rect 6800 3420 6850 3430
rect 8400 3420 8500 3430
rect 1350 3410 1450 3420
rect 3000 3410 3050 3420
rect 3350 3410 3450 3420
rect 3900 3410 3950 3420
rect 4500 3410 4600 3420
rect 5850 3410 6050 3420
rect 6100 3410 6200 3420
rect 6800 3410 6850 3420
rect 8400 3410 8500 3420
rect 1350 3400 1450 3410
rect 3000 3400 3050 3410
rect 3350 3400 3450 3410
rect 3900 3400 3950 3410
rect 4500 3400 4600 3410
rect 5850 3400 6050 3410
rect 6100 3400 6200 3410
rect 6800 3400 6850 3410
rect 8400 3400 8500 3410
rect 1350 3390 1450 3400
rect 2100 3390 2150 3400
rect 3450 3390 3500 3400
rect 4800 3390 4850 3400
rect 5650 3390 5750 3400
rect 5850 3390 6050 3400
rect 6100 3390 6150 3400
rect 6750 3390 6800 3400
rect 8450 3390 8500 3400
rect 1350 3380 1450 3390
rect 2100 3380 2150 3390
rect 3450 3380 3500 3390
rect 4800 3380 4850 3390
rect 5650 3380 5750 3390
rect 5850 3380 6050 3390
rect 6100 3380 6150 3390
rect 6750 3380 6800 3390
rect 8450 3380 8500 3390
rect 1350 3370 1450 3380
rect 2100 3370 2150 3380
rect 3450 3370 3500 3380
rect 4800 3370 4850 3380
rect 5650 3370 5750 3380
rect 5850 3370 6050 3380
rect 6100 3370 6150 3380
rect 6750 3370 6800 3380
rect 8450 3370 8500 3380
rect 1350 3360 1450 3370
rect 2100 3360 2150 3370
rect 3450 3360 3500 3370
rect 4800 3360 4850 3370
rect 5650 3360 5750 3370
rect 5850 3360 6050 3370
rect 6100 3360 6150 3370
rect 6750 3360 6800 3370
rect 8450 3360 8500 3370
rect 1350 3350 1450 3360
rect 2100 3350 2150 3360
rect 3450 3350 3500 3360
rect 4800 3350 4850 3360
rect 5650 3350 5750 3360
rect 5850 3350 6050 3360
rect 6100 3350 6150 3360
rect 6750 3350 6800 3360
rect 8450 3350 8500 3360
rect 1300 3340 1400 3350
rect 3450 3340 3500 3350
rect 3600 3340 3650 3350
rect 3950 3340 4000 3350
rect 4250 3340 4300 3350
rect 4700 3340 4750 3350
rect 5600 3340 6150 3350
rect 6700 3340 6750 3350
rect 1300 3330 1400 3340
rect 3450 3330 3500 3340
rect 3600 3330 3650 3340
rect 3950 3330 4000 3340
rect 4250 3330 4300 3340
rect 4700 3330 4750 3340
rect 5600 3330 6150 3340
rect 6700 3330 6750 3340
rect 1300 3320 1400 3330
rect 3450 3320 3500 3330
rect 3600 3320 3650 3330
rect 3950 3320 4000 3330
rect 4250 3320 4300 3330
rect 4700 3320 4750 3330
rect 5600 3320 6150 3330
rect 6700 3320 6750 3330
rect 1300 3310 1400 3320
rect 3450 3310 3500 3320
rect 3600 3310 3650 3320
rect 3950 3310 4000 3320
rect 4250 3310 4300 3320
rect 4700 3310 4750 3320
rect 5600 3310 6150 3320
rect 6700 3310 6750 3320
rect 1300 3300 1400 3310
rect 3450 3300 3500 3310
rect 3600 3300 3650 3310
rect 3950 3300 4000 3310
rect 4250 3300 4300 3310
rect 4700 3300 4750 3310
rect 5600 3300 6150 3310
rect 6700 3300 6750 3310
rect 1300 3290 1400 3300
rect 2050 3290 2100 3300
rect 3150 3290 3200 3300
rect 3500 3290 3550 3300
rect 3600 3290 3650 3300
rect 4000 3290 4050 3300
rect 4250 3290 4300 3300
rect 4550 3290 4650 3300
rect 5300 3290 5350 3300
rect 5600 3290 6150 3300
rect 6650 3290 6700 3300
rect 8400 3290 8450 3300
rect 1300 3280 1400 3290
rect 2050 3280 2100 3290
rect 3150 3280 3200 3290
rect 3500 3280 3550 3290
rect 3600 3280 3650 3290
rect 4000 3280 4050 3290
rect 4250 3280 4300 3290
rect 4550 3280 4650 3290
rect 5300 3280 5350 3290
rect 5600 3280 6150 3290
rect 6650 3280 6700 3290
rect 8400 3280 8450 3290
rect 1300 3270 1400 3280
rect 2050 3270 2100 3280
rect 3150 3270 3200 3280
rect 3500 3270 3550 3280
rect 3600 3270 3650 3280
rect 4000 3270 4050 3280
rect 4250 3270 4300 3280
rect 4550 3270 4650 3280
rect 5300 3270 5350 3280
rect 5600 3270 6150 3280
rect 6650 3270 6700 3280
rect 8400 3270 8450 3280
rect 1300 3260 1400 3270
rect 2050 3260 2100 3270
rect 3150 3260 3200 3270
rect 3500 3260 3550 3270
rect 3600 3260 3650 3270
rect 4000 3260 4050 3270
rect 4250 3260 4300 3270
rect 4550 3260 4650 3270
rect 5300 3260 5350 3270
rect 5600 3260 6150 3270
rect 6650 3260 6700 3270
rect 8400 3260 8450 3270
rect 1300 3250 1400 3260
rect 2050 3250 2100 3260
rect 3150 3250 3200 3260
rect 3500 3250 3550 3260
rect 3600 3250 3650 3260
rect 4000 3250 4050 3260
rect 4250 3250 4300 3260
rect 4550 3250 4650 3260
rect 5300 3250 5350 3260
rect 5600 3250 6150 3260
rect 6650 3250 6700 3260
rect 8400 3250 8450 3260
rect 1300 3240 1400 3250
rect 4050 3240 4100 3250
rect 4350 3240 4600 3250
rect 5300 3240 5350 3250
rect 5650 3240 6200 3250
rect 6550 3240 6600 3250
rect 6650 3240 6700 3250
rect 1300 3230 1400 3240
rect 4050 3230 4100 3240
rect 4350 3230 4600 3240
rect 5300 3230 5350 3240
rect 5650 3230 6200 3240
rect 6550 3230 6600 3240
rect 6650 3230 6700 3240
rect 1300 3220 1400 3230
rect 4050 3220 4100 3230
rect 4350 3220 4600 3230
rect 5300 3220 5350 3230
rect 5650 3220 6200 3230
rect 6550 3220 6600 3230
rect 6650 3220 6700 3230
rect 1300 3210 1400 3220
rect 4050 3210 4100 3220
rect 4350 3210 4600 3220
rect 5300 3210 5350 3220
rect 5650 3210 6200 3220
rect 6550 3210 6600 3220
rect 6650 3210 6700 3220
rect 1300 3200 1400 3210
rect 4050 3200 4100 3210
rect 4350 3200 4600 3210
rect 5300 3200 5350 3210
rect 5650 3200 6200 3210
rect 6550 3200 6600 3210
rect 6650 3200 6700 3210
rect 1250 3190 1350 3200
rect 2000 3190 2050 3200
rect 4050 3190 4150 3200
rect 4400 3190 4500 3200
rect 5700 3190 6200 3200
rect 6400 3190 6500 3200
rect 6550 3190 6600 3200
rect 6650 3190 6700 3200
rect 8350 3190 8400 3200
rect 9100 3190 9200 3200
rect 1250 3180 1350 3190
rect 2000 3180 2050 3190
rect 4050 3180 4150 3190
rect 4400 3180 4500 3190
rect 5700 3180 6200 3190
rect 6400 3180 6500 3190
rect 6550 3180 6600 3190
rect 6650 3180 6700 3190
rect 8350 3180 8400 3190
rect 9100 3180 9200 3190
rect 1250 3170 1350 3180
rect 2000 3170 2050 3180
rect 4050 3170 4150 3180
rect 4400 3170 4500 3180
rect 5700 3170 6200 3180
rect 6400 3170 6500 3180
rect 6550 3170 6600 3180
rect 6650 3170 6700 3180
rect 8350 3170 8400 3180
rect 9100 3170 9200 3180
rect 1250 3160 1350 3170
rect 2000 3160 2050 3170
rect 4050 3160 4150 3170
rect 4400 3160 4500 3170
rect 5700 3160 6200 3170
rect 6400 3160 6500 3170
rect 6550 3160 6600 3170
rect 6650 3160 6700 3170
rect 8350 3160 8400 3170
rect 9100 3160 9200 3170
rect 1250 3150 1350 3160
rect 2000 3150 2050 3160
rect 4050 3150 4150 3160
rect 4400 3150 4500 3160
rect 5700 3150 6200 3160
rect 6400 3150 6500 3160
rect 6550 3150 6600 3160
rect 6650 3150 6700 3160
rect 8350 3150 8400 3160
rect 9100 3150 9200 3160
rect 1250 3140 1350 3150
rect 2000 3140 2050 3150
rect 3200 3140 3250 3150
rect 3750 3140 4000 3150
rect 4050 3140 4150 3150
rect 5800 3140 6350 3150
rect 6550 3140 6650 3150
rect 9100 3140 9150 3150
rect 1250 3130 1350 3140
rect 2000 3130 2050 3140
rect 3200 3130 3250 3140
rect 3750 3130 4000 3140
rect 4050 3130 4150 3140
rect 5800 3130 6350 3140
rect 6550 3130 6650 3140
rect 9100 3130 9150 3140
rect 1250 3120 1350 3130
rect 2000 3120 2050 3130
rect 3200 3120 3250 3130
rect 3750 3120 4000 3130
rect 4050 3120 4150 3130
rect 5800 3120 6350 3130
rect 6550 3120 6650 3130
rect 9100 3120 9150 3130
rect 1250 3110 1350 3120
rect 2000 3110 2050 3120
rect 3200 3110 3250 3120
rect 3750 3110 4000 3120
rect 4050 3110 4150 3120
rect 5800 3110 6350 3120
rect 6550 3110 6650 3120
rect 9100 3110 9150 3120
rect 1250 3100 1350 3110
rect 2000 3100 2050 3110
rect 3200 3100 3250 3110
rect 3750 3100 4000 3110
rect 4050 3100 4150 3110
rect 5800 3100 6350 3110
rect 6550 3100 6650 3110
rect 9100 3100 9150 3110
rect 1200 3090 1350 3100
rect 3750 3090 3800 3100
rect 4100 3090 4150 3100
rect 4550 3090 4600 3100
rect 4800 3090 4850 3100
rect 5250 3090 5300 3100
rect 6600 3090 6650 3100
rect 8300 3090 8350 3100
rect 9050 3090 9100 3100
rect 9200 3090 9250 3100
rect 9400 3090 9450 3100
rect 1200 3080 1350 3090
rect 3750 3080 3800 3090
rect 4100 3080 4150 3090
rect 4550 3080 4600 3090
rect 4800 3080 4850 3090
rect 5250 3080 5300 3090
rect 6600 3080 6650 3090
rect 8300 3080 8350 3090
rect 9050 3080 9100 3090
rect 9200 3080 9250 3090
rect 9400 3080 9450 3090
rect 1200 3070 1350 3080
rect 3750 3070 3800 3080
rect 4100 3070 4150 3080
rect 4550 3070 4600 3080
rect 4800 3070 4850 3080
rect 5250 3070 5300 3080
rect 6600 3070 6650 3080
rect 8300 3070 8350 3080
rect 9050 3070 9100 3080
rect 9200 3070 9250 3080
rect 9400 3070 9450 3080
rect 1200 3060 1350 3070
rect 3750 3060 3800 3070
rect 4100 3060 4150 3070
rect 4550 3060 4600 3070
rect 4800 3060 4850 3070
rect 5250 3060 5300 3070
rect 6600 3060 6650 3070
rect 8300 3060 8350 3070
rect 9050 3060 9100 3070
rect 9200 3060 9250 3070
rect 9400 3060 9450 3070
rect 1200 3050 1350 3060
rect 3750 3050 3800 3060
rect 4100 3050 4150 3060
rect 4550 3050 4600 3060
rect 4800 3050 4850 3060
rect 5250 3050 5300 3060
rect 6600 3050 6650 3060
rect 8300 3050 8350 3060
rect 9050 3050 9100 3060
rect 9200 3050 9250 3060
rect 9400 3050 9450 3060
rect 1200 3040 1300 3050
rect 3700 3040 3750 3050
rect 4050 3040 4200 3050
rect 4650 3040 4750 3050
rect 6500 3040 6550 3050
rect 6600 3040 6650 3050
rect 9050 3040 9400 3050
rect 1200 3030 1300 3040
rect 3700 3030 3750 3040
rect 4050 3030 4200 3040
rect 4650 3030 4750 3040
rect 6500 3030 6550 3040
rect 6600 3030 6650 3040
rect 9050 3030 9400 3040
rect 1200 3020 1300 3030
rect 3700 3020 3750 3030
rect 4050 3020 4200 3030
rect 4650 3020 4750 3030
rect 6500 3020 6550 3030
rect 6600 3020 6650 3030
rect 9050 3020 9400 3030
rect 1200 3010 1300 3020
rect 3700 3010 3750 3020
rect 4050 3010 4200 3020
rect 4650 3010 4750 3020
rect 6500 3010 6550 3020
rect 6600 3010 6650 3020
rect 9050 3010 9400 3020
rect 1200 3000 1300 3010
rect 3700 3000 3750 3010
rect 4050 3000 4200 3010
rect 4650 3000 4750 3010
rect 6500 3000 6550 3010
rect 6600 3000 6650 3010
rect 9050 3000 9400 3010
rect 1150 2990 1300 3000
rect 1950 2990 2000 3000
rect 3750 2990 3850 3000
rect 4200 2990 4300 3000
rect 5200 2990 5250 3000
rect 6500 2990 6650 3000
rect 8250 2990 8300 3000
rect 9050 2990 9150 3000
rect 9200 2990 9250 3000
rect 1150 2980 1300 2990
rect 1950 2980 2000 2990
rect 3750 2980 3850 2990
rect 4200 2980 4300 2990
rect 5200 2980 5250 2990
rect 6500 2980 6650 2990
rect 8250 2980 8300 2990
rect 9050 2980 9150 2990
rect 9200 2980 9250 2990
rect 1150 2970 1300 2980
rect 1950 2970 2000 2980
rect 3750 2970 3850 2980
rect 4200 2970 4300 2980
rect 5200 2970 5250 2980
rect 6500 2970 6650 2980
rect 8250 2970 8300 2980
rect 9050 2970 9150 2980
rect 9200 2970 9250 2980
rect 1150 2960 1300 2970
rect 1950 2960 2000 2970
rect 3750 2960 3850 2970
rect 4200 2960 4300 2970
rect 5200 2960 5250 2970
rect 6500 2960 6650 2970
rect 8250 2960 8300 2970
rect 9050 2960 9150 2970
rect 9200 2960 9250 2970
rect 1150 2950 1300 2960
rect 1950 2950 2000 2960
rect 3750 2950 3850 2960
rect 4200 2950 4300 2960
rect 5200 2950 5250 2960
rect 6500 2950 6650 2960
rect 8250 2950 8300 2960
rect 9050 2950 9150 2960
rect 9200 2950 9250 2960
rect 1150 2940 1300 2950
rect 1950 2940 2000 2950
rect 3150 2940 3200 2950
rect 3800 2940 3850 2950
rect 4250 2940 4350 2950
rect 6500 2940 6600 2950
rect 9000 2940 9100 2950
rect 1150 2930 1300 2940
rect 1950 2930 2000 2940
rect 3150 2930 3200 2940
rect 3800 2930 3850 2940
rect 4250 2930 4350 2940
rect 6500 2930 6600 2940
rect 9000 2930 9100 2940
rect 1150 2920 1300 2930
rect 1950 2920 2000 2930
rect 3150 2920 3200 2930
rect 3800 2920 3850 2930
rect 4250 2920 4350 2930
rect 6500 2920 6600 2930
rect 9000 2920 9100 2930
rect 1150 2910 1300 2920
rect 1950 2910 2000 2920
rect 3150 2910 3200 2920
rect 3800 2910 3850 2920
rect 4250 2910 4350 2920
rect 6500 2910 6600 2920
rect 9000 2910 9100 2920
rect 1150 2900 1300 2910
rect 1950 2900 2000 2910
rect 3150 2900 3200 2910
rect 3800 2900 3850 2910
rect 4250 2900 4350 2910
rect 6500 2900 6600 2910
rect 9000 2900 9100 2910
rect 1150 2890 1250 2900
rect 1950 2890 2000 2900
rect 3150 2890 3200 2900
rect 3850 2890 3950 2900
rect 4250 2890 4300 2900
rect 4350 2890 4450 2900
rect 5150 2890 5200 2900
rect 6500 2890 6600 2900
rect 7200 2890 7250 2900
rect 1150 2880 1250 2890
rect 1950 2880 2000 2890
rect 3150 2880 3200 2890
rect 3850 2880 3950 2890
rect 4250 2880 4300 2890
rect 4350 2880 4450 2890
rect 5150 2880 5200 2890
rect 6500 2880 6600 2890
rect 7200 2880 7250 2890
rect 1150 2870 1250 2880
rect 1950 2870 2000 2880
rect 3150 2870 3200 2880
rect 3850 2870 3950 2880
rect 4250 2870 4300 2880
rect 4350 2870 4450 2880
rect 5150 2870 5200 2880
rect 6500 2870 6600 2880
rect 7200 2870 7250 2880
rect 1150 2860 1250 2870
rect 1950 2860 2000 2870
rect 3150 2860 3200 2870
rect 3850 2860 3950 2870
rect 4250 2860 4300 2870
rect 4350 2860 4450 2870
rect 5150 2860 5200 2870
rect 6500 2860 6600 2870
rect 7200 2860 7250 2870
rect 1150 2850 1250 2860
rect 1950 2850 2000 2860
rect 3150 2850 3200 2860
rect 3850 2850 3950 2860
rect 4250 2850 4300 2860
rect 4350 2850 4450 2860
rect 5150 2850 5200 2860
rect 6500 2850 6600 2860
rect 7200 2850 7250 2860
rect 1100 2840 1250 2850
rect 1950 2840 2000 2850
rect 3150 2840 3200 2850
rect 3900 2840 3950 2850
rect 4450 2840 4500 2850
rect 5100 2840 5200 2850
rect 5850 2840 6100 2850
rect 6500 2840 6600 2850
rect 7100 2840 7150 2850
rect 8150 2840 8200 2850
rect 1100 2830 1250 2840
rect 1950 2830 2000 2840
rect 3150 2830 3200 2840
rect 3900 2830 3950 2840
rect 4450 2830 4500 2840
rect 5100 2830 5200 2840
rect 5850 2830 6100 2840
rect 6500 2830 6600 2840
rect 7100 2830 7150 2840
rect 8150 2830 8200 2840
rect 1100 2820 1250 2830
rect 1950 2820 2000 2830
rect 3150 2820 3200 2830
rect 3900 2820 3950 2830
rect 4450 2820 4500 2830
rect 5100 2820 5200 2830
rect 5850 2820 6100 2830
rect 6500 2820 6600 2830
rect 7100 2820 7150 2830
rect 8150 2820 8200 2830
rect 1100 2810 1250 2820
rect 1950 2810 2000 2820
rect 3150 2810 3200 2820
rect 3900 2810 3950 2820
rect 4450 2810 4500 2820
rect 5100 2810 5200 2820
rect 5850 2810 6100 2820
rect 6500 2810 6600 2820
rect 7100 2810 7150 2820
rect 8150 2810 8200 2820
rect 1100 2800 1250 2810
rect 1950 2800 2000 2810
rect 3150 2800 3200 2810
rect 3900 2800 3950 2810
rect 4450 2800 4500 2810
rect 5100 2800 5200 2810
rect 5850 2800 6100 2810
rect 6500 2800 6600 2810
rect 7100 2800 7150 2810
rect 8150 2800 8200 2810
rect 1100 2790 1200 2800
rect 1950 2790 2000 2800
rect 3150 2790 3200 2800
rect 4500 2790 4750 2800
rect 5150 2790 5200 2800
rect 5550 2790 6000 2800
rect 6100 2790 6150 2800
rect 6500 2790 6550 2800
rect 7000 2790 7050 2800
rect 7650 2790 7700 2800
rect 8100 2790 8150 2800
rect 1100 2780 1200 2790
rect 1950 2780 2000 2790
rect 3150 2780 3200 2790
rect 4500 2780 4750 2790
rect 5150 2780 5200 2790
rect 5550 2780 6000 2790
rect 6100 2780 6150 2790
rect 6500 2780 6550 2790
rect 7000 2780 7050 2790
rect 7650 2780 7700 2790
rect 8100 2780 8150 2790
rect 1100 2770 1200 2780
rect 1950 2770 2000 2780
rect 3150 2770 3200 2780
rect 4500 2770 4750 2780
rect 5150 2770 5200 2780
rect 5550 2770 6000 2780
rect 6100 2770 6150 2780
rect 6500 2770 6550 2780
rect 7000 2770 7050 2780
rect 7650 2770 7700 2780
rect 8100 2770 8150 2780
rect 1100 2760 1200 2770
rect 1950 2760 2000 2770
rect 3150 2760 3200 2770
rect 4500 2760 4750 2770
rect 5150 2760 5200 2770
rect 5550 2760 6000 2770
rect 6100 2760 6150 2770
rect 6500 2760 6550 2770
rect 7000 2760 7050 2770
rect 7650 2760 7700 2770
rect 8100 2760 8150 2770
rect 1100 2750 1200 2760
rect 1950 2750 2000 2760
rect 3150 2750 3200 2760
rect 4500 2750 4750 2760
rect 5150 2750 5200 2760
rect 5550 2750 6000 2760
rect 6100 2750 6150 2760
rect 6500 2750 6550 2760
rect 7000 2750 7050 2760
rect 7650 2750 7700 2760
rect 8100 2750 8150 2760
rect 1050 2740 1200 2750
rect 1950 2740 2000 2750
rect 3150 2740 3200 2750
rect 3850 2740 3900 2750
rect 4650 2740 5000 2750
rect 5150 2740 5200 2750
rect 5250 2740 5350 2750
rect 5450 2740 5900 2750
rect 6150 2740 6200 2750
rect 6500 2740 6550 2750
rect 8050 2740 8100 2750
rect 8750 2740 8800 2750
rect 1050 2730 1200 2740
rect 1950 2730 2000 2740
rect 3150 2730 3200 2740
rect 3850 2730 3900 2740
rect 4650 2730 5000 2740
rect 5150 2730 5200 2740
rect 5250 2730 5350 2740
rect 5450 2730 5900 2740
rect 6150 2730 6200 2740
rect 6500 2730 6550 2740
rect 8050 2730 8100 2740
rect 8750 2730 8800 2740
rect 1050 2720 1200 2730
rect 1950 2720 2000 2730
rect 3150 2720 3200 2730
rect 3850 2720 3900 2730
rect 4650 2720 5000 2730
rect 5150 2720 5200 2730
rect 5250 2720 5350 2730
rect 5450 2720 5900 2730
rect 6150 2720 6200 2730
rect 6500 2720 6550 2730
rect 8050 2720 8100 2730
rect 8750 2720 8800 2730
rect 1050 2710 1200 2720
rect 1950 2710 2000 2720
rect 3150 2710 3200 2720
rect 3850 2710 3900 2720
rect 4650 2710 5000 2720
rect 5150 2710 5200 2720
rect 5250 2710 5350 2720
rect 5450 2710 5900 2720
rect 6150 2710 6200 2720
rect 6500 2710 6550 2720
rect 8050 2710 8100 2720
rect 8750 2710 8800 2720
rect 1050 2700 1200 2710
rect 1950 2700 2000 2710
rect 3150 2700 3200 2710
rect 3850 2700 3900 2710
rect 4650 2700 5000 2710
rect 5150 2700 5200 2710
rect 5250 2700 5350 2710
rect 5450 2700 5900 2710
rect 6150 2700 6200 2710
rect 6500 2700 6550 2710
rect 8050 2700 8100 2710
rect 8750 2700 8800 2710
rect 1050 2690 1150 2700
rect 3150 2690 3200 2700
rect 3850 2690 3900 2700
rect 4800 2690 4950 2700
rect 5100 2690 5850 2700
rect 6200 2690 6250 2700
rect 6500 2690 6550 2700
rect 6850 2690 6900 2700
rect 7700 2690 7750 2700
rect 8000 2690 8050 2700
rect 1050 2680 1150 2690
rect 3150 2680 3200 2690
rect 3850 2680 3900 2690
rect 4800 2680 4950 2690
rect 5100 2680 5850 2690
rect 6200 2680 6250 2690
rect 6500 2680 6550 2690
rect 6850 2680 6900 2690
rect 7700 2680 7750 2690
rect 8000 2680 8050 2690
rect 1050 2670 1150 2680
rect 3150 2670 3200 2680
rect 3850 2670 3900 2680
rect 4800 2670 4950 2680
rect 5100 2670 5850 2680
rect 6200 2670 6250 2680
rect 6500 2670 6550 2680
rect 6850 2670 6900 2680
rect 7700 2670 7750 2680
rect 8000 2670 8050 2680
rect 1050 2660 1150 2670
rect 3150 2660 3200 2670
rect 3850 2660 3900 2670
rect 4800 2660 4950 2670
rect 5100 2660 5850 2670
rect 6200 2660 6250 2670
rect 6500 2660 6550 2670
rect 6850 2660 6900 2670
rect 7700 2660 7750 2670
rect 8000 2660 8050 2670
rect 1050 2650 1150 2660
rect 3150 2650 3200 2660
rect 3850 2650 3900 2660
rect 4800 2650 4950 2660
rect 5100 2650 5850 2660
rect 6200 2650 6250 2660
rect 6500 2650 6550 2660
rect 6850 2650 6900 2660
rect 7700 2650 7750 2660
rect 8000 2650 8050 2660
rect 1000 2640 1100 2650
rect 1900 2640 1950 2650
rect 2250 2640 2400 2650
rect 2850 2640 2900 2650
rect 3100 2640 3150 2650
rect 3850 2640 3900 2650
rect 4800 2640 4950 2650
rect 5050 2640 5800 2650
rect 6250 2640 6300 2650
rect 7750 2640 7800 2650
rect 7950 2640 8000 2650
rect 9050 2640 9150 2650
rect 1000 2630 1100 2640
rect 1900 2630 1950 2640
rect 2250 2630 2400 2640
rect 2850 2630 2900 2640
rect 3100 2630 3150 2640
rect 3850 2630 3900 2640
rect 4800 2630 4950 2640
rect 5050 2630 5800 2640
rect 6250 2630 6300 2640
rect 7750 2630 7800 2640
rect 7950 2630 8000 2640
rect 9050 2630 9150 2640
rect 1000 2620 1100 2630
rect 1900 2620 1950 2630
rect 2250 2620 2400 2630
rect 2850 2620 2900 2630
rect 3100 2620 3150 2630
rect 3850 2620 3900 2630
rect 4800 2620 4950 2630
rect 5050 2620 5800 2630
rect 6250 2620 6300 2630
rect 7750 2620 7800 2630
rect 7950 2620 8000 2630
rect 9050 2620 9150 2630
rect 1000 2610 1100 2620
rect 1900 2610 1950 2620
rect 2250 2610 2400 2620
rect 2850 2610 2900 2620
rect 3100 2610 3150 2620
rect 3850 2610 3900 2620
rect 4800 2610 4950 2620
rect 5050 2610 5800 2620
rect 6250 2610 6300 2620
rect 7750 2610 7800 2620
rect 7950 2610 8000 2620
rect 9050 2610 9150 2620
rect 1000 2600 1100 2610
rect 1900 2600 1950 2610
rect 2250 2600 2400 2610
rect 2850 2600 2900 2610
rect 3100 2600 3150 2610
rect 3850 2600 3900 2610
rect 4800 2600 4950 2610
rect 5050 2600 5800 2610
rect 6250 2600 6300 2610
rect 7750 2600 7800 2610
rect 7950 2600 8000 2610
rect 9050 2600 9150 2610
rect 1000 2590 1100 2600
rect 2050 2590 2250 2600
rect 2300 2590 2400 2600
rect 2850 2590 3150 2600
rect 3850 2590 3900 2600
rect 4500 2590 5750 2600
rect 6250 2590 6300 2600
rect 7900 2590 7950 2600
rect 9050 2590 9150 2600
rect 1000 2580 1100 2590
rect 2050 2580 2250 2590
rect 2300 2580 2400 2590
rect 2850 2580 3150 2590
rect 3850 2580 3900 2590
rect 4500 2580 5750 2590
rect 6250 2580 6300 2590
rect 7900 2580 7950 2590
rect 9050 2580 9150 2590
rect 1000 2570 1100 2580
rect 2050 2570 2250 2580
rect 2300 2570 2400 2580
rect 2850 2570 3150 2580
rect 3850 2570 3900 2580
rect 4500 2570 5750 2580
rect 6250 2570 6300 2580
rect 7900 2570 7950 2580
rect 9050 2570 9150 2580
rect 1000 2560 1100 2570
rect 2050 2560 2250 2570
rect 2300 2560 2400 2570
rect 2850 2560 3150 2570
rect 3850 2560 3900 2570
rect 4500 2560 5750 2570
rect 6250 2560 6300 2570
rect 7900 2560 7950 2570
rect 9050 2560 9150 2570
rect 1000 2550 1100 2560
rect 2050 2550 2250 2560
rect 2300 2550 2400 2560
rect 2850 2550 3150 2560
rect 3850 2550 3900 2560
rect 4500 2550 5750 2560
rect 6250 2550 6300 2560
rect 7900 2550 7950 2560
rect 9050 2550 9150 2560
rect 950 2540 1050 2550
rect 3200 2540 3250 2550
rect 3900 2540 3950 2550
rect 4200 2540 4250 2550
rect 4650 2540 5750 2550
rect 6300 2540 6350 2550
rect 7800 2540 7850 2550
rect 950 2530 1050 2540
rect 3200 2530 3250 2540
rect 3900 2530 3950 2540
rect 4200 2530 4250 2540
rect 4650 2530 5750 2540
rect 6300 2530 6350 2540
rect 7800 2530 7850 2540
rect 950 2520 1050 2530
rect 3200 2520 3250 2530
rect 3900 2520 3950 2530
rect 4200 2520 4250 2530
rect 4650 2520 5750 2530
rect 6300 2520 6350 2530
rect 7800 2520 7850 2530
rect 950 2510 1050 2520
rect 3200 2510 3250 2520
rect 3900 2510 3950 2520
rect 4200 2510 4250 2520
rect 4650 2510 5750 2520
rect 6300 2510 6350 2520
rect 7800 2510 7850 2520
rect 950 2500 1050 2510
rect 3200 2500 3250 2510
rect 3900 2500 3950 2510
rect 4200 2500 4250 2510
rect 4650 2500 5750 2510
rect 6300 2500 6350 2510
rect 7800 2500 7850 2510
rect 950 2490 1050 2500
rect 1850 2490 1900 2500
rect 3250 2490 3300 2500
rect 3950 2490 4000 2500
rect 4050 2490 4150 2500
rect 4600 2490 5550 2500
rect 6700 2490 6750 2500
rect 9400 2490 9450 2500
rect 950 2480 1050 2490
rect 1850 2480 1900 2490
rect 3250 2480 3300 2490
rect 3950 2480 4000 2490
rect 4050 2480 4150 2490
rect 4600 2480 5550 2490
rect 6700 2480 6750 2490
rect 9400 2480 9450 2490
rect 950 2470 1050 2480
rect 1850 2470 1900 2480
rect 3250 2470 3300 2480
rect 3950 2470 4000 2480
rect 4050 2470 4150 2480
rect 4600 2470 5550 2480
rect 6700 2470 6750 2480
rect 9400 2470 9450 2480
rect 950 2460 1050 2470
rect 1850 2460 1900 2470
rect 3250 2460 3300 2470
rect 3950 2460 4000 2470
rect 4050 2460 4150 2470
rect 4600 2460 5550 2470
rect 6700 2460 6750 2470
rect 9400 2460 9450 2470
rect 950 2450 1050 2460
rect 1850 2450 1900 2460
rect 3250 2450 3300 2460
rect 3950 2450 4000 2460
rect 4050 2450 4150 2460
rect 4600 2450 5550 2460
rect 6700 2450 6750 2460
rect 9400 2450 9450 2460
rect 900 2440 1050 2450
rect 1850 2440 1900 2450
rect 3250 2440 3300 2450
rect 4000 2440 4050 2450
rect 4550 2440 5550 2450
rect 6350 2440 6400 2450
rect 6700 2440 6750 2450
rect 900 2430 1050 2440
rect 1850 2430 1900 2440
rect 3250 2430 3300 2440
rect 4000 2430 4050 2440
rect 4550 2430 5550 2440
rect 6350 2430 6400 2440
rect 6700 2430 6750 2440
rect 900 2420 1050 2430
rect 1850 2420 1900 2430
rect 3250 2420 3300 2430
rect 4000 2420 4050 2430
rect 4550 2420 5550 2430
rect 6350 2420 6400 2430
rect 6700 2420 6750 2430
rect 900 2410 1050 2420
rect 1850 2410 1900 2420
rect 3250 2410 3300 2420
rect 4000 2410 4050 2420
rect 4550 2410 5550 2420
rect 6350 2410 6400 2420
rect 6700 2410 6750 2420
rect 900 2400 1050 2410
rect 1850 2400 1900 2410
rect 3250 2400 3300 2410
rect 4000 2400 4050 2410
rect 4550 2400 5550 2410
rect 6350 2400 6400 2410
rect 6700 2400 6750 2410
rect 900 2390 1050 2400
rect 1850 2390 1900 2400
rect 4500 2390 5650 2400
rect 6700 2390 6750 2400
rect 900 2380 1050 2390
rect 1850 2380 1900 2390
rect 4500 2380 5650 2390
rect 6700 2380 6750 2390
rect 900 2370 1050 2380
rect 1850 2370 1900 2380
rect 4500 2370 5650 2380
rect 6700 2370 6750 2380
rect 900 2360 1050 2370
rect 1850 2360 1900 2370
rect 4500 2360 5650 2370
rect 6700 2360 6750 2370
rect 900 2350 1050 2360
rect 1850 2350 1900 2360
rect 4500 2350 5650 2360
rect 6700 2350 6750 2360
rect 850 2340 1000 2350
rect 3300 2340 3350 2350
rect 4450 2340 5650 2350
rect 6400 2340 6450 2350
rect 6700 2340 6750 2350
rect 9650 2340 9750 2350
rect 850 2330 1000 2340
rect 3300 2330 3350 2340
rect 4450 2330 5650 2340
rect 6400 2330 6450 2340
rect 6700 2330 6750 2340
rect 9650 2330 9750 2340
rect 850 2320 1000 2330
rect 3300 2320 3350 2330
rect 4450 2320 5650 2330
rect 6400 2320 6450 2330
rect 6700 2320 6750 2330
rect 9650 2320 9750 2330
rect 850 2310 1000 2320
rect 3300 2310 3350 2320
rect 4450 2310 5650 2320
rect 6400 2310 6450 2320
rect 6700 2310 6750 2320
rect 9650 2310 9750 2320
rect 850 2300 1000 2310
rect 3300 2300 3350 2310
rect 4450 2300 5650 2310
rect 6400 2300 6450 2310
rect 6700 2300 6750 2310
rect 9650 2300 9750 2310
rect 850 2290 1000 2300
rect 1800 2290 1850 2300
rect 3300 2290 3350 2300
rect 4100 2290 5400 2300
rect 5550 2290 5600 2300
rect 6450 2290 6500 2300
rect 6700 2290 6750 2300
rect 6850 2290 6950 2300
rect 8500 2290 8550 2300
rect 9150 2290 9250 2300
rect 9350 2290 9450 2300
rect 9600 2290 9750 2300
rect 850 2280 1000 2290
rect 1800 2280 1850 2290
rect 3300 2280 3350 2290
rect 4100 2280 5400 2290
rect 5550 2280 5600 2290
rect 6450 2280 6500 2290
rect 6700 2280 6750 2290
rect 6850 2280 6950 2290
rect 8500 2280 8550 2290
rect 9150 2280 9250 2290
rect 9350 2280 9450 2290
rect 9600 2280 9750 2290
rect 850 2270 1000 2280
rect 1800 2270 1850 2280
rect 3300 2270 3350 2280
rect 4100 2270 5400 2280
rect 5550 2270 5600 2280
rect 6450 2270 6500 2280
rect 6700 2270 6750 2280
rect 6850 2270 6950 2280
rect 8500 2270 8550 2280
rect 9150 2270 9250 2280
rect 9350 2270 9450 2280
rect 9600 2270 9750 2280
rect 850 2260 1000 2270
rect 1800 2260 1850 2270
rect 3300 2260 3350 2270
rect 4100 2260 5400 2270
rect 5550 2260 5600 2270
rect 6450 2260 6500 2270
rect 6700 2260 6750 2270
rect 6850 2260 6950 2270
rect 8500 2260 8550 2270
rect 9150 2260 9250 2270
rect 9350 2260 9450 2270
rect 9600 2260 9750 2270
rect 850 2250 1000 2260
rect 1800 2250 1850 2260
rect 3300 2250 3350 2260
rect 4100 2250 5400 2260
rect 5550 2250 5600 2260
rect 6450 2250 6500 2260
rect 6700 2250 6750 2260
rect 6850 2250 6950 2260
rect 8500 2250 8550 2260
rect 9150 2250 9250 2260
rect 9350 2250 9450 2260
rect 9600 2250 9750 2260
rect 800 2240 1000 2250
rect 1800 2240 1850 2250
rect 3300 2240 3350 2250
rect 4350 2240 5350 2250
rect 6700 2240 6750 2250
rect 6900 2240 7250 2250
rect 7550 2240 7600 2250
rect 8600 2240 8650 2250
rect 9100 2240 9150 2250
rect 9450 2240 9500 2250
rect 9550 2240 9750 2250
rect 800 2230 1000 2240
rect 1800 2230 1850 2240
rect 3300 2230 3350 2240
rect 4350 2230 5350 2240
rect 6700 2230 6750 2240
rect 6900 2230 7250 2240
rect 7550 2230 7600 2240
rect 8600 2230 8650 2240
rect 9100 2230 9150 2240
rect 9450 2230 9500 2240
rect 9550 2230 9750 2240
rect 800 2220 1000 2230
rect 1800 2220 1850 2230
rect 3300 2220 3350 2230
rect 4350 2220 5350 2230
rect 6700 2220 6750 2230
rect 6900 2220 7250 2230
rect 7550 2220 7600 2230
rect 8600 2220 8650 2230
rect 9100 2220 9150 2230
rect 9450 2220 9500 2230
rect 9550 2220 9750 2230
rect 800 2210 1000 2220
rect 1800 2210 1850 2220
rect 3300 2210 3350 2220
rect 4350 2210 5350 2220
rect 6700 2210 6750 2220
rect 6900 2210 7250 2220
rect 7550 2210 7600 2220
rect 8600 2210 8650 2220
rect 9100 2210 9150 2220
rect 9450 2210 9500 2220
rect 9550 2210 9750 2220
rect 800 2200 1000 2210
rect 1800 2200 1850 2210
rect 3300 2200 3350 2210
rect 4350 2200 5350 2210
rect 6700 2200 6750 2210
rect 6900 2200 7250 2210
rect 7550 2200 7600 2210
rect 8600 2200 8650 2210
rect 9100 2200 9150 2210
rect 9450 2200 9500 2210
rect 9550 2200 9750 2210
rect 800 2190 1000 2200
rect 1800 2190 1850 2200
rect 3300 2190 3350 2200
rect 4350 2190 5300 2200
rect 6500 2190 6550 2200
rect 6700 2190 6750 2200
rect 7000 2190 7100 2200
rect 7250 2190 7350 2200
rect 7500 2190 7550 2200
rect 7600 2190 7650 2200
rect 8800 2190 9050 2200
rect 9600 2190 9650 2200
rect 800 2180 1000 2190
rect 1800 2180 1850 2190
rect 3300 2180 3350 2190
rect 4350 2180 5300 2190
rect 6500 2180 6550 2190
rect 6700 2180 6750 2190
rect 7000 2180 7100 2190
rect 7250 2180 7350 2190
rect 7500 2180 7550 2190
rect 7600 2180 7650 2190
rect 8800 2180 9050 2190
rect 9600 2180 9650 2190
rect 800 2170 1000 2180
rect 1800 2170 1850 2180
rect 3300 2170 3350 2180
rect 4350 2170 5300 2180
rect 6500 2170 6550 2180
rect 6700 2170 6750 2180
rect 7000 2170 7100 2180
rect 7250 2170 7350 2180
rect 7500 2170 7550 2180
rect 7600 2170 7650 2180
rect 8800 2170 9050 2180
rect 9600 2170 9650 2180
rect 800 2160 1000 2170
rect 1800 2160 1850 2170
rect 3300 2160 3350 2170
rect 4350 2160 5300 2170
rect 6500 2160 6550 2170
rect 6700 2160 6750 2170
rect 7000 2160 7100 2170
rect 7250 2160 7350 2170
rect 7500 2160 7550 2170
rect 7600 2160 7650 2170
rect 8800 2160 9050 2170
rect 9600 2160 9650 2170
rect 800 2150 1000 2160
rect 1800 2150 1850 2160
rect 3300 2150 3350 2160
rect 4350 2150 5300 2160
rect 6500 2150 6550 2160
rect 6700 2150 6750 2160
rect 7000 2150 7100 2160
rect 7250 2150 7350 2160
rect 7500 2150 7550 2160
rect 7600 2150 7650 2160
rect 8800 2150 9050 2160
rect 9600 2150 9650 2160
rect 750 2140 1000 2150
rect 1800 2140 1850 2150
rect 3300 2140 3350 2150
rect 4350 2140 5250 2150
rect 6500 2140 6550 2150
rect 6700 2140 6750 2150
rect 7050 2140 7250 2150
rect 7350 2140 7500 2150
rect 7700 2140 7750 2150
rect 8400 2140 8450 2150
rect 750 2130 1000 2140
rect 1800 2130 1850 2140
rect 3300 2130 3350 2140
rect 4350 2130 5250 2140
rect 6500 2130 6550 2140
rect 6700 2130 6750 2140
rect 7050 2130 7250 2140
rect 7350 2130 7500 2140
rect 7700 2130 7750 2140
rect 8400 2130 8450 2140
rect 750 2120 1000 2130
rect 1800 2120 1850 2130
rect 3300 2120 3350 2130
rect 4350 2120 5250 2130
rect 6500 2120 6550 2130
rect 6700 2120 6750 2130
rect 7050 2120 7250 2130
rect 7350 2120 7500 2130
rect 7700 2120 7750 2130
rect 8400 2120 8450 2130
rect 750 2110 1000 2120
rect 1800 2110 1850 2120
rect 3300 2110 3350 2120
rect 4350 2110 5250 2120
rect 6500 2110 6550 2120
rect 6700 2110 6750 2120
rect 7050 2110 7250 2120
rect 7350 2110 7500 2120
rect 7700 2110 7750 2120
rect 8400 2110 8450 2120
rect 750 2100 1000 2110
rect 1800 2100 1850 2110
rect 3300 2100 3350 2110
rect 4350 2100 5250 2110
rect 6500 2100 6550 2110
rect 6700 2100 6750 2110
rect 7050 2100 7250 2110
rect 7350 2100 7500 2110
rect 7700 2100 7750 2110
rect 8400 2100 8450 2110
rect 750 2090 950 2100
rect 1800 2090 1850 2100
rect 3300 2090 3350 2100
rect 4350 2090 5100 2100
rect 5150 2090 5250 2100
rect 7800 2090 7850 2100
rect 8450 2090 8550 2100
rect 9100 2090 9150 2100
rect 750 2080 950 2090
rect 1800 2080 1850 2090
rect 3300 2080 3350 2090
rect 4350 2080 5100 2090
rect 5150 2080 5250 2090
rect 7800 2080 7850 2090
rect 8450 2080 8550 2090
rect 9100 2080 9150 2090
rect 750 2070 950 2080
rect 1800 2070 1850 2080
rect 3300 2070 3350 2080
rect 4350 2070 5100 2080
rect 5150 2070 5250 2080
rect 7800 2070 7850 2080
rect 8450 2070 8550 2080
rect 9100 2070 9150 2080
rect 750 2060 950 2070
rect 1800 2060 1850 2070
rect 3300 2060 3350 2070
rect 4350 2060 5100 2070
rect 5150 2060 5250 2070
rect 7800 2060 7850 2070
rect 8450 2060 8550 2070
rect 9100 2060 9150 2070
rect 750 2050 950 2060
rect 1800 2050 1850 2060
rect 3300 2050 3350 2060
rect 4350 2050 5100 2060
rect 5150 2050 5250 2060
rect 7800 2050 7850 2060
rect 8450 2050 8550 2060
rect 9100 2050 9150 2060
rect 700 2040 950 2050
rect 1800 2040 1850 2050
rect 3300 2040 3350 2050
rect 4350 2040 5100 2050
rect 7750 2040 7900 2050
rect 8550 2040 8650 2050
rect 700 2030 950 2040
rect 1800 2030 1850 2040
rect 3300 2030 3350 2040
rect 4350 2030 5100 2040
rect 7750 2030 7900 2040
rect 8550 2030 8650 2040
rect 700 2020 950 2030
rect 1800 2020 1850 2030
rect 3300 2020 3350 2030
rect 4350 2020 5100 2030
rect 7750 2020 7900 2030
rect 8550 2020 8650 2030
rect 700 2010 950 2020
rect 1800 2010 1850 2020
rect 3300 2010 3350 2020
rect 4350 2010 5100 2020
rect 7750 2010 7900 2020
rect 8550 2010 8650 2020
rect 700 2000 950 2010
rect 1800 2000 1850 2010
rect 3300 2000 3350 2010
rect 4350 2000 5100 2010
rect 7750 2000 7900 2010
rect 8550 2000 8650 2010
rect 700 1990 950 2000
rect 1800 1990 1850 2000
rect 4350 1990 4800 2000
rect 4850 1990 5000 2000
rect 6750 1990 6800 2000
rect 7350 1990 7400 2000
rect 7700 1990 7750 2000
rect 700 1980 950 1990
rect 1800 1980 1850 1990
rect 4350 1980 4800 1990
rect 4850 1980 5000 1990
rect 6750 1980 6800 1990
rect 7350 1980 7400 1990
rect 7700 1980 7750 1990
rect 700 1970 950 1980
rect 1800 1970 1850 1980
rect 4350 1970 4800 1980
rect 4850 1970 5000 1980
rect 6750 1970 6800 1980
rect 7350 1970 7400 1980
rect 7700 1970 7750 1980
rect 700 1960 950 1970
rect 1800 1960 1850 1970
rect 4350 1960 4800 1970
rect 4850 1960 5000 1970
rect 6750 1960 6800 1970
rect 7350 1960 7400 1970
rect 7700 1960 7750 1970
rect 700 1950 950 1960
rect 1800 1950 1850 1960
rect 4350 1950 4800 1960
rect 4850 1950 5000 1960
rect 6750 1950 6800 1960
rect 7350 1950 7400 1960
rect 7700 1950 7750 1960
rect 650 1940 950 1950
rect 1800 1940 1850 1950
rect 4350 1940 4450 1950
rect 4700 1940 4750 1950
rect 4900 1940 4950 1950
rect 6200 1940 6300 1950
rect 6550 1940 6600 1950
rect 6750 1940 6800 1950
rect 7350 1940 7400 1950
rect 7700 1940 7750 1950
rect 650 1930 950 1940
rect 1800 1930 1850 1940
rect 4350 1930 4450 1940
rect 4700 1930 4750 1940
rect 4900 1930 4950 1940
rect 6200 1930 6300 1940
rect 6550 1930 6600 1940
rect 6750 1930 6800 1940
rect 7350 1930 7400 1940
rect 7700 1930 7750 1940
rect 650 1920 950 1930
rect 1800 1920 1850 1930
rect 4350 1920 4450 1930
rect 4700 1920 4750 1930
rect 4900 1920 4950 1930
rect 6200 1920 6300 1930
rect 6550 1920 6600 1930
rect 6750 1920 6800 1930
rect 7350 1920 7400 1930
rect 7700 1920 7750 1930
rect 650 1910 950 1920
rect 1800 1910 1850 1920
rect 4350 1910 4450 1920
rect 4700 1910 4750 1920
rect 4900 1910 4950 1920
rect 6200 1910 6300 1920
rect 6550 1910 6600 1920
rect 6750 1910 6800 1920
rect 7350 1910 7400 1920
rect 7700 1910 7750 1920
rect 650 1900 950 1910
rect 1800 1900 1850 1910
rect 4350 1900 4450 1910
rect 4700 1900 4750 1910
rect 4900 1900 4950 1910
rect 6200 1900 6300 1910
rect 6550 1900 6600 1910
rect 6750 1900 6800 1910
rect 7350 1900 7400 1910
rect 7700 1900 7750 1910
rect 650 1890 950 1900
rect 1800 1890 1850 1900
rect 4250 1890 4350 1900
rect 6200 1890 6300 1900
rect 6550 1890 6600 1900
rect 6750 1890 6800 1900
rect 7350 1890 7400 1900
rect 7700 1890 7750 1900
rect 650 1880 950 1890
rect 1800 1880 1850 1890
rect 4250 1880 4350 1890
rect 6200 1880 6300 1890
rect 6550 1880 6600 1890
rect 6750 1880 6800 1890
rect 7350 1880 7400 1890
rect 7700 1880 7750 1890
rect 650 1870 950 1880
rect 1800 1870 1850 1880
rect 4250 1870 4350 1880
rect 6200 1870 6300 1880
rect 6550 1870 6600 1880
rect 6750 1870 6800 1880
rect 7350 1870 7400 1880
rect 7700 1870 7750 1880
rect 650 1860 950 1870
rect 1800 1860 1850 1870
rect 4250 1860 4350 1870
rect 6200 1860 6300 1870
rect 6550 1860 6600 1870
rect 6750 1860 6800 1870
rect 7350 1860 7400 1870
rect 7700 1860 7750 1870
rect 650 1850 950 1860
rect 1800 1850 1850 1860
rect 4250 1850 4350 1860
rect 6200 1850 6300 1860
rect 6550 1850 6600 1860
rect 6750 1850 6800 1860
rect 7350 1850 7400 1860
rect 7700 1850 7750 1860
rect 600 1840 900 1850
rect 1800 1840 1850 1850
rect 2450 1840 2750 1850
rect 3300 1840 3350 1850
rect 4050 1840 4100 1850
rect 4200 1840 4450 1850
rect 6150 1840 6250 1850
rect 6500 1840 6600 1850
rect 6750 1840 6800 1850
rect 7350 1840 7400 1850
rect 600 1830 900 1840
rect 1800 1830 1850 1840
rect 2450 1830 2750 1840
rect 3300 1830 3350 1840
rect 4050 1830 4100 1840
rect 4200 1830 4450 1840
rect 6150 1830 6250 1840
rect 6500 1830 6600 1840
rect 6750 1830 6800 1840
rect 7350 1830 7400 1840
rect 600 1820 900 1830
rect 1800 1820 1850 1830
rect 2450 1820 2750 1830
rect 3300 1820 3350 1830
rect 4050 1820 4100 1830
rect 4200 1820 4450 1830
rect 6150 1820 6250 1830
rect 6500 1820 6600 1830
rect 6750 1820 6800 1830
rect 7350 1820 7400 1830
rect 600 1810 900 1820
rect 1800 1810 1850 1820
rect 2450 1810 2750 1820
rect 3300 1810 3350 1820
rect 4050 1810 4100 1820
rect 4200 1810 4450 1820
rect 6150 1810 6250 1820
rect 6500 1810 6600 1820
rect 6750 1810 6800 1820
rect 7350 1810 7400 1820
rect 600 1800 900 1810
rect 1800 1800 1850 1810
rect 2450 1800 2750 1810
rect 3300 1800 3350 1810
rect 4050 1800 4100 1810
rect 4200 1800 4450 1810
rect 6150 1800 6250 1810
rect 6500 1800 6600 1810
rect 6750 1800 6800 1810
rect 7350 1800 7400 1810
rect 600 1790 900 1800
rect 1800 1790 1850 1800
rect 3300 1790 3350 1800
rect 4250 1790 4350 1800
rect 4400 1790 4450 1800
rect 6100 1790 6250 1800
rect 6550 1790 6650 1800
rect 6750 1790 6800 1800
rect 7350 1790 7400 1800
rect 7750 1790 7800 1800
rect 600 1780 900 1790
rect 1800 1780 1850 1790
rect 3300 1780 3350 1790
rect 4250 1780 4350 1790
rect 4400 1780 4450 1790
rect 6100 1780 6250 1790
rect 6550 1780 6650 1790
rect 6750 1780 6800 1790
rect 7350 1780 7400 1790
rect 7750 1780 7800 1790
rect 600 1770 900 1780
rect 1800 1770 1850 1780
rect 3300 1770 3350 1780
rect 4250 1770 4350 1780
rect 4400 1770 4450 1780
rect 6100 1770 6250 1780
rect 6550 1770 6650 1780
rect 6750 1770 6800 1780
rect 7350 1770 7400 1780
rect 7750 1770 7800 1780
rect 600 1760 900 1770
rect 1800 1760 1850 1770
rect 3300 1760 3350 1770
rect 4250 1760 4350 1770
rect 4400 1760 4450 1770
rect 6100 1760 6250 1770
rect 6550 1760 6650 1770
rect 6750 1760 6800 1770
rect 7350 1760 7400 1770
rect 7750 1760 7800 1770
rect 600 1750 900 1760
rect 1800 1750 1850 1760
rect 3300 1750 3350 1760
rect 4250 1750 4350 1760
rect 4400 1750 4450 1760
rect 6100 1750 6250 1760
rect 6550 1750 6650 1760
rect 6750 1750 6800 1760
rect 7350 1750 7400 1760
rect 7750 1750 7800 1760
rect 550 1740 900 1750
rect 3300 1740 3350 1750
rect 4000 1740 4050 1750
rect 4300 1740 4350 1750
rect 4400 1740 4450 1750
rect 6050 1740 6300 1750
rect 6550 1740 6650 1750
rect 6750 1740 6800 1750
rect 7350 1740 7400 1750
rect 7750 1740 7800 1750
rect 550 1730 900 1740
rect 3300 1730 3350 1740
rect 4000 1730 4050 1740
rect 4300 1730 4350 1740
rect 4400 1730 4450 1740
rect 6050 1730 6300 1740
rect 6550 1730 6650 1740
rect 6750 1730 6800 1740
rect 7350 1730 7400 1740
rect 7750 1730 7800 1740
rect 550 1720 900 1730
rect 3300 1720 3350 1730
rect 4000 1720 4050 1730
rect 4300 1720 4350 1730
rect 4400 1720 4450 1730
rect 6050 1720 6300 1730
rect 6550 1720 6650 1730
rect 6750 1720 6800 1730
rect 7350 1720 7400 1730
rect 7750 1720 7800 1730
rect 550 1710 900 1720
rect 3300 1710 3350 1720
rect 4000 1710 4050 1720
rect 4300 1710 4350 1720
rect 4400 1710 4450 1720
rect 6050 1710 6300 1720
rect 6550 1710 6650 1720
rect 6750 1710 6800 1720
rect 7350 1710 7400 1720
rect 7750 1710 7800 1720
rect 550 1700 900 1710
rect 3300 1700 3350 1710
rect 4000 1700 4050 1710
rect 4300 1700 4350 1710
rect 4400 1700 4450 1710
rect 6050 1700 6300 1710
rect 6550 1700 6650 1710
rect 6750 1700 6800 1710
rect 7350 1700 7400 1710
rect 7750 1700 7800 1710
rect 550 1690 900 1700
rect 1850 1690 1900 1700
rect 3250 1690 3300 1700
rect 4300 1690 4350 1700
rect 6050 1690 6300 1700
rect 6550 1690 6650 1700
rect 6750 1690 6800 1700
rect 7750 1690 7800 1700
rect 550 1680 900 1690
rect 1850 1680 1900 1690
rect 3250 1680 3300 1690
rect 4300 1680 4350 1690
rect 6050 1680 6300 1690
rect 6550 1680 6650 1690
rect 6750 1680 6800 1690
rect 7750 1680 7800 1690
rect 550 1670 900 1680
rect 1850 1670 1900 1680
rect 3250 1670 3300 1680
rect 4300 1670 4350 1680
rect 6050 1670 6300 1680
rect 6550 1670 6650 1680
rect 6750 1670 6800 1680
rect 7750 1670 7800 1680
rect 550 1660 900 1670
rect 1850 1660 1900 1670
rect 3250 1660 3300 1670
rect 4300 1660 4350 1670
rect 6050 1660 6300 1670
rect 6550 1660 6650 1670
rect 6750 1660 6800 1670
rect 7750 1660 7800 1670
rect 550 1650 900 1660
rect 1850 1650 1900 1660
rect 3250 1650 3300 1660
rect 4300 1650 4350 1660
rect 6050 1650 6300 1660
rect 6550 1650 6650 1660
rect 6750 1650 6800 1660
rect 7750 1650 7800 1660
rect 550 1640 900 1650
rect 3250 1640 3300 1650
rect 4050 1640 4100 1650
rect 4550 1640 4600 1650
rect 6000 1640 6200 1650
rect 6250 1640 6300 1650
rect 6500 1640 6700 1650
rect 6750 1640 6800 1650
rect 7750 1640 7800 1650
rect 550 1630 900 1640
rect 3250 1630 3300 1640
rect 4050 1630 4100 1640
rect 4550 1630 4600 1640
rect 6000 1630 6200 1640
rect 6250 1630 6300 1640
rect 6500 1630 6700 1640
rect 6750 1630 6800 1640
rect 7750 1630 7800 1640
rect 550 1620 900 1630
rect 3250 1620 3300 1630
rect 4050 1620 4100 1630
rect 4550 1620 4600 1630
rect 6000 1620 6200 1630
rect 6250 1620 6300 1630
rect 6500 1620 6700 1630
rect 6750 1620 6800 1630
rect 7750 1620 7800 1630
rect 550 1610 900 1620
rect 3250 1610 3300 1620
rect 4050 1610 4100 1620
rect 4550 1610 4600 1620
rect 6000 1610 6200 1620
rect 6250 1610 6300 1620
rect 6500 1610 6700 1620
rect 6750 1610 6800 1620
rect 7750 1610 7800 1620
rect 550 1600 900 1610
rect 3250 1600 3300 1610
rect 4050 1600 4100 1610
rect 4550 1600 4600 1610
rect 6000 1600 6200 1610
rect 6250 1600 6300 1610
rect 6500 1600 6700 1610
rect 6750 1600 6800 1610
rect 7750 1600 7800 1610
rect 500 1590 850 1600
rect 1900 1590 1950 1600
rect 3200 1590 3250 1600
rect 4050 1590 4100 1600
rect 4350 1590 4800 1600
rect 6000 1590 6300 1600
rect 6450 1590 6800 1600
rect 7750 1590 7800 1600
rect 500 1580 850 1590
rect 1900 1580 1950 1590
rect 3200 1580 3250 1590
rect 4050 1580 4100 1590
rect 4350 1580 4800 1590
rect 6000 1580 6300 1590
rect 6450 1580 6800 1590
rect 7750 1580 7800 1590
rect 500 1570 850 1580
rect 1900 1570 1950 1580
rect 3200 1570 3250 1580
rect 4050 1570 4100 1580
rect 4350 1570 4800 1580
rect 6000 1570 6300 1580
rect 6450 1570 6800 1580
rect 7750 1570 7800 1580
rect 500 1560 850 1570
rect 1900 1560 1950 1570
rect 3200 1560 3250 1570
rect 4050 1560 4100 1570
rect 4350 1560 4800 1570
rect 6000 1560 6300 1570
rect 6450 1560 6800 1570
rect 7750 1560 7800 1570
rect 500 1550 850 1560
rect 1900 1550 1950 1560
rect 3200 1550 3250 1560
rect 4050 1550 4100 1560
rect 4350 1550 4800 1560
rect 6000 1550 6300 1560
rect 6450 1550 6800 1560
rect 7750 1550 7800 1560
rect 500 1540 850 1550
rect 3150 1540 3200 1550
rect 4350 1540 4850 1550
rect 6000 1540 6250 1550
rect 6400 1540 6800 1550
rect 7750 1540 7800 1550
rect 500 1530 850 1540
rect 3150 1530 3200 1540
rect 4350 1530 4850 1540
rect 6000 1530 6250 1540
rect 6400 1530 6800 1540
rect 7750 1530 7800 1540
rect 500 1520 850 1530
rect 3150 1520 3200 1530
rect 4350 1520 4850 1530
rect 6000 1520 6250 1530
rect 6400 1520 6800 1530
rect 7750 1520 7800 1530
rect 500 1510 850 1520
rect 3150 1510 3200 1520
rect 4350 1510 4850 1520
rect 6000 1510 6250 1520
rect 6400 1510 6800 1520
rect 7750 1510 7800 1520
rect 500 1500 850 1510
rect 3150 1500 3200 1510
rect 4350 1500 4850 1510
rect 6000 1500 6250 1510
rect 6400 1500 6800 1510
rect 7750 1500 7800 1510
rect 500 1490 900 1500
rect 950 1490 1000 1500
rect 1950 1490 2000 1500
rect 3100 1490 3150 1500
rect 4400 1490 4950 1500
rect 5950 1490 6200 1500
rect 6300 1490 6350 1500
rect 6400 1490 6800 1500
rect 500 1480 900 1490
rect 950 1480 1000 1490
rect 1950 1480 2000 1490
rect 3100 1480 3150 1490
rect 4400 1480 4950 1490
rect 5950 1480 6200 1490
rect 6300 1480 6350 1490
rect 6400 1480 6800 1490
rect 500 1470 900 1480
rect 950 1470 1000 1480
rect 1950 1470 2000 1480
rect 3100 1470 3150 1480
rect 4400 1470 4950 1480
rect 5950 1470 6200 1480
rect 6300 1470 6350 1480
rect 6400 1470 6800 1480
rect 500 1460 900 1470
rect 950 1460 1000 1470
rect 1950 1460 2000 1470
rect 3100 1460 3150 1470
rect 4400 1460 4950 1470
rect 5950 1460 6200 1470
rect 6300 1460 6350 1470
rect 6400 1460 6800 1470
rect 500 1450 900 1460
rect 950 1450 1000 1460
rect 1950 1450 2000 1460
rect 3100 1450 3150 1460
rect 4400 1450 4950 1460
rect 5950 1450 6200 1460
rect 6300 1450 6350 1460
rect 6400 1450 6800 1460
rect 450 1440 850 1450
rect 1000 1440 1050 1450
rect 2000 1440 2050 1450
rect 3050 1440 3100 1450
rect 4100 1440 4150 1450
rect 4400 1440 4950 1450
rect 5950 1440 6200 1450
rect 6300 1440 6800 1450
rect 7400 1440 7450 1450
rect 7800 1440 7850 1450
rect 450 1430 850 1440
rect 1000 1430 1050 1440
rect 2000 1430 2050 1440
rect 3050 1430 3100 1440
rect 4100 1430 4150 1440
rect 4400 1430 4950 1440
rect 5950 1430 6200 1440
rect 6300 1430 6800 1440
rect 7400 1430 7450 1440
rect 7800 1430 7850 1440
rect 450 1420 850 1430
rect 1000 1420 1050 1430
rect 2000 1420 2050 1430
rect 3050 1420 3100 1430
rect 4100 1420 4150 1430
rect 4400 1420 4950 1430
rect 5950 1420 6200 1430
rect 6300 1420 6800 1430
rect 7400 1420 7450 1430
rect 7800 1420 7850 1430
rect 450 1410 850 1420
rect 1000 1410 1050 1420
rect 2000 1410 2050 1420
rect 3050 1410 3100 1420
rect 4100 1410 4150 1420
rect 4400 1410 4950 1420
rect 5950 1410 6200 1420
rect 6300 1410 6800 1420
rect 7400 1410 7450 1420
rect 7800 1410 7850 1420
rect 450 1400 850 1410
rect 1000 1400 1050 1410
rect 2000 1400 2050 1410
rect 3050 1400 3100 1410
rect 4100 1400 4150 1410
rect 4400 1400 4950 1410
rect 5950 1400 6200 1410
rect 6300 1400 6800 1410
rect 7400 1400 7450 1410
rect 7800 1400 7850 1410
rect 450 1390 800 1400
rect 1000 1390 1050 1400
rect 2050 1390 2100 1400
rect 3000 1390 3050 1400
rect 3500 1390 3550 1400
rect 3650 1390 3700 1400
rect 4450 1390 5100 1400
rect 5950 1390 6200 1400
rect 6300 1390 6800 1400
rect 7400 1390 7450 1400
rect 7800 1390 7850 1400
rect 450 1380 800 1390
rect 1000 1380 1050 1390
rect 2050 1380 2100 1390
rect 3000 1380 3050 1390
rect 3500 1380 3550 1390
rect 3650 1380 3700 1390
rect 4450 1380 5100 1390
rect 5950 1380 6200 1390
rect 6300 1380 6800 1390
rect 7400 1380 7450 1390
rect 7800 1380 7850 1390
rect 450 1370 800 1380
rect 1000 1370 1050 1380
rect 2050 1370 2100 1380
rect 3000 1370 3050 1380
rect 3500 1370 3550 1380
rect 3650 1370 3700 1380
rect 4450 1370 5100 1380
rect 5950 1370 6200 1380
rect 6300 1370 6800 1380
rect 7400 1370 7450 1380
rect 7800 1370 7850 1380
rect 450 1360 800 1370
rect 1000 1360 1050 1370
rect 2050 1360 2100 1370
rect 3000 1360 3050 1370
rect 3500 1360 3550 1370
rect 3650 1360 3700 1370
rect 4450 1360 5100 1370
rect 5950 1360 6200 1370
rect 6300 1360 6800 1370
rect 7400 1360 7450 1370
rect 7800 1360 7850 1370
rect 450 1350 800 1360
rect 1000 1350 1050 1360
rect 2050 1350 2100 1360
rect 3000 1350 3050 1360
rect 3500 1350 3550 1360
rect 3650 1350 3700 1360
rect 4450 1350 5100 1360
rect 5950 1350 6200 1360
rect 6300 1350 6800 1360
rect 7400 1350 7450 1360
rect 7800 1350 7850 1360
rect 450 1340 800 1350
rect 950 1340 1050 1350
rect 2050 1340 2100 1350
rect 2850 1340 3000 1350
rect 3450 1340 3500 1350
rect 3700 1340 3750 1350
rect 4450 1340 4950 1350
rect 5950 1340 6200 1350
rect 6300 1340 6800 1350
rect 7400 1340 7450 1350
rect 7800 1340 7850 1350
rect 450 1330 800 1340
rect 950 1330 1050 1340
rect 2050 1330 2100 1340
rect 2850 1330 3000 1340
rect 3450 1330 3500 1340
rect 3700 1330 3750 1340
rect 4450 1330 4950 1340
rect 5950 1330 6200 1340
rect 6300 1330 6800 1340
rect 7400 1330 7450 1340
rect 7800 1330 7850 1340
rect 450 1320 800 1330
rect 950 1320 1050 1330
rect 2050 1320 2100 1330
rect 2850 1320 3000 1330
rect 3450 1320 3500 1330
rect 3700 1320 3750 1330
rect 4450 1320 4950 1330
rect 5950 1320 6200 1330
rect 6300 1320 6800 1330
rect 7400 1320 7450 1330
rect 7800 1320 7850 1330
rect 450 1310 800 1320
rect 950 1310 1050 1320
rect 2050 1310 2100 1320
rect 2850 1310 3000 1320
rect 3450 1310 3500 1320
rect 3700 1310 3750 1320
rect 4450 1310 4950 1320
rect 5950 1310 6200 1320
rect 6300 1310 6800 1320
rect 7400 1310 7450 1320
rect 7800 1310 7850 1320
rect 450 1300 800 1310
rect 950 1300 1050 1310
rect 2050 1300 2100 1310
rect 2850 1300 3000 1310
rect 3450 1300 3500 1310
rect 3700 1300 3750 1310
rect 4450 1300 4950 1310
rect 5950 1300 6200 1310
rect 6300 1300 6800 1310
rect 7400 1300 7450 1310
rect 7800 1300 7850 1310
rect 400 1290 800 1300
rect 950 1290 1050 1300
rect 2050 1290 2150 1300
rect 2800 1290 2900 1300
rect 3450 1290 3500 1300
rect 3750 1290 3800 1300
rect 4450 1290 4950 1300
rect 5950 1290 6250 1300
rect 6300 1290 6800 1300
rect 7400 1290 7450 1300
rect 7800 1290 7850 1300
rect 400 1280 800 1290
rect 950 1280 1050 1290
rect 2050 1280 2150 1290
rect 2800 1280 2900 1290
rect 3450 1280 3500 1290
rect 3750 1280 3800 1290
rect 4450 1280 4950 1290
rect 5950 1280 6250 1290
rect 6300 1280 6800 1290
rect 7400 1280 7450 1290
rect 7800 1280 7850 1290
rect 400 1270 800 1280
rect 950 1270 1050 1280
rect 2050 1270 2150 1280
rect 2800 1270 2900 1280
rect 3450 1270 3500 1280
rect 3750 1270 3800 1280
rect 4450 1270 4950 1280
rect 5950 1270 6250 1280
rect 6300 1270 6800 1280
rect 7400 1270 7450 1280
rect 7800 1270 7850 1280
rect 400 1260 800 1270
rect 950 1260 1050 1270
rect 2050 1260 2150 1270
rect 2800 1260 2900 1270
rect 3450 1260 3500 1270
rect 3750 1260 3800 1270
rect 4450 1260 4950 1270
rect 5950 1260 6250 1270
rect 6300 1260 6800 1270
rect 7400 1260 7450 1270
rect 7800 1260 7850 1270
rect 400 1250 800 1260
rect 950 1250 1050 1260
rect 2050 1250 2150 1260
rect 2800 1250 2900 1260
rect 3450 1250 3500 1260
rect 3750 1250 3800 1260
rect 4450 1250 4950 1260
rect 5950 1250 6250 1260
rect 6300 1250 6800 1260
rect 7400 1250 7450 1260
rect 7800 1250 7850 1260
rect 400 1240 800 1250
rect 950 1240 1000 1250
rect 2000 1240 2100 1250
rect 2700 1240 2800 1250
rect 3450 1240 3500 1250
rect 3850 1240 3900 1250
rect 4150 1240 4200 1250
rect 4500 1240 4750 1250
rect 5950 1240 6250 1250
rect 6300 1240 6700 1250
rect 7400 1240 7450 1250
rect 400 1230 800 1240
rect 950 1230 1000 1240
rect 2000 1230 2100 1240
rect 2700 1230 2800 1240
rect 3450 1230 3500 1240
rect 3850 1230 3900 1240
rect 4150 1230 4200 1240
rect 4500 1230 4750 1240
rect 5950 1230 6250 1240
rect 6300 1230 6700 1240
rect 7400 1230 7450 1240
rect 400 1220 800 1230
rect 950 1220 1000 1230
rect 2000 1220 2100 1230
rect 2700 1220 2800 1230
rect 3450 1220 3500 1230
rect 3850 1220 3900 1230
rect 4150 1220 4200 1230
rect 4500 1220 4750 1230
rect 5950 1220 6250 1230
rect 6300 1220 6700 1230
rect 7400 1220 7450 1230
rect 400 1210 800 1220
rect 950 1210 1000 1220
rect 2000 1210 2100 1220
rect 2700 1210 2800 1220
rect 3450 1210 3500 1220
rect 3850 1210 3900 1220
rect 4150 1210 4200 1220
rect 4500 1210 4750 1220
rect 5950 1210 6250 1220
rect 6300 1210 6700 1220
rect 7400 1210 7450 1220
rect 400 1200 800 1210
rect 950 1200 1000 1210
rect 2000 1200 2100 1210
rect 2700 1200 2800 1210
rect 3450 1200 3500 1210
rect 3850 1200 3900 1210
rect 4150 1200 4200 1210
rect 4500 1200 4750 1210
rect 5950 1200 6250 1210
rect 6300 1200 6700 1210
rect 7400 1200 7450 1210
rect 400 1190 750 1200
rect 900 1190 1000 1200
rect 2000 1190 2050 1200
rect 2600 1190 2850 1200
rect 3500 1190 3550 1200
rect 3900 1190 3950 1200
rect 4150 1190 4200 1200
rect 4500 1190 4550 1200
rect 5950 1190 6250 1200
rect 6350 1190 6600 1200
rect 7400 1190 7450 1200
rect 7850 1190 7900 1200
rect 400 1180 750 1190
rect 900 1180 1000 1190
rect 2000 1180 2050 1190
rect 2600 1180 2850 1190
rect 3500 1180 3550 1190
rect 3900 1180 3950 1190
rect 4150 1180 4200 1190
rect 4500 1180 4550 1190
rect 5950 1180 6250 1190
rect 6350 1180 6600 1190
rect 7400 1180 7450 1190
rect 7850 1180 7900 1190
rect 400 1170 750 1180
rect 900 1170 1000 1180
rect 2000 1170 2050 1180
rect 2600 1170 2850 1180
rect 3500 1170 3550 1180
rect 3900 1170 3950 1180
rect 4150 1170 4200 1180
rect 4500 1170 4550 1180
rect 5950 1170 6250 1180
rect 6350 1170 6600 1180
rect 7400 1170 7450 1180
rect 7850 1170 7900 1180
rect 400 1160 750 1170
rect 900 1160 1000 1170
rect 2000 1160 2050 1170
rect 2600 1160 2850 1170
rect 3500 1160 3550 1170
rect 3900 1160 3950 1170
rect 4150 1160 4200 1170
rect 4500 1160 4550 1170
rect 5950 1160 6250 1170
rect 6350 1160 6600 1170
rect 7400 1160 7450 1170
rect 7850 1160 7900 1170
rect 400 1150 750 1160
rect 900 1150 1000 1160
rect 2000 1150 2050 1160
rect 2600 1150 2850 1160
rect 3500 1150 3550 1160
rect 3900 1150 3950 1160
rect 4150 1150 4200 1160
rect 4500 1150 4550 1160
rect 5950 1150 6250 1160
rect 6350 1150 6600 1160
rect 7400 1150 7450 1160
rect 7850 1150 7900 1160
rect 350 1140 650 1150
rect 700 1140 750 1150
rect 900 1140 1000 1150
rect 1500 1140 1650 1150
rect 2400 1140 2550 1150
rect 2800 1140 2900 1150
rect 3550 1140 3600 1150
rect 4150 1140 4200 1150
rect 4500 1140 4550 1150
rect 4900 1140 5350 1150
rect 5950 1140 6300 1150
rect 6400 1140 6500 1150
rect 7850 1140 7900 1150
rect 350 1130 650 1140
rect 700 1130 750 1140
rect 900 1130 1000 1140
rect 1500 1130 1650 1140
rect 2400 1130 2550 1140
rect 2800 1130 2900 1140
rect 3550 1130 3600 1140
rect 4150 1130 4200 1140
rect 4500 1130 4550 1140
rect 4900 1130 5350 1140
rect 5950 1130 6300 1140
rect 6400 1130 6500 1140
rect 7850 1130 7900 1140
rect 350 1120 650 1130
rect 700 1120 750 1130
rect 900 1120 1000 1130
rect 1500 1120 1650 1130
rect 2400 1120 2550 1130
rect 2800 1120 2900 1130
rect 3550 1120 3600 1130
rect 4150 1120 4200 1130
rect 4500 1120 4550 1130
rect 4900 1120 5350 1130
rect 5950 1120 6300 1130
rect 6400 1120 6500 1130
rect 7850 1120 7900 1130
rect 350 1110 650 1120
rect 700 1110 750 1120
rect 900 1110 1000 1120
rect 1500 1110 1650 1120
rect 2400 1110 2550 1120
rect 2800 1110 2900 1120
rect 3550 1110 3600 1120
rect 4150 1110 4200 1120
rect 4500 1110 4550 1120
rect 4900 1110 5350 1120
rect 5950 1110 6300 1120
rect 6400 1110 6500 1120
rect 7850 1110 7900 1120
rect 350 1100 650 1110
rect 700 1100 750 1110
rect 900 1100 1000 1110
rect 1500 1100 1650 1110
rect 2400 1100 2550 1110
rect 2800 1100 2900 1110
rect 3550 1100 3600 1110
rect 4150 1100 4200 1110
rect 4500 1100 4550 1110
rect 4900 1100 5350 1110
rect 5950 1100 6300 1110
rect 6400 1100 6500 1110
rect 7850 1100 7900 1110
rect 350 1090 650 1100
rect 700 1090 750 1100
rect 900 1090 1000 1100
rect 1450 1090 1500 1100
rect 1650 1090 1700 1100
rect 1950 1090 2000 1100
rect 2850 1090 2900 1100
rect 3600 1090 3650 1100
rect 4050 1090 4100 1100
rect 4150 1090 4200 1100
rect 4650 1090 5450 1100
rect 5700 1090 5800 1100
rect 6000 1090 6300 1100
rect 6400 1090 6450 1100
rect 7850 1090 7900 1100
rect 350 1080 650 1090
rect 700 1080 750 1090
rect 900 1080 1000 1090
rect 1450 1080 1500 1090
rect 1650 1080 1700 1090
rect 1950 1080 2000 1090
rect 2850 1080 2900 1090
rect 3600 1080 3650 1090
rect 4050 1080 4100 1090
rect 4150 1080 4200 1090
rect 4650 1080 5450 1090
rect 5700 1080 5800 1090
rect 6000 1080 6300 1090
rect 6400 1080 6450 1090
rect 7850 1080 7900 1090
rect 350 1070 650 1080
rect 700 1070 750 1080
rect 900 1070 1000 1080
rect 1450 1070 1500 1080
rect 1650 1070 1700 1080
rect 1950 1070 2000 1080
rect 2850 1070 2900 1080
rect 3600 1070 3650 1080
rect 4050 1070 4100 1080
rect 4150 1070 4200 1080
rect 4650 1070 5450 1080
rect 5700 1070 5800 1080
rect 6000 1070 6300 1080
rect 6400 1070 6450 1080
rect 7850 1070 7900 1080
rect 350 1060 650 1070
rect 700 1060 750 1070
rect 900 1060 1000 1070
rect 1450 1060 1500 1070
rect 1650 1060 1700 1070
rect 1950 1060 2000 1070
rect 2850 1060 2900 1070
rect 3600 1060 3650 1070
rect 4050 1060 4100 1070
rect 4150 1060 4200 1070
rect 4650 1060 5450 1070
rect 5700 1060 5800 1070
rect 6000 1060 6300 1070
rect 6400 1060 6450 1070
rect 7850 1060 7900 1070
rect 350 1050 650 1060
rect 700 1050 750 1060
rect 900 1050 1000 1060
rect 1450 1050 1500 1060
rect 1650 1050 1700 1060
rect 1950 1050 2000 1060
rect 2850 1050 2900 1060
rect 3600 1050 3650 1060
rect 4050 1050 4100 1060
rect 4150 1050 4200 1060
rect 4650 1050 5450 1060
rect 5700 1050 5800 1060
rect 6000 1050 6300 1060
rect 6400 1050 6450 1060
rect 7850 1050 7900 1060
rect 300 1040 700 1050
rect 850 1040 1000 1050
rect 1400 1040 1450 1050
rect 1650 1040 1700 1050
rect 1950 1040 2000 1050
rect 2850 1040 2900 1050
rect 3650 1040 3700 1050
rect 4150 1040 4200 1050
rect 4750 1040 5450 1050
rect 5650 1040 5800 1050
rect 5950 1040 6300 1050
rect 6350 1040 6400 1050
rect 300 1030 700 1040
rect 850 1030 1000 1040
rect 1400 1030 1450 1040
rect 1650 1030 1700 1040
rect 1950 1030 2000 1040
rect 2850 1030 2900 1040
rect 3650 1030 3700 1040
rect 4150 1030 4200 1040
rect 4750 1030 5450 1040
rect 5650 1030 5800 1040
rect 5950 1030 6300 1040
rect 6350 1030 6400 1040
rect 300 1020 700 1030
rect 850 1020 1000 1030
rect 1400 1020 1450 1030
rect 1650 1020 1700 1030
rect 1950 1020 2000 1030
rect 2850 1020 2900 1030
rect 3650 1020 3700 1030
rect 4150 1020 4200 1030
rect 4750 1020 5450 1030
rect 5650 1020 5800 1030
rect 5950 1020 6300 1030
rect 6350 1020 6400 1030
rect 300 1010 700 1020
rect 850 1010 1000 1020
rect 1400 1010 1450 1020
rect 1650 1010 1700 1020
rect 1950 1010 2000 1020
rect 2850 1010 2900 1020
rect 3650 1010 3700 1020
rect 4150 1010 4200 1020
rect 4750 1010 5450 1020
rect 5650 1010 5800 1020
rect 5950 1010 6300 1020
rect 6350 1010 6400 1020
rect 300 1000 700 1010
rect 850 1000 1000 1010
rect 1400 1000 1450 1010
rect 1650 1000 1700 1010
rect 1950 1000 2000 1010
rect 2850 1000 2900 1010
rect 3650 1000 3700 1010
rect 4150 1000 4200 1010
rect 4750 1000 5450 1010
rect 5650 1000 5800 1010
rect 5950 1000 6300 1010
rect 6350 1000 6400 1010
rect 300 990 700 1000
rect 850 990 950 1000
rect 1350 990 1400 1000
rect 1550 990 1650 1000
rect 1950 990 2000 1000
rect 2850 990 2900 1000
rect 3700 990 3750 1000
rect 4850 990 5300 1000
rect 6000 990 6400 1000
rect 300 980 700 990
rect 850 980 950 990
rect 1350 980 1400 990
rect 1550 980 1650 990
rect 1950 980 2000 990
rect 2850 980 2900 990
rect 3700 980 3750 990
rect 4850 980 5300 990
rect 6000 980 6400 990
rect 300 970 700 980
rect 850 970 950 980
rect 1350 970 1400 980
rect 1550 970 1650 980
rect 1950 970 2000 980
rect 2850 970 2900 980
rect 3700 970 3750 980
rect 4850 970 5300 980
rect 6000 970 6400 980
rect 300 960 700 970
rect 850 960 950 970
rect 1350 960 1400 970
rect 1550 960 1650 970
rect 1950 960 2000 970
rect 2850 960 2900 970
rect 3700 960 3750 970
rect 4850 960 5300 970
rect 6000 960 6400 970
rect 300 950 700 960
rect 850 950 950 960
rect 1350 950 1400 960
rect 1550 950 1650 960
rect 1950 950 2000 960
rect 2850 950 2900 960
rect 3700 950 3750 960
rect 4850 950 5300 960
rect 6000 950 6400 960
rect 250 940 650 950
rect 850 940 950 950
rect 1250 940 1300 950
rect 1500 940 1600 950
rect 1950 940 2000 950
rect 2800 940 2850 950
rect 3750 940 3800 950
rect 4850 940 5300 950
rect 6050 940 6200 950
rect 6300 940 6400 950
rect 7900 940 7950 950
rect 8950 940 9050 950
rect 250 930 650 940
rect 850 930 950 940
rect 1250 930 1300 940
rect 1500 930 1600 940
rect 1950 930 2000 940
rect 2800 930 2850 940
rect 3750 930 3800 940
rect 4850 930 5300 940
rect 6050 930 6200 940
rect 6300 930 6400 940
rect 7900 930 7950 940
rect 8950 930 9050 940
rect 250 920 650 930
rect 850 920 950 930
rect 1250 920 1300 930
rect 1500 920 1600 930
rect 1950 920 2000 930
rect 2800 920 2850 930
rect 3750 920 3800 930
rect 4850 920 5300 930
rect 6050 920 6200 930
rect 6300 920 6400 930
rect 7900 920 7950 930
rect 8950 920 9050 930
rect 250 910 650 920
rect 850 910 950 920
rect 1250 910 1300 920
rect 1500 910 1600 920
rect 1950 910 2000 920
rect 2800 910 2850 920
rect 3750 910 3800 920
rect 4850 910 5300 920
rect 6050 910 6200 920
rect 6300 910 6400 920
rect 7900 910 7950 920
rect 8950 910 9050 920
rect 250 900 650 910
rect 850 900 950 910
rect 1250 900 1300 910
rect 1500 900 1600 910
rect 1950 900 2000 910
rect 2800 900 2850 910
rect 3750 900 3800 910
rect 4850 900 5300 910
rect 6050 900 6200 910
rect 6300 900 6400 910
rect 7900 900 7950 910
rect 8950 900 9050 910
rect 250 890 650 900
rect 900 890 950 900
rect 1200 890 1250 900
rect 1450 890 1550 900
rect 1950 890 2000 900
rect 2750 890 2800 900
rect 5100 890 5150 900
rect 5200 890 5300 900
rect 6050 890 6200 900
rect 6350 890 6400 900
rect 7900 890 7950 900
rect 8900 890 9050 900
rect 250 880 650 890
rect 900 880 950 890
rect 1200 880 1250 890
rect 1450 880 1550 890
rect 1950 880 2000 890
rect 2750 880 2800 890
rect 5100 880 5150 890
rect 5200 880 5300 890
rect 6050 880 6200 890
rect 6350 880 6400 890
rect 7900 880 7950 890
rect 8900 880 9050 890
rect 250 870 650 880
rect 900 870 950 880
rect 1200 870 1250 880
rect 1450 870 1550 880
rect 1950 870 2000 880
rect 2750 870 2800 880
rect 5100 870 5150 880
rect 5200 870 5300 880
rect 6050 870 6200 880
rect 6350 870 6400 880
rect 7900 870 7950 880
rect 8900 870 9050 880
rect 250 860 650 870
rect 900 860 950 870
rect 1200 860 1250 870
rect 1450 860 1550 870
rect 1950 860 2000 870
rect 2750 860 2800 870
rect 5100 860 5150 870
rect 5200 860 5300 870
rect 6050 860 6200 870
rect 6350 860 6400 870
rect 7900 860 7950 870
rect 8900 860 9050 870
rect 250 850 650 860
rect 900 850 950 860
rect 1200 850 1250 860
rect 1450 850 1550 860
rect 1950 850 2000 860
rect 2750 850 2800 860
rect 5100 850 5150 860
rect 5200 850 5300 860
rect 6050 850 6200 860
rect 6350 850 6400 860
rect 7900 850 7950 860
rect 8900 850 9050 860
rect 200 840 600 850
rect 900 840 950 850
rect 1150 840 1200 850
rect 1400 840 1500 850
rect 2650 840 2700 850
rect 3800 840 3850 850
rect 4900 840 4950 850
rect 5200 840 5350 850
rect 5600 840 5750 850
rect 6050 840 6150 850
rect 6300 840 6350 850
rect 6400 840 6450 850
rect 7900 840 7950 850
rect 8900 840 9050 850
rect 200 830 600 840
rect 900 830 950 840
rect 1150 830 1200 840
rect 1400 830 1500 840
rect 2650 830 2700 840
rect 3800 830 3850 840
rect 4900 830 4950 840
rect 5200 830 5350 840
rect 5600 830 5750 840
rect 6050 830 6150 840
rect 6300 830 6350 840
rect 6400 830 6450 840
rect 7900 830 7950 840
rect 8900 830 9050 840
rect 200 820 600 830
rect 900 820 950 830
rect 1150 820 1200 830
rect 1400 820 1500 830
rect 2650 820 2700 830
rect 3800 820 3850 830
rect 4900 820 4950 830
rect 5200 820 5350 830
rect 5600 820 5750 830
rect 6050 820 6150 830
rect 6300 820 6350 830
rect 6400 820 6450 830
rect 7900 820 7950 830
rect 8900 820 9050 830
rect 200 810 600 820
rect 900 810 950 820
rect 1150 810 1200 820
rect 1400 810 1500 820
rect 2650 810 2700 820
rect 3800 810 3850 820
rect 4900 810 4950 820
rect 5200 810 5350 820
rect 5600 810 5750 820
rect 6050 810 6150 820
rect 6300 810 6350 820
rect 6400 810 6450 820
rect 7900 810 7950 820
rect 8900 810 9050 820
rect 200 800 600 810
rect 900 800 950 810
rect 1150 800 1200 810
rect 1400 800 1500 810
rect 2650 800 2700 810
rect 3800 800 3850 810
rect 4900 800 4950 810
rect 5200 800 5350 810
rect 5600 800 5750 810
rect 6050 800 6150 810
rect 6300 800 6350 810
rect 6400 800 6450 810
rect 7900 800 7950 810
rect 8900 800 9050 810
rect 150 790 600 800
rect 850 790 950 800
rect 1050 790 1100 800
rect 1350 790 1500 800
rect 2000 790 2050 800
rect 2600 790 2650 800
rect 3400 790 3550 800
rect 5200 790 5450 800
rect 5550 790 5750 800
rect 6300 790 6350 800
rect 6400 790 6450 800
rect 7400 790 7450 800
rect 8150 790 8200 800
rect 8850 790 9150 800
rect 150 780 600 790
rect 850 780 950 790
rect 1050 780 1100 790
rect 1350 780 1500 790
rect 2000 780 2050 790
rect 2600 780 2650 790
rect 3400 780 3550 790
rect 5200 780 5450 790
rect 5550 780 5750 790
rect 6300 780 6350 790
rect 6400 780 6450 790
rect 7400 780 7450 790
rect 8150 780 8200 790
rect 8850 780 9150 790
rect 150 770 600 780
rect 850 770 950 780
rect 1050 770 1100 780
rect 1350 770 1500 780
rect 2000 770 2050 780
rect 2600 770 2650 780
rect 3400 770 3550 780
rect 5200 770 5450 780
rect 5550 770 5750 780
rect 6300 770 6350 780
rect 6400 770 6450 780
rect 7400 770 7450 780
rect 8150 770 8200 780
rect 8850 770 9150 780
rect 150 760 600 770
rect 850 760 950 770
rect 1050 760 1100 770
rect 1350 760 1500 770
rect 2000 760 2050 770
rect 2600 760 2650 770
rect 3400 760 3550 770
rect 5200 760 5450 770
rect 5550 760 5750 770
rect 6300 760 6350 770
rect 6400 760 6450 770
rect 7400 760 7450 770
rect 8150 760 8200 770
rect 8850 760 9150 770
rect 150 750 600 760
rect 850 750 950 760
rect 1050 750 1100 760
rect 1350 750 1500 760
rect 2000 750 2050 760
rect 2600 750 2650 760
rect 3400 750 3550 760
rect 5200 750 5450 760
rect 5550 750 5750 760
rect 6300 750 6350 760
rect 6400 750 6450 760
rect 7400 750 7450 760
rect 8150 750 8200 760
rect 8850 750 9150 760
rect 100 740 600 750
rect 800 740 900 750
rect 1000 740 1050 750
rect 1300 740 1450 750
rect 2500 740 2550 750
rect 3300 740 3350 750
rect 5150 740 5200 750
rect 5400 740 5500 750
rect 5550 740 5750 750
rect 6300 740 6350 750
rect 6400 740 6450 750
rect 7400 740 7450 750
rect 8150 740 8200 750
rect 8800 740 9150 750
rect 100 730 600 740
rect 800 730 900 740
rect 1000 730 1050 740
rect 1300 730 1450 740
rect 2500 730 2550 740
rect 3300 730 3350 740
rect 5150 730 5200 740
rect 5400 730 5500 740
rect 5550 730 5750 740
rect 6300 730 6350 740
rect 6400 730 6450 740
rect 7400 730 7450 740
rect 8150 730 8200 740
rect 8800 730 9150 740
rect 100 720 600 730
rect 800 720 900 730
rect 1000 720 1050 730
rect 1300 720 1450 730
rect 2500 720 2550 730
rect 3300 720 3350 730
rect 5150 720 5200 730
rect 5400 720 5500 730
rect 5550 720 5750 730
rect 6300 720 6350 730
rect 6400 720 6450 730
rect 7400 720 7450 730
rect 8150 720 8200 730
rect 8800 720 9150 730
rect 100 710 600 720
rect 800 710 900 720
rect 1000 710 1050 720
rect 1300 710 1450 720
rect 2500 710 2550 720
rect 3300 710 3350 720
rect 5150 710 5200 720
rect 5400 710 5500 720
rect 5550 710 5750 720
rect 6300 710 6350 720
rect 6400 710 6450 720
rect 7400 710 7450 720
rect 8150 710 8200 720
rect 8800 710 9150 720
rect 100 700 600 710
rect 800 700 900 710
rect 1000 700 1050 710
rect 1300 700 1450 710
rect 2500 700 2550 710
rect 3300 700 3350 710
rect 5150 700 5200 710
rect 5400 700 5500 710
rect 5550 700 5750 710
rect 6300 700 6350 710
rect 6400 700 6450 710
rect 7400 700 7450 710
rect 8150 700 8200 710
rect 8800 700 9150 710
rect 0 690 550 700
rect 900 690 950 700
rect 1300 690 1400 700
rect 2050 690 2100 700
rect 2400 690 2450 700
rect 3200 690 3250 700
rect 4950 690 5000 700
rect 5150 690 5200 700
rect 5400 690 5500 700
rect 5700 690 5750 700
rect 6300 690 6350 700
rect 6450 690 6500 700
rect 7400 690 7450 700
rect 7950 690 8000 700
rect 8150 690 8250 700
rect 8750 690 9100 700
rect 0 680 550 690
rect 900 680 950 690
rect 1300 680 1400 690
rect 2050 680 2100 690
rect 2400 680 2450 690
rect 3200 680 3250 690
rect 4950 680 5000 690
rect 5150 680 5200 690
rect 5400 680 5500 690
rect 5700 680 5750 690
rect 6300 680 6350 690
rect 6450 680 6500 690
rect 7400 680 7450 690
rect 7950 680 8000 690
rect 8150 680 8250 690
rect 8750 680 9100 690
rect 0 670 550 680
rect 900 670 950 680
rect 1300 670 1400 680
rect 2050 670 2100 680
rect 2400 670 2450 680
rect 3200 670 3250 680
rect 4950 670 5000 680
rect 5150 670 5200 680
rect 5400 670 5500 680
rect 5700 670 5750 680
rect 6300 670 6350 680
rect 6450 670 6500 680
rect 7400 670 7450 680
rect 7950 670 8000 680
rect 8150 670 8250 680
rect 8750 670 9100 680
rect 0 660 550 670
rect 900 660 950 670
rect 1300 660 1400 670
rect 2050 660 2100 670
rect 2400 660 2450 670
rect 3200 660 3250 670
rect 4950 660 5000 670
rect 5150 660 5200 670
rect 5400 660 5500 670
rect 5700 660 5750 670
rect 6300 660 6350 670
rect 6450 660 6500 670
rect 7400 660 7450 670
rect 7950 660 8000 670
rect 8150 660 8250 670
rect 8750 660 9100 670
rect 0 650 550 660
rect 900 650 950 660
rect 1300 650 1400 660
rect 2050 650 2100 660
rect 2400 650 2450 660
rect 3200 650 3250 660
rect 4950 650 5000 660
rect 5150 650 5200 660
rect 5400 650 5500 660
rect 5700 650 5750 660
rect 6300 650 6350 660
rect 6450 650 6500 660
rect 7400 650 7450 660
rect 7950 650 8000 660
rect 8150 650 8250 660
rect 8750 650 9100 660
rect 0 640 350 650
rect 1350 640 1450 650
rect 2050 640 2100 650
rect 3050 640 3100 650
rect 4950 640 5000 650
rect 5400 640 5450 650
rect 5500 640 5550 650
rect 5700 640 5750 650
rect 6300 640 6350 650
rect 7400 640 7450 650
rect 8150 640 8300 650
rect 8750 640 9100 650
rect 0 630 350 640
rect 1350 630 1450 640
rect 2050 630 2100 640
rect 3050 630 3100 640
rect 4950 630 5000 640
rect 5400 630 5450 640
rect 5500 630 5550 640
rect 5700 630 5750 640
rect 6300 630 6350 640
rect 7400 630 7450 640
rect 8150 630 8300 640
rect 8750 630 9100 640
rect 0 620 350 630
rect 1350 620 1450 630
rect 2050 620 2100 630
rect 3050 620 3100 630
rect 4950 620 5000 630
rect 5400 620 5450 630
rect 5500 620 5550 630
rect 5700 620 5750 630
rect 6300 620 6350 630
rect 7400 620 7450 630
rect 8150 620 8300 630
rect 8750 620 9100 630
rect 0 610 350 620
rect 1350 610 1450 620
rect 2050 610 2100 620
rect 3050 610 3100 620
rect 4950 610 5000 620
rect 5400 610 5450 620
rect 5500 610 5550 620
rect 5700 610 5750 620
rect 6300 610 6350 620
rect 7400 610 7450 620
rect 8150 610 8300 620
rect 8750 610 9100 620
rect 0 600 350 610
rect 1350 600 1450 610
rect 2050 600 2100 610
rect 3050 600 3100 610
rect 4950 600 5000 610
rect 5400 600 5450 610
rect 5500 600 5550 610
rect 5700 600 5750 610
rect 6300 600 6350 610
rect 7400 600 7450 610
rect 8150 600 8300 610
rect 8750 600 9100 610
rect 0 590 300 600
rect 1450 590 1500 600
rect 2250 590 2300 600
rect 2950 590 3000 600
rect 5550 590 5600 600
rect 5700 590 5850 600
rect 6500 590 6550 600
rect 7400 590 7450 600
rect 8000 590 8050 600
rect 8150 590 8350 600
rect 8700 590 9050 600
rect 0 580 300 590
rect 1450 580 1500 590
rect 2250 580 2300 590
rect 2950 580 3000 590
rect 5550 580 5600 590
rect 5700 580 5850 590
rect 6500 580 6550 590
rect 7400 580 7450 590
rect 8000 580 8050 590
rect 8150 580 8350 590
rect 8700 580 9050 590
rect 0 570 300 580
rect 1450 570 1500 580
rect 2250 570 2300 580
rect 2950 570 3000 580
rect 5550 570 5600 580
rect 5700 570 5850 580
rect 6500 570 6550 580
rect 7400 570 7450 580
rect 8000 570 8050 580
rect 8150 570 8350 580
rect 8700 570 9050 580
rect 0 560 300 570
rect 1450 560 1500 570
rect 2250 560 2300 570
rect 2950 560 3000 570
rect 5550 560 5600 570
rect 5700 560 5850 570
rect 6500 560 6550 570
rect 7400 560 7450 570
rect 8000 560 8050 570
rect 8150 560 8350 570
rect 8700 560 9050 570
rect 0 550 300 560
rect 1450 550 1500 560
rect 2250 550 2300 560
rect 2950 550 3000 560
rect 5550 550 5600 560
rect 5700 550 5850 560
rect 6500 550 6550 560
rect 7400 550 7450 560
rect 8000 550 8050 560
rect 8150 550 8350 560
rect 8700 550 9050 560
rect 0 540 150 550
rect 2150 540 2200 550
rect 2800 540 2850 550
rect 5400 540 5500 550
rect 5600 540 5850 550
rect 6550 540 6600 550
rect 7400 540 7450 550
rect 8050 540 8450 550
rect 8550 540 9050 550
rect 0 530 150 540
rect 2150 530 2200 540
rect 2800 530 2850 540
rect 5400 530 5500 540
rect 5600 530 5850 540
rect 6550 530 6600 540
rect 7400 530 7450 540
rect 8050 530 8450 540
rect 8550 530 9050 540
rect 0 520 150 530
rect 2150 520 2200 530
rect 2800 520 2850 530
rect 5400 520 5500 530
rect 5600 520 5850 530
rect 6550 520 6600 530
rect 7400 520 7450 530
rect 8050 520 8450 530
rect 8550 520 9050 530
rect 0 510 150 520
rect 2150 510 2200 520
rect 2800 510 2850 520
rect 5400 510 5500 520
rect 5600 510 5850 520
rect 6550 510 6600 520
rect 7400 510 7450 520
rect 8050 510 8450 520
rect 8550 510 9050 520
rect 0 500 150 510
rect 2150 500 2200 510
rect 2800 500 2850 510
rect 5400 500 5500 510
rect 5600 500 5850 510
rect 6550 500 6600 510
rect 7400 500 7450 510
rect 8050 500 8450 510
rect 8550 500 9050 510
rect 0 490 100 500
rect 650 490 900 500
rect 1550 490 1750 500
rect 1800 490 2000 500
rect 2250 490 2350 500
rect 2550 490 2700 500
rect 4350 490 4550 500
rect 5400 490 5450 500
rect 5650 490 5800 500
rect 6300 490 6350 500
rect 6550 490 6600 500
rect 7400 490 7450 500
rect 8100 490 9000 500
rect 0 480 100 490
rect 650 480 900 490
rect 1550 480 1750 490
rect 1800 480 2000 490
rect 2250 480 2350 490
rect 2550 480 2700 490
rect 4350 480 4550 490
rect 5400 480 5450 490
rect 5650 480 5800 490
rect 6300 480 6350 490
rect 6550 480 6600 490
rect 7400 480 7450 490
rect 8100 480 9000 490
rect 0 470 100 480
rect 650 470 900 480
rect 1550 470 1750 480
rect 1800 470 2000 480
rect 2250 470 2350 480
rect 2550 470 2700 480
rect 4350 470 4550 480
rect 5400 470 5450 480
rect 5650 470 5800 480
rect 6300 470 6350 480
rect 6550 470 6600 480
rect 7400 470 7450 480
rect 8100 470 9000 480
rect 0 460 100 470
rect 650 460 900 470
rect 1550 460 1750 470
rect 1800 460 2000 470
rect 2250 460 2350 470
rect 2550 460 2700 470
rect 4350 460 4550 470
rect 5400 460 5450 470
rect 5650 460 5800 470
rect 6300 460 6350 470
rect 6550 460 6600 470
rect 7400 460 7450 470
rect 8100 460 9000 470
rect 0 450 100 460
rect 650 450 900 460
rect 1550 450 1750 460
rect 1800 450 2000 460
rect 2250 450 2350 460
rect 2550 450 2700 460
rect 4350 450 4550 460
rect 5400 450 5450 460
rect 5650 450 5800 460
rect 6300 450 6350 460
rect 6550 450 6600 460
rect 7400 450 7450 460
rect 8100 450 9000 460
rect 0 440 50 450
rect 750 440 1000 450
rect 4300 440 4550 450
rect 4650 440 4700 450
rect 5700 440 5800 450
rect 5900 440 5950 450
rect 6300 440 6350 450
rect 6600 440 6650 450
rect 7350 440 7450 450
rect 8200 440 8950 450
rect 0 430 50 440
rect 750 430 1000 440
rect 4300 430 4550 440
rect 4650 430 4700 440
rect 5700 430 5800 440
rect 5900 430 5950 440
rect 6300 430 6350 440
rect 6600 430 6650 440
rect 7350 430 7450 440
rect 8200 430 8950 440
rect 0 420 50 430
rect 750 420 1000 430
rect 4300 420 4550 430
rect 4650 420 4700 430
rect 5700 420 5800 430
rect 5900 420 5950 430
rect 6300 420 6350 430
rect 6600 420 6650 430
rect 7350 420 7450 430
rect 8200 420 8950 430
rect 0 410 50 420
rect 750 410 1000 420
rect 4300 410 4550 420
rect 4650 410 4700 420
rect 5700 410 5800 420
rect 5900 410 5950 420
rect 6300 410 6350 420
rect 6600 410 6650 420
rect 7350 410 7450 420
rect 8200 410 8950 420
rect 0 400 50 410
rect 750 400 1000 410
rect 4300 400 4550 410
rect 4650 400 4700 410
rect 5700 400 5800 410
rect 5900 400 5950 410
rect 6300 400 6350 410
rect 6600 400 6650 410
rect 7350 400 7450 410
rect 8200 400 8950 410
rect 700 390 1050 400
rect 4400 390 4550 400
rect 4600 390 4700 400
rect 5200 390 5250 400
rect 5300 390 5400 400
rect 5750 390 5800 400
rect 5850 390 5950 400
rect 6300 390 6350 400
rect 6600 390 6700 400
rect 7350 390 7450 400
rect 8250 390 8800 400
rect 8850 390 8950 400
rect 700 380 1050 390
rect 4400 380 4550 390
rect 4600 380 4700 390
rect 5200 380 5250 390
rect 5300 380 5400 390
rect 5750 380 5800 390
rect 5850 380 5950 390
rect 6300 380 6350 390
rect 6600 380 6700 390
rect 7350 380 7450 390
rect 8250 380 8800 390
rect 8850 380 8950 390
rect 700 370 1050 380
rect 4400 370 4550 380
rect 4600 370 4700 380
rect 5200 370 5250 380
rect 5300 370 5400 380
rect 5750 370 5800 380
rect 5850 370 5950 380
rect 6300 370 6350 380
rect 6600 370 6700 380
rect 7350 370 7450 380
rect 8250 370 8800 380
rect 8850 370 8950 380
rect 700 360 1050 370
rect 4400 360 4550 370
rect 4600 360 4700 370
rect 5200 360 5250 370
rect 5300 360 5400 370
rect 5750 360 5800 370
rect 5850 360 5950 370
rect 6300 360 6350 370
rect 6600 360 6700 370
rect 7350 360 7450 370
rect 8250 360 8800 370
rect 8850 360 8950 370
rect 700 350 1050 360
rect 4400 350 4550 360
rect 4600 350 4700 360
rect 5200 350 5250 360
rect 5300 350 5400 360
rect 5750 350 5800 360
rect 5850 350 5950 360
rect 6300 350 6350 360
rect 6600 350 6700 360
rect 7350 350 7450 360
rect 8250 350 8800 360
rect 8850 350 8950 360
rect 800 340 1000 350
rect 4600 340 4650 350
rect 5000 340 5050 350
rect 5700 340 6000 350
rect 6300 340 6350 350
rect 6650 340 6700 350
rect 7350 340 7450 350
rect 8300 340 8800 350
rect 8850 340 9000 350
rect 800 330 1000 340
rect 4600 330 4650 340
rect 5000 330 5050 340
rect 5700 330 6000 340
rect 6300 330 6350 340
rect 6650 330 6700 340
rect 7350 330 7450 340
rect 8300 330 8800 340
rect 8850 330 9000 340
rect 800 320 1000 330
rect 4600 320 4650 330
rect 5000 320 5050 330
rect 5700 320 6000 330
rect 6300 320 6350 330
rect 6650 320 6700 330
rect 7350 320 7450 330
rect 8300 320 8800 330
rect 8850 320 9000 330
rect 800 310 1000 320
rect 4600 310 4650 320
rect 5000 310 5050 320
rect 5700 310 6000 320
rect 6300 310 6350 320
rect 6650 310 6700 320
rect 7350 310 7450 320
rect 8300 310 8800 320
rect 8850 310 9000 320
rect 800 300 1000 310
rect 4600 300 4650 310
rect 5000 300 5050 310
rect 5700 300 6000 310
rect 6300 300 6350 310
rect 6650 300 6700 310
rect 7350 300 7450 310
rect 8300 300 8800 310
rect 8850 300 9000 310
rect 5000 290 5050 300
rect 5700 290 6000 300
rect 6300 290 6350 300
rect 6700 290 6750 300
rect 7350 290 7450 300
rect 8350 290 8850 300
rect 8950 290 9000 300
rect 5000 280 5050 290
rect 5700 280 6000 290
rect 6300 280 6350 290
rect 6700 280 6750 290
rect 7350 280 7450 290
rect 8350 280 8850 290
rect 8950 280 9000 290
rect 5000 270 5050 280
rect 5700 270 6000 280
rect 6300 270 6350 280
rect 6700 270 6750 280
rect 7350 270 7450 280
rect 8350 270 8850 280
rect 8950 270 9000 280
rect 5000 260 5050 270
rect 5700 260 6000 270
rect 6300 260 6350 270
rect 6700 260 6750 270
rect 7350 260 7450 270
rect 8350 260 8850 270
rect 8950 260 9000 270
rect 5000 250 5050 260
rect 5700 250 6000 260
rect 6300 250 6350 260
rect 6700 250 6750 260
rect 7350 250 7450 260
rect 8350 250 8850 260
rect 8950 250 9000 260
rect 5950 240 6100 250
rect 6300 240 6400 250
rect 6750 240 6800 250
rect 7350 240 7400 250
rect 8400 240 8850 250
rect 5950 230 6100 240
rect 6300 230 6400 240
rect 6750 230 6800 240
rect 7350 230 7400 240
rect 8400 230 8850 240
rect 5950 220 6100 230
rect 6300 220 6400 230
rect 6750 220 6800 230
rect 7350 220 7400 230
rect 8400 220 8850 230
rect 5950 210 6100 220
rect 6300 210 6400 220
rect 6750 210 6800 220
rect 7350 210 7400 220
rect 8400 210 8850 220
rect 5950 200 6100 210
rect 6300 200 6400 210
rect 6750 200 6800 210
rect 7350 200 7400 210
rect 8400 200 8850 210
rect 150 190 200 200
rect 5350 190 5700 200
rect 5950 190 6050 200
rect 6350 190 6400 200
rect 6800 190 6900 200
rect 7350 190 7400 200
rect 8450 190 8550 200
rect 8750 190 8800 200
rect 150 180 200 190
rect 5350 180 5700 190
rect 5950 180 6050 190
rect 6350 180 6400 190
rect 6800 180 6900 190
rect 7350 180 7400 190
rect 8450 180 8550 190
rect 8750 180 8800 190
rect 150 170 200 180
rect 5350 170 5700 180
rect 5950 170 6050 180
rect 6350 170 6400 180
rect 6800 170 6900 180
rect 7350 170 7400 180
rect 8450 170 8550 180
rect 8750 170 8800 180
rect 150 160 200 170
rect 5350 160 5700 170
rect 5950 160 6050 170
rect 6350 160 6400 170
rect 6800 160 6900 170
rect 7350 160 7400 170
rect 8450 160 8550 170
rect 8750 160 8800 170
rect 150 150 200 160
rect 5350 150 5700 160
rect 5950 150 6050 160
rect 6350 150 6400 160
rect 6800 150 6900 160
rect 7350 150 7400 160
rect 8450 150 8550 160
rect 8750 150 8800 160
rect 350 140 500 150
rect 5050 140 5100 150
rect 5350 140 5950 150
rect 6350 140 6450 150
rect 6800 140 7000 150
rect 7350 140 7400 150
rect 8500 140 8550 150
rect 8950 140 9050 150
rect 9200 140 9300 150
rect 9800 140 9850 150
rect 350 130 500 140
rect 5050 130 5100 140
rect 5350 130 5950 140
rect 6350 130 6450 140
rect 6800 130 7000 140
rect 7350 130 7400 140
rect 8500 130 8550 140
rect 8950 130 9050 140
rect 9200 130 9300 140
rect 9800 130 9850 140
rect 350 120 500 130
rect 5050 120 5100 130
rect 5350 120 5950 130
rect 6350 120 6450 130
rect 6800 120 7000 130
rect 7350 120 7400 130
rect 8500 120 8550 130
rect 8950 120 9050 130
rect 9200 120 9300 130
rect 9800 120 9850 130
rect 350 110 500 120
rect 5050 110 5100 120
rect 5350 110 5950 120
rect 6350 110 6450 120
rect 6800 110 7000 120
rect 7350 110 7400 120
rect 8500 110 8550 120
rect 8950 110 9050 120
rect 9200 110 9300 120
rect 9800 110 9850 120
rect 350 100 500 110
rect 5050 100 5100 110
rect 5350 100 5950 110
rect 6350 100 6450 110
rect 6800 100 7000 110
rect 7350 100 7400 110
rect 8500 100 8550 110
rect 8950 100 9050 110
rect 9200 100 9300 110
rect 9800 100 9850 110
rect 200 90 250 100
rect 350 90 400 100
rect 500 90 600 100
rect 750 90 800 100
rect 4350 90 4450 100
rect 5050 90 5100 100
rect 5350 90 5850 100
rect 6000 90 6050 100
rect 6400 90 6450 100
rect 6800 90 7050 100
rect 7350 90 7400 100
rect 8550 90 8600 100
rect 9200 90 9350 100
rect 9800 90 9850 100
rect 200 80 250 90
rect 350 80 400 90
rect 500 80 600 90
rect 750 80 800 90
rect 4350 80 4450 90
rect 5050 80 5100 90
rect 5350 80 5850 90
rect 6000 80 6050 90
rect 6400 80 6450 90
rect 6800 80 7050 90
rect 7350 80 7400 90
rect 8550 80 8600 90
rect 9200 80 9350 90
rect 9800 80 9850 90
rect 200 70 250 80
rect 350 70 400 80
rect 500 70 600 80
rect 750 70 800 80
rect 4350 70 4450 80
rect 5050 70 5100 80
rect 5350 70 5850 80
rect 6000 70 6050 80
rect 6400 70 6450 80
rect 6800 70 7050 80
rect 7350 70 7400 80
rect 8550 70 8600 80
rect 9200 70 9350 80
rect 9800 70 9850 80
rect 200 60 250 70
rect 350 60 400 70
rect 500 60 600 70
rect 750 60 800 70
rect 4350 60 4450 70
rect 5050 60 5100 70
rect 5350 60 5850 70
rect 6000 60 6050 70
rect 6400 60 6450 70
rect 6800 60 7050 70
rect 7350 60 7400 70
rect 8550 60 8600 70
rect 9200 60 9350 70
rect 9800 60 9850 70
rect 200 50 250 60
rect 350 50 400 60
rect 500 50 600 60
rect 750 50 800 60
rect 4350 50 4450 60
rect 5050 50 5100 60
rect 5350 50 5850 60
rect 6000 50 6050 60
rect 6400 50 6450 60
rect 6800 50 7050 60
rect 7350 50 7400 60
rect 8550 50 8600 60
rect 9200 50 9350 60
rect 9800 50 9850 60
rect 200 40 350 50
rect 600 40 650 50
rect 750 40 850 50
rect 4400 40 4550 50
rect 5350 40 5700 50
rect 5800 40 6050 50
rect 6450 40 6500 50
rect 6850 40 7100 50
rect 7350 40 7400 50
rect 8950 40 9000 50
rect 9200 40 9250 50
rect 9350 40 9450 50
rect 9800 40 9900 50
rect 200 30 350 40
rect 600 30 650 40
rect 750 30 850 40
rect 4400 30 4550 40
rect 5350 30 5700 40
rect 5800 30 6050 40
rect 6450 30 6500 40
rect 6850 30 7100 40
rect 7350 30 7400 40
rect 8950 30 9000 40
rect 9200 30 9250 40
rect 9350 30 9450 40
rect 9800 30 9900 40
rect 200 20 350 30
rect 600 20 650 30
rect 750 20 850 30
rect 4400 20 4550 30
rect 5350 20 5700 30
rect 5800 20 6050 30
rect 6450 20 6500 30
rect 6850 20 7100 30
rect 7350 20 7400 30
rect 8950 20 9000 30
rect 9200 20 9250 30
rect 9350 20 9450 30
rect 9800 20 9900 30
rect 200 10 350 20
rect 600 10 650 20
rect 750 10 850 20
rect 4400 10 4550 20
rect 5350 10 5700 20
rect 5800 10 6050 20
rect 6450 10 6500 20
rect 6850 10 7100 20
rect 7350 10 7400 20
rect 8950 10 9000 20
rect 9200 10 9250 20
rect 9350 10 9450 20
rect 9800 10 9900 20
rect 200 0 350 10
rect 600 0 650 10
rect 750 0 850 10
rect 4400 0 4550 10
rect 5350 0 5700 10
rect 5800 0 6050 10
rect 6450 0 6500 10
rect 6850 0 7100 10
rect 7350 0 7400 10
rect 8950 0 9000 10
rect 9200 0 9250 10
rect 9350 0 9450 10
rect 9800 0 9900 10
<< metal2 >>
rect 3600 7440 3650 7450
rect 9650 7440 9750 7450
rect 9950 7440 9990 7450
rect 3600 7430 3650 7440
rect 9650 7430 9750 7440
rect 9950 7430 9990 7440
rect 3600 7420 3650 7430
rect 9650 7420 9750 7430
rect 9950 7420 9990 7430
rect 3600 7410 3650 7420
rect 9650 7410 9750 7420
rect 9950 7410 9990 7420
rect 3600 7400 3650 7410
rect 9650 7400 9750 7410
rect 9950 7400 9990 7410
rect 3300 7390 3350 7400
rect 9950 7390 9990 7400
rect 3300 7380 3350 7390
rect 9950 7380 9990 7390
rect 3300 7370 3350 7380
rect 9950 7370 9990 7380
rect 3300 7360 3350 7370
rect 9950 7360 9990 7370
rect 3300 7350 3350 7360
rect 9950 7350 9990 7360
rect 2050 7340 2100 7350
rect 9650 7340 9750 7350
rect 9800 7340 9850 7350
rect 9950 7340 9990 7350
rect 2050 7330 2100 7340
rect 9650 7330 9750 7340
rect 9800 7330 9850 7340
rect 9950 7330 9990 7340
rect 2050 7320 2100 7330
rect 9650 7320 9750 7330
rect 9800 7320 9850 7330
rect 9950 7320 9990 7330
rect 2050 7310 2100 7320
rect 9650 7310 9750 7320
rect 9800 7310 9850 7320
rect 9950 7310 9990 7320
rect 2050 7300 2100 7310
rect 9650 7300 9750 7310
rect 9800 7300 9850 7310
rect 9950 7300 9990 7310
rect 2000 7290 2050 7300
rect 9650 7290 9800 7300
rect 9900 7290 9990 7300
rect 2000 7280 2050 7290
rect 9650 7280 9800 7290
rect 9900 7280 9990 7290
rect 2000 7270 2050 7280
rect 9650 7270 9800 7280
rect 9900 7270 9990 7280
rect 2000 7260 2050 7270
rect 9650 7260 9800 7270
rect 9900 7260 9990 7270
rect 2000 7250 2050 7260
rect 9650 7250 9800 7260
rect 9900 7250 9990 7260
rect 3350 7240 3400 7250
rect 9800 7240 9900 7250
rect 9950 7240 9990 7250
rect 3350 7230 3400 7240
rect 9800 7230 9900 7240
rect 9950 7230 9990 7240
rect 3350 7220 3400 7230
rect 9800 7220 9900 7230
rect 9950 7220 9990 7230
rect 3350 7210 3400 7220
rect 9800 7210 9900 7220
rect 9950 7210 9990 7220
rect 3350 7200 3400 7210
rect 9800 7200 9900 7210
rect 9950 7200 9990 7210
rect 1950 7190 2000 7200
rect 3850 7190 3900 7200
rect 9650 7190 9850 7200
rect 9950 7190 9990 7200
rect 1950 7180 2000 7190
rect 3850 7180 3900 7190
rect 9650 7180 9850 7190
rect 9950 7180 9990 7190
rect 1950 7170 2000 7180
rect 3850 7170 3900 7180
rect 9650 7170 9850 7180
rect 9950 7170 9990 7180
rect 1950 7160 2000 7170
rect 3850 7160 3900 7170
rect 9650 7160 9850 7170
rect 9950 7160 9990 7170
rect 1950 7150 2000 7160
rect 3850 7150 3900 7160
rect 9650 7150 9850 7160
rect 9950 7150 9990 7160
rect 3350 7140 3400 7150
rect 3850 7140 3900 7150
rect 9650 7140 9850 7150
rect 3350 7130 3400 7140
rect 3850 7130 3900 7140
rect 9650 7130 9850 7140
rect 3350 7120 3400 7130
rect 3850 7120 3900 7130
rect 9650 7120 9850 7130
rect 3350 7110 3400 7120
rect 3850 7110 3900 7120
rect 9650 7110 9850 7120
rect 3350 7100 3400 7110
rect 3850 7100 3900 7110
rect 9650 7100 9850 7110
rect 1950 7090 2100 7100
rect 3450 7090 3500 7100
rect 3650 7090 3700 7100
rect 3850 7090 3900 7100
rect 9600 7090 9800 7100
rect 1950 7080 2100 7090
rect 3450 7080 3500 7090
rect 3650 7080 3700 7090
rect 3850 7080 3900 7090
rect 9600 7080 9800 7090
rect 1950 7070 2100 7080
rect 3450 7070 3500 7080
rect 3650 7070 3700 7080
rect 3850 7070 3900 7080
rect 9600 7070 9800 7080
rect 1950 7060 2100 7070
rect 3450 7060 3500 7070
rect 3650 7060 3700 7070
rect 3850 7060 3900 7070
rect 9600 7060 9800 7070
rect 1950 7050 2100 7060
rect 3450 7050 3500 7060
rect 3650 7050 3700 7060
rect 3850 7050 3900 7060
rect 9600 7050 9800 7060
rect 1950 7040 2100 7050
rect 2250 7040 2400 7050
rect 2850 7040 2900 7050
rect 3000 7040 3100 7050
rect 3500 7040 3550 7050
rect 3650 7040 3700 7050
rect 9650 7040 9700 7050
rect 1950 7030 2100 7040
rect 2250 7030 2400 7040
rect 2850 7030 2900 7040
rect 3000 7030 3100 7040
rect 3500 7030 3550 7040
rect 3650 7030 3700 7040
rect 9650 7030 9700 7040
rect 1950 7020 2100 7030
rect 2250 7020 2400 7030
rect 2850 7020 2900 7030
rect 3000 7020 3100 7030
rect 3500 7020 3550 7030
rect 3650 7020 3700 7030
rect 9650 7020 9700 7030
rect 1950 7010 2100 7020
rect 2250 7010 2400 7020
rect 2850 7010 2900 7020
rect 3000 7010 3100 7020
rect 3500 7010 3550 7020
rect 3650 7010 3700 7020
rect 9650 7010 9700 7020
rect 1950 7000 2100 7010
rect 2250 7000 2400 7010
rect 2850 7000 2900 7010
rect 3000 7000 3100 7010
rect 3500 7000 3550 7010
rect 3650 7000 3700 7010
rect 9650 7000 9700 7010
rect 1950 6990 2000 7000
rect 2250 6990 3150 7000
rect 3300 6990 3350 7000
rect 3550 6990 3600 7000
rect 1950 6980 2000 6990
rect 2250 6980 3150 6990
rect 3300 6980 3350 6990
rect 3550 6980 3600 6990
rect 1950 6970 2000 6980
rect 2250 6970 3150 6980
rect 3300 6970 3350 6980
rect 3550 6970 3600 6980
rect 1950 6960 2000 6970
rect 2250 6960 3150 6970
rect 3300 6960 3350 6970
rect 3550 6960 3600 6970
rect 1950 6950 2000 6960
rect 2250 6950 3150 6960
rect 3300 6950 3350 6960
rect 3550 6950 3600 6960
rect 2300 6940 2400 6950
rect 2650 6940 2750 6950
rect 3450 6940 3500 6950
rect 3650 6940 3750 6950
rect 9650 6940 9700 6950
rect 2300 6930 2400 6940
rect 2650 6930 2750 6940
rect 3450 6930 3500 6940
rect 3650 6930 3750 6940
rect 9650 6930 9700 6940
rect 2300 6920 2400 6930
rect 2650 6920 2750 6930
rect 3450 6920 3500 6930
rect 3650 6920 3750 6930
rect 9650 6920 9700 6930
rect 2300 6910 2400 6920
rect 2650 6910 2750 6920
rect 3450 6910 3500 6920
rect 3650 6910 3750 6920
rect 9650 6910 9700 6920
rect 2300 6900 2400 6910
rect 2650 6900 2750 6910
rect 3450 6900 3500 6910
rect 3650 6900 3750 6910
rect 9650 6900 9700 6910
rect 1900 6890 1950 6900
rect 2350 6890 2500 6900
rect 3550 6890 3600 6900
rect 3750 6890 3800 6900
rect 9650 6890 9700 6900
rect 1900 6880 1950 6890
rect 2350 6880 2500 6890
rect 3550 6880 3600 6890
rect 3750 6880 3800 6890
rect 9650 6880 9700 6890
rect 1900 6870 1950 6880
rect 2350 6870 2500 6880
rect 3550 6870 3600 6880
rect 3750 6870 3800 6880
rect 9650 6870 9700 6880
rect 1900 6860 1950 6870
rect 2350 6860 2500 6870
rect 3550 6860 3600 6870
rect 3750 6860 3800 6870
rect 9650 6860 9700 6870
rect 1900 6850 1950 6860
rect 2350 6850 2500 6860
rect 3550 6850 3600 6860
rect 3750 6850 3800 6860
rect 9650 6850 9700 6860
rect 2450 6840 2550 6850
rect 3800 6840 3850 6850
rect 9650 6840 9700 6850
rect 2450 6830 2550 6840
rect 3800 6830 3850 6840
rect 9650 6830 9700 6840
rect 2450 6820 2550 6830
rect 3800 6820 3850 6830
rect 9650 6820 9700 6830
rect 2450 6810 2550 6820
rect 3800 6810 3850 6820
rect 9650 6810 9700 6820
rect 2450 6800 2550 6810
rect 3800 6800 3850 6810
rect 9650 6800 9700 6810
rect 1950 6790 2000 6800
rect 2300 6790 2450 6800
rect 2650 6790 2800 6800
rect 3700 6790 3750 6800
rect 3850 6790 3900 6800
rect 9600 6790 9700 6800
rect 1950 6780 2000 6790
rect 2300 6780 2450 6790
rect 2650 6780 2800 6790
rect 3700 6780 3750 6790
rect 3850 6780 3900 6790
rect 9600 6780 9700 6790
rect 1950 6770 2000 6780
rect 2300 6770 2450 6780
rect 2650 6770 2800 6780
rect 3700 6770 3750 6780
rect 3850 6770 3900 6780
rect 9600 6770 9700 6780
rect 1950 6760 2000 6770
rect 2300 6760 2450 6770
rect 2650 6760 2800 6770
rect 3700 6760 3750 6770
rect 3850 6760 3900 6770
rect 9600 6760 9700 6770
rect 1950 6750 2000 6760
rect 2300 6750 2450 6760
rect 2650 6750 2800 6760
rect 3700 6750 3750 6760
rect 3850 6750 3900 6760
rect 9600 6750 9700 6760
rect 2500 6740 2550 6750
rect 3050 6740 3200 6750
rect 3850 6740 3900 6750
rect 9600 6740 9700 6750
rect 2500 6730 2550 6740
rect 3050 6730 3200 6740
rect 3850 6730 3900 6740
rect 9600 6730 9700 6740
rect 2500 6720 2550 6730
rect 3050 6720 3200 6730
rect 3850 6720 3900 6730
rect 9600 6720 9700 6730
rect 2500 6710 2550 6720
rect 3050 6710 3200 6720
rect 3850 6710 3900 6720
rect 9600 6710 9700 6720
rect 2500 6700 2550 6710
rect 3050 6700 3200 6710
rect 3850 6700 3900 6710
rect 9600 6700 9700 6710
rect 2200 6690 2250 6700
rect 2550 6690 2600 6700
rect 3350 6690 3450 6700
rect 3900 6690 3950 6700
rect 9650 6690 9700 6700
rect 9850 6690 9900 6700
rect 2200 6680 2250 6690
rect 2550 6680 2600 6690
rect 3350 6680 3450 6690
rect 3900 6680 3950 6690
rect 9650 6680 9700 6690
rect 9850 6680 9900 6690
rect 2200 6670 2250 6680
rect 2550 6670 2600 6680
rect 3350 6670 3450 6680
rect 3900 6670 3950 6680
rect 9650 6670 9700 6680
rect 9850 6670 9900 6680
rect 2200 6660 2250 6670
rect 2550 6660 2600 6670
rect 3350 6660 3450 6670
rect 3900 6660 3950 6670
rect 9650 6660 9700 6670
rect 9850 6660 9900 6670
rect 2200 6650 2250 6660
rect 2550 6650 2600 6660
rect 3350 6650 3450 6660
rect 3900 6650 3950 6660
rect 9650 6650 9700 6660
rect 9850 6650 9900 6660
rect 1800 6640 1850 6650
rect 2600 6640 2650 6650
rect 3550 6640 3600 6650
rect 3900 6640 3950 6650
rect 9650 6640 9750 6650
rect 1800 6630 1850 6640
rect 2600 6630 2650 6640
rect 3550 6630 3600 6640
rect 3900 6630 3950 6640
rect 9650 6630 9750 6640
rect 1800 6620 1850 6630
rect 2600 6620 2650 6630
rect 3550 6620 3600 6630
rect 3900 6620 3950 6630
rect 9650 6620 9750 6630
rect 1800 6610 1850 6620
rect 2600 6610 2650 6620
rect 3550 6610 3600 6620
rect 3900 6610 3950 6620
rect 9650 6610 9750 6620
rect 1800 6600 1850 6610
rect 2600 6600 2650 6610
rect 3550 6600 3600 6610
rect 3900 6600 3950 6610
rect 9650 6600 9750 6610
rect 2600 6590 2650 6600
rect 3650 6590 3700 6600
rect 2600 6580 2650 6590
rect 3650 6580 3700 6590
rect 2600 6570 2650 6580
rect 3650 6570 3700 6580
rect 2600 6560 2650 6570
rect 3650 6560 3700 6570
rect 2600 6550 2650 6560
rect 3650 6550 3700 6560
rect 1450 6540 1500 6550
rect 1650 6540 1750 6550
rect 1800 6540 1850 6550
rect 3750 6540 3800 6550
rect 1450 6530 1500 6540
rect 1650 6530 1750 6540
rect 1800 6530 1850 6540
rect 3750 6530 3800 6540
rect 1450 6520 1500 6530
rect 1650 6520 1750 6530
rect 1800 6520 1850 6530
rect 3750 6520 3800 6530
rect 1450 6510 1500 6520
rect 1650 6510 1750 6520
rect 1800 6510 1850 6520
rect 3750 6510 3800 6520
rect 1450 6500 1500 6510
rect 1650 6500 1750 6510
rect 1800 6500 1850 6510
rect 3750 6500 3800 6510
rect 1300 6490 1400 6500
rect 1650 6490 1900 6500
rect 2400 6490 2600 6500
rect 3850 6490 3900 6500
rect 6150 6490 6200 6500
rect 6350 6490 6550 6500
rect 9900 6490 9950 6500
rect 1300 6480 1400 6490
rect 1650 6480 1900 6490
rect 2400 6480 2600 6490
rect 3850 6480 3900 6490
rect 6150 6480 6200 6490
rect 6350 6480 6550 6490
rect 9900 6480 9950 6490
rect 1300 6470 1400 6480
rect 1650 6470 1900 6480
rect 2400 6470 2600 6480
rect 3850 6470 3900 6480
rect 6150 6470 6200 6480
rect 6350 6470 6550 6480
rect 9900 6470 9950 6480
rect 1300 6460 1400 6470
rect 1650 6460 1900 6470
rect 2400 6460 2600 6470
rect 3850 6460 3900 6470
rect 6150 6460 6200 6470
rect 6350 6460 6550 6470
rect 9900 6460 9950 6470
rect 1300 6450 1400 6460
rect 1650 6450 1900 6460
rect 2400 6450 2600 6460
rect 3850 6450 3900 6460
rect 6150 6450 6200 6460
rect 6350 6450 6550 6460
rect 9900 6450 9950 6460
rect 1350 6440 1450 6450
rect 1600 6440 1650 6450
rect 1950 6440 2050 6450
rect 2500 6440 2550 6450
rect 6100 6440 6400 6450
rect 6550 6440 6600 6450
rect 9700 6440 9750 6450
rect 9950 6440 9990 6450
rect 1350 6430 1450 6440
rect 1600 6430 1650 6440
rect 1950 6430 2050 6440
rect 2500 6430 2550 6440
rect 6100 6430 6400 6440
rect 6550 6430 6600 6440
rect 9700 6430 9750 6440
rect 9950 6430 9990 6440
rect 1350 6420 1450 6430
rect 1600 6420 1650 6430
rect 1950 6420 2050 6430
rect 2500 6420 2550 6430
rect 6100 6420 6400 6430
rect 6550 6420 6600 6430
rect 9700 6420 9750 6430
rect 9950 6420 9990 6430
rect 1350 6410 1450 6420
rect 1600 6410 1650 6420
rect 1950 6410 2050 6420
rect 2500 6410 2550 6420
rect 6100 6410 6400 6420
rect 6550 6410 6600 6420
rect 9700 6410 9750 6420
rect 9950 6410 9990 6420
rect 1350 6400 1450 6410
rect 1600 6400 1650 6410
rect 1950 6400 2050 6410
rect 2500 6400 2550 6410
rect 6100 6400 6400 6410
rect 6550 6400 6600 6410
rect 9700 6400 9750 6410
rect 9950 6400 9990 6410
rect 2400 6390 2450 6400
rect 4000 6390 4050 6400
rect 6400 6390 6450 6400
rect 6550 6390 6650 6400
rect 9650 6390 9700 6400
rect 9950 6390 9990 6400
rect 2400 6380 2450 6390
rect 4000 6380 4050 6390
rect 6400 6380 6450 6390
rect 6550 6380 6650 6390
rect 9650 6380 9700 6390
rect 9950 6380 9990 6390
rect 2400 6370 2450 6380
rect 4000 6370 4050 6380
rect 6400 6370 6450 6380
rect 6550 6370 6650 6380
rect 9650 6370 9700 6380
rect 9950 6370 9990 6380
rect 2400 6360 2450 6370
rect 4000 6360 4050 6370
rect 6400 6360 6450 6370
rect 6550 6360 6650 6370
rect 9650 6360 9700 6370
rect 9950 6360 9990 6370
rect 2400 6350 2450 6360
rect 4000 6350 4050 6360
rect 6400 6350 6450 6360
rect 6550 6350 6650 6360
rect 9650 6350 9700 6360
rect 9950 6350 9990 6360
rect 1550 6340 1600 6350
rect 1800 6340 1850 6350
rect 2450 6340 2500 6350
rect 6500 6340 6750 6350
rect 9950 6340 9990 6350
rect 1550 6330 1600 6340
rect 1800 6330 1850 6340
rect 2450 6330 2500 6340
rect 6500 6330 6750 6340
rect 9950 6330 9990 6340
rect 1550 6320 1600 6330
rect 1800 6320 1850 6330
rect 2450 6320 2500 6330
rect 6500 6320 6750 6330
rect 9950 6320 9990 6330
rect 1550 6310 1600 6320
rect 1800 6310 1850 6320
rect 2450 6310 2500 6320
rect 6500 6310 6750 6320
rect 9950 6310 9990 6320
rect 1550 6300 1600 6310
rect 1800 6300 1850 6310
rect 2450 6300 2500 6310
rect 6500 6300 6750 6310
rect 9950 6300 9990 6310
rect 1400 6290 1450 6300
rect 1550 6290 1650 6300
rect 2450 6290 2500 6300
rect 5500 6290 5550 6300
rect 6550 6290 6650 6300
rect 6750 6290 6800 6300
rect 9650 6290 9700 6300
rect 9800 6290 9850 6300
rect 1400 6280 1450 6290
rect 1550 6280 1650 6290
rect 2450 6280 2500 6290
rect 5500 6280 5550 6290
rect 6550 6280 6650 6290
rect 6750 6280 6800 6290
rect 9650 6280 9700 6290
rect 9800 6280 9850 6290
rect 1400 6270 1450 6280
rect 1550 6270 1650 6280
rect 2450 6270 2500 6280
rect 5500 6270 5550 6280
rect 6550 6270 6650 6280
rect 6750 6270 6800 6280
rect 9650 6270 9700 6280
rect 9800 6270 9850 6280
rect 1400 6260 1450 6270
rect 1550 6260 1650 6270
rect 2450 6260 2500 6270
rect 5500 6260 5550 6270
rect 6550 6260 6650 6270
rect 6750 6260 6800 6270
rect 9650 6260 9700 6270
rect 9800 6260 9850 6270
rect 1400 6250 1450 6260
rect 1550 6250 1650 6260
rect 2450 6250 2500 6260
rect 5500 6250 5550 6260
rect 6550 6250 6650 6260
rect 6750 6250 6800 6260
rect 9650 6250 9700 6260
rect 9800 6250 9850 6260
rect 1400 6240 1450 6250
rect 1600 6240 1650 6250
rect 5450 6240 5500 6250
rect 6600 6240 6700 6250
rect 6750 6240 6800 6250
rect 9500 6240 9600 6250
rect 9650 6240 9700 6250
rect 1400 6230 1450 6240
rect 1600 6230 1650 6240
rect 5450 6230 5500 6240
rect 6600 6230 6700 6240
rect 6750 6230 6800 6240
rect 9500 6230 9600 6240
rect 9650 6230 9700 6240
rect 1400 6220 1450 6230
rect 1600 6220 1650 6230
rect 5450 6220 5500 6230
rect 6600 6220 6700 6230
rect 6750 6220 6800 6230
rect 9500 6220 9600 6230
rect 9650 6220 9700 6230
rect 1400 6210 1450 6220
rect 1600 6210 1650 6220
rect 5450 6210 5500 6220
rect 6600 6210 6700 6220
rect 6750 6210 6800 6220
rect 9500 6210 9600 6220
rect 9650 6210 9700 6220
rect 1400 6200 1450 6210
rect 1600 6200 1650 6210
rect 5450 6200 5500 6210
rect 6600 6200 6700 6210
rect 6750 6200 6800 6210
rect 9500 6200 9600 6210
rect 9650 6200 9700 6210
rect 1400 6190 1450 6200
rect 1600 6190 1750 6200
rect 5300 6190 5350 6200
rect 5400 6190 5450 6200
rect 6700 6190 6800 6200
rect 9300 6190 9400 6200
rect 1400 6180 1450 6190
rect 1600 6180 1750 6190
rect 5300 6180 5350 6190
rect 5400 6180 5450 6190
rect 6700 6180 6800 6190
rect 9300 6180 9400 6190
rect 1400 6170 1450 6180
rect 1600 6170 1750 6180
rect 5300 6170 5350 6180
rect 5400 6170 5450 6180
rect 6700 6170 6800 6180
rect 9300 6170 9400 6180
rect 1400 6160 1450 6170
rect 1600 6160 1750 6170
rect 5300 6160 5350 6170
rect 5400 6160 5450 6170
rect 6700 6160 6800 6170
rect 9300 6160 9400 6170
rect 1400 6150 1450 6160
rect 1600 6150 1750 6160
rect 5300 6150 5350 6160
rect 5400 6150 5450 6160
rect 6700 6150 6800 6160
rect 9300 6150 9400 6160
rect 1300 6140 1450 6150
rect 1600 6140 1650 6150
rect 3900 6140 3950 6150
rect 4250 6140 4300 6150
rect 6700 6140 6850 6150
rect 9200 6140 9250 6150
rect 9350 6140 9500 6150
rect 9800 6140 9850 6150
rect 1300 6130 1450 6140
rect 1600 6130 1650 6140
rect 3900 6130 3950 6140
rect 4250 6130 4300 6140
rect 6700 6130 6850 6140
rect 9200 6130 9250 6140
rect 9350 6130 9500 6140
rect 9800 6130 9850 6140
rect 1300 6120 1450 6130
rect 1600 6120 1650 6130
rect 3900 6120 3950 6130
rect 4250 6120 4300 6130
rect 6700 6120 6850 6130
rect 9200 6120 9250 6130
rect 9350 6120 9500 6130
rect 9800 6120 9850 6130
rect 1300 6110 1450 6120
rect 1600 6110 1650 6120
rect 3900 6110 3950 6120
rect 4250 6110 4300 6120
rect 6700 6110 6850 6120
rect 9200 6110 9250 6120
rect 9350 6110 9500 6120
rect 9800 6110 9850 6120
rect 1300 6100 1450 6110
rect 1600 6100 1650 6110
rect 3900 6100 3950 6110
rect 4250 6100 4300 6110
rect 6700 6100 6850 6110
rect 9200 6100 9250 6110
rect 9350 6100 9500 6110
rect 9800 6100 9850 6110
rect 1300 6090 1350 6100
rect 1600 6090 1650 6100
rect 2450 6090 2500 6100
rect 3800 6090 3850 6100
rect 5250 6090 5300 6100
rect 6750 6090 6900 6100
rect 9100 6090 9350 6100
rect 1300 6080 1350 6090
rect 1600 6080 1650 6090
rect 2450 6080 2500 6090
rect 3800 6080 3850 6090
rect 5250 6080 5300 6090
rect 6750 6080 6900 6090
rect 9100 6080 9350 6090
rect 1300 6070 1350 6080
rect 1600 6070 1650 6080
rect 2450 6070 2500 6080
rect 3800 6070 3850 6080
rect 5250 6070 5300 6080
rect 6750 6070 6900 6080
rect 9100 6070 9350 6080
rect 1300 6060 1350 6070
rect 1600 6060 1650 6070
rect 2450 6060 2500 6070
rect 3800 6060 3850 6070
rect 5250 6060 5300 6070
rect 6750 6060 6900 6070
rect 9100 6060 9350 6070
rect 1300 6050 1350 6060
rect 1600 6050 1650 6060
rect 2450 6050 2500 6060
rect 3800 6050 3850 6060
rect 5250 6050 5300 6060
rect 6750 6050 6900 6060
rect 9100 6050 9350 6060
rect 1200 6040 1300 6050
rect 1600 6040 1700 6050
rect 3750 6040 3800 6050
rect 4300 6040 4350 6050
rect 5200 6040 5250 6050
rect 6750 6040 6950 6050
rect 8950 6040 9100 6050
rect 9300 6040 9350 6050
rect 1200 6030 1300 6040
rect 1600 6030 1700 6040
rect 3750 6030 3800 6040
rect 4300 6030 4350 6040
rect 5200 6030 5250 6040
rect 6750 6030 6950 6040
rect 8950 6030 9100 6040
rect 9300 6030 9350 6040
rect 1200 6020 1300 6030
rect 1600 6020 1700 6030
rect 3750 6020 3800 6030
rect 4300 6020 4350 6030
rect 5200 6020 5250 6030
rect 6750 6020 6950 6030
rect 8950 6020 9100 6030
rect 9300 6020 9350 6030
rect 1200 6010 1300 6020
rect 1600 6010 1700 6020
rect 3750 6010 3800 6020
rect 4300 6010 4350 6020
rect 5200 6010 5250 6020
rect 6750 6010 6950 6020
rect 8950 6010 9100 6020
rect 9300 6010 9350 6020
rect 1200 6000 1300 6010
rect 1600 6000 1700 6010
rect 3750 6000 3800 6010
rect 4300 6000 4350 6010
rect 5200 6000 5250 6010
rect 6750 6000 6950 6010
rect 8950 6000 9100 6010
rect 9300 6000 9350 6010
rect 1150 5990 1200 6000
rect 1650 5990 1700 6000
rect 3150 5990 3250 6000
rect 4100 5990 4150 6000
rect 4300 5990 4350 6000
rect 6800 5990 6950 6000
rect 8750 5990 8950 6000
rect 9300 5990 9350 6000
rect 9850 5990 9900 6000
rect 1150 5980 1200 5990
rect 1650 5980 1700 5990
rect 3150 5980 3250 5990
rect 4100 5980 4150 5990
rect 4300 5980 4350 5990
rect 6800 5980 6950 5990
rect 8750 5980 8950 5990
rect 9300 5980 9350 5990
rect 9850 5980 9900 5990
rect 1150 5970 1200 5980
rect 1650 5970 1700 5980
rect 3150 5970 3250 5980
rect 4100 5970 4150 5980
rect 4300 5970 4350 5980
rect 6800 5970 6950 5980
rect 8750 5970 8950 5980
rect 9300 5970 9350 5980
rect 9850 5970 9900 5980
rect 1150 5960 1200 5970
rect 1650 5960 1700 5970
rect 3150 5960 3250 5970
rect 4100 5960 4150 5970
rect 4300 5960 4350 5970
rect 6800 5960 6950 5970
rect 8750 5960 8950 5970
rect 9300 5960 9350 5970
rect 9850 5960 9900 5970
rect 1150 5950 1200 5960
rect 1650 5950 1700 5960
rect 3150 5950 3250 5960
rect 4100 5950 4150 5960
rect 4300 5950 4350 5960
rect 6800 5950 6950 5960
rect 8750 5950 8950 5960
rect 9300 5950 9350 5960
rect 9850 5950 9900 5960
rect 950 5940 1050 5950
rect 2550 5940 2600 5950
rect 3100 5940 3150 5950
rect 4200 5940 4300 5950
rect 5150 5940 5200 5950
rect 5300 5940 5350 5950
rect 6800 5940 6850 5950
rect 8600 5940 8800 5950
rect 9300 5940 9350 5950
rect 9500 5940 9550 5950
rect 9850 5940 9900 5950
rect 950 5930 1050 5940
rect 2550 5930 2600 5940
rect 3100 5930 3150 5940
rect 4200 5930 4300 5940
rect 5150 5930 5200 5940
rect 5300 5930 5350 5940
rect 6800 5930 6850 5940
rect 8600 5930 8800 5940
rect 9300 5930 9350 5940
rect 9500 5930 9550 5940
rect 9850 5930 9900 5940
rect 950 5920 1050 5930
rect 2550 5920 2600 5930
rect 3100 5920 3150 5930
rect 4200 5920 4300 5930
rect 5150 5920 5200 5930
rect 5300 5920 5350 5930
rect 6800 5920 6850 5930
rect 8600 5920 8800 5930
rect 9300 5920 9350 5930
rect 9500 5920 9550 5930
rect 9850 5920 9900 5930
rect 950 5910 1050 5920
rect 2550 5910 2600 5920
rect 3100 5910 3150 5920
rect 4200 5910 4300 5920
rect 5150 5910 5200 5920
rect 5300 5910 5350 5920
rect 6800 5910 6850 5920
rect 8600 5910 8800 5920
rect 9300 5910 9350 5920
rect 9500 5910 9550 5920
rect 9850 5910 9900 5920
rect 950 5900 1050 5910
rect 2550 5900 2600 5910
rect 3100 5900 3150 5910
rect 4200 5900 4300 5910
rect 5150 5900 5200 5910
rect 5300 5900 5350 5910
rect 6800 5900 6850 5910
rect 8600 5900 8800 5910
rect 9300 5900 9350 5910
rect 9500 5900 9550 5910
rect 9850 5900 9900 5910
rect 700 5890 750 5900
rect 1750 5890 1800 5900
rect 2600 5890 2650 5900
rect 3000 5890 3050 5900
rect 3250 5890 3300 5900
rect 6800 5890 6850 5900
rect 8400 5890 8500 5900
rect 8600 5890 8650 5900
rect 700 5880 750 5890
rect 1750 5880 1800 5890
rect 2600 5880 2650 5890
rect 3000 5880 3050 5890
rect 3250 5880 3300 5890
rect 6800 5880 6850 5890
rect 8400 5880 8500 5890
rect 8600 5880 8650 5890
rect 700 5870 750 5880
rect 1750 5870 1800 5880
rect 2600 5870 2650 5880
rect 3000 5870 3050 5880
rect 3250 5870 3300 5880
rect 6800 5870 6850 5880
rect 8400 5870 8500 5880
rect 8600 5870 8650 5880
rect 700 5860 750 5870
rect 1750 5860 1800 5870
rect 2600 5860 2650 5870
rect 3000 5860 3050 5870
rect 3250 5860 3300 5870
rect 6800 5860 6850 5870
rect 8400 5860 8500 5870
rect 8600 5860 8650 5870
rect 700 5850 750 5860
rect 1750 5850 1800 5860
rect 2600 5850 2650 5860
rect 3000 5850 3050 5860
rect 3250 5850 3300 5860
rect 6800 5850 6850 5860
rect 8400 5850 8500 5860
rect 8600 5850 8650 5860
rect 650 5840 700 5850
rect 800 5840 1000 5850
rect 2650 5840 2700 5850
rect 2850 5840 3000 5850
rect 3250 5840 3300 5850
rect 3700 5840 3750 5850
rect 5100 5840 5150 5850
rect 6800 5840 6850 5850
rect 6950 5840 7000 5850
rect 8250 5840 8400 5850
rect 8600 5840 8650 5850
rect 8750 5840 8800 5850
rect 9200 5840 9300 5850
rect 650 5830 700 5840
rect 800 5830 1000 5840
rect 2650 5830 2700 5840
rect 2850 5830 3000 5840
rect 3250 5830 3300 5840
rect 3700 5830 3750 5840
rect 5100 5830 5150 5840
rect 6800 5830 6850 5840
rect 6950 5830 7000 5840
rect 8250 5830 8400 5840
rect 8600 5830 8650 5840
rect 8750 5830 8800 5840
rect 9200 5830 9300 5840
rect 650 5820 700 5830
rect 800 5820 1000 5830
rect 2650 5820 2700 5830
rect 2850 5820 3000 5830
rect 3250 5820 3300 5830
rect 3700 5820 3750 5830
rect 5100 5820 5150 5830
rect 6800 5820 6850 5830
rect 6950 5820 7000 5830
rect 8250 5820 8400 5830
rect 8600 5820 8650 5830
rect 8750 5820 8800 5830
rect 9200 5820 9300 5830
rect 650 5810 700 5820
rect 800 5810 1000 5820
rect 2650 5810 2700 5820
rect 2850 5810 3000 5820
rect 3250 5810 3300 5820
rect 3700 5810 3750 5820
rect 5100 5810 5150 5820
rect 6800 5810 6850 5820
rect 6950 5810 7000 5820
rect 8250 5810 8400 5820
rect 8600 5810 8650 5820
rect 8750 5810 8800 5820
rect 9200 5810 9300 5820
rect 650 5800 700 5810
rect 800 5800 1000 5810
rect 2650 5800 2700 5810
rect 2850 5800 3000 5810
rect 3250 5800 3300 5810
rect 3700 5800 3750 5810
rect 5100 5800 5150 5810
rect 6800 5800 6850 5810
rect 6950 5800 7000 5810
rect 8250 5800 8400 5810
rect 8600 5800 8650 5810
rect 8750 5800 8800 5810
rect 9200 5800 9300 5810
rect 2650 5790 2700 5800
rect 2800 5790 2900 5800
rect 3250 5790 3300 5800
rect 3750 5790 3850 5800
rect 8100 5790 8300 5800
rect 8750 5790 8800 5800
rect 8950 5790 9100 5800
rect 9900 5790 9950 5800
rect 2650 5780 2700 5790
rect 2800 5780 2900 5790
rect 3250 5780 3300 5790
rect 3750 5780 3850 5790
rect 8100 5780 8300 5790
rect 8750 5780 8800 5790
rect 8950 5780 9100 5790
rect 9900 5780 9950 5790
rect 2650 5770 2700 5780
rect 2800 5770 2900 5780
rect 3250 5770 3300 5780
rect 3750 5770 3850 5780
rect 8100 5770 8300 5780
rect 8750 5770 8800 5780
rect 8950 5770 9100 5780
rect 9900 5770 9950 5780
rect 2650 5760 2700 5770
rect 2800 5760 2900 5770
rect 3250 5760 3300 5770
rect 3750 5760 3850 5770
rect 8100 5760 8300 5770
rect 8750 5760 8800 5770
rect 8950 5760 9100 5770
rect 9900 5760 9950 5770
rect 2650 5750 2700 5760
rect 2800 5750 2900 5760
rect 3250 5750 3300 5760
rect 3750 5750 3850 5760
rect 8100 5750 8300 5760
rect 8750 5750 8800 5760
rect 8950 5750 9100 5760
rect 9900 5750 9950 5760
rect 800 5740 850 5750
rect 1850 5740 1900 5750
rect 2550 5740 2600 5750
rect 2750 5740 2800 5750
rect 3250 5740 3300 5750
rect 3750 5740 3850 5750
rect 3900 5740 3950 5750
rect 5250 5740 5300 5750
rect 6850 5740 6950 5750
rect 7950 5740 8150 5750
rect 8300 5740 8350 5750
rect 8450 5740 8500 5750
rect 8650 5740 8700 5750
rect 8850 5740 8950 5750
rect 800 5730 850 5740
rect 1850 5730 1900 5740
rect 2550 5730 2600 5740
rect 2750 5730 2800 5740
rect 3250 5730 3300 5740
rect 3750 5730 3850 5740
rect 3900 5730 3950 5740
rect 5250 5730 5300 5740
rect 6850 5730 6950 5740
rect 7950 5730 8150 5740
rect 8300 5730 8350 5740
rect 8450 5730 8500 5740
rect 8650 5730 8700 5740
rect 8850 5730 8950 5740
rect 800 5720 850 5730
rect 1850 5720 1900 5730
rect 2550 5720 2600 5730
rect 2750 5720 2800 5730
rect 3250 5720 3300 5730
rect 3750 5720 3850 5730
rect 3900 5720 3950 5730
rect 5250 5720 5300 5730
rect 6850 5720 6950 5730
rect 7950 5720 8150 5730
rect 8300 5720 8350 5730
rect 8450 5720 8500 5730
rect 8650 5720 8700 5730
rect 8850 5720 8950 5730
rect 800 5710 850 5720
rect 1850 5710 1900 5720
rect 2550 5710 2600 5720
rect 2750 5710 2800 5720
rect 3250 5710 3300 5720
rect 3750 5710 3850 5720
rect 3900 5710 3950 5720
rect 5250 5710 5300 5720
rect 6850 5710 6950 5720
rect 7950 5710 8150 5720
rect 8300 5710 8350 5720
rect 8450 5710 8500 5720
rect 8650 5710 8700 5720
rect 8850 5710 8950 5720
rect 800 5700 850 5710
rect 1850 5700 1900 5710
rect 2550 5700 2600 5710
rect 2750 5700 2800 5710
rect 3250 5700 3300 5710
rect 3750 5700 3850 5710
rect 3900 5700 3950 5710
rect 5250 5700 5300 5710
rect 6850 5700 6950 5710
rect 7950 5700 8150 5710
rect 8300 5700 8350 5710
rect 8450 5700 8500 5710
rect 8650 5700 8700 5710
rect 8850 5700 8950 5710
rect 800 5690 850 5700
rect 1100 5690 1150 5700
rect 1850 5690 1900 5700
rect 2200 5690 2250 5700
rect 2500 5690 2550 5700
rect 2650 5690 2750 5700
rect 3250 5690 3300 5700
rect 3700 5690 3950 5700
rect 5100 5690 5150 5700
rect 5250 5690 5300 5700
rect 6850 5690 6950 5700
rect 7750 5690 7850 5700
rect 7900 5690 7950 5700
rect 8300 5690 8400 5700
rect 8500 5690 8550 5700
rect 8700 5690 8750 5700
rect 9950 5690 9990 5700
rect 800 5680 850 5690
rect 1100 5680 1150 5690
rect 1850 5680 1900 5690
rect 2200 5680 2250 5690
rect 2500 5680 2550 5690
rect 2650 5680 2750 5690
rect 3250 5680 3300 5690
rect 3700 5680 3950 5690
rect 5100 5680 5150 5690
rect 5250 5680 5300 5690
rect 6850 5680 6950 5690
rect 7750 5680 7850 5690
rect 7900 5680 7950 5690
rect 8300 5680 8400 5690
rect 8500 5680 8550 5690
rect 8700 5680 8750 5690
rect 9950 5680 9990 5690
rect 800 5670 850 5680
rect 1100 5670 1150 5680
rect 1850 5670 1900 5680
rect 2200 5670 2250 5680
rect 2500 5670 2550 5680
rect 2650 5670 2750 5680
rect 3250 5670 3300 5680
rect 3700 5670 3950 5680
rect 5100 5670 5150 5680
rect 5250 5670 5300 5680
rect 6850 5670 6950 5680
rect 7750 5670 7850 5680
rect 7900 5670 7950 5680
rect 8300 5670 8400 5680
rect 8500 5670 8550 5680
rect 8700 5670 8750 5680
rect 9950 5670 9990 5680
rect 800 5660 850 5670
rect 1100 5660 1150 5670
rect 1850 5660 1900 5670
rect 2200 5660 2250 5670
rect 2500 5660 2550 5670
rect 2650 5660 2750 5670
rect 3250 5660 3300 5670
rect 3700 5660 3950 5670
rect 5100 5660 5150 5670
rect 5250 5660 5300 5670
rect 6850 5660 6950 5670
rect 7750 5660 7850 5670
rect 7900 5660 7950 5670
rect 8300 5660 8400 5670
rect 8500 5660 8550 5670
rect 8700 5660 8750 5670
rect 9950 5660 9990 5670
rect 800 5650 850 5660
rect 1100 5650 1150 5660
rect 1850 5650 1900 5660
rect 2200 5650 2250 5660
rect 2500 5650 2550 5660
rect 2650 5650 2750 5660
rect 3250 5650 3300 5660
rect 3700 5650 3950 5660
rect 5100 5650 5150 5660
rect 5250 5650 5300 5660
rect 6850 5650 6950 5660
rect 7750 5650 7850 5660
rect 7900 5650 7950 5660
rect 8300 5650 8400 5660
rect 8500 5650 8550 5660
rect 8700 5650 8750 5660
rect 9950 5650 9990 5660
rect 750 5640 800 5650
rect 1900 5640 1950 5650
rect 2200 5640 2250 5650
rect 2500 5640 2550 5650
rect 2600 5640 2700 5650
rect 3250 5640 3300 5650
rect 3700 5640 3800 5650
rect 7700 5640 7800 5650
rect 7950 5640 8000 5650
rect 8500 5640 8550 5650
rect 9000 5640 9050 5650
rect 9950 5640 9990 5650
rect 750 5630 800 5640
rect 1900 5630 1950 5640
rect 2200 5630 2250 5640
rect 2500 5630 2550 5640
rect 2600 5630 2700 5640
rect 3250 5630 3300 5640
rect 3700 5630 3800 5640
rect 7700 5630 7800 5640
rect 7950 5630 8000 5640
rect 8500 5630 8550 5640
rect 9000 5630 9050 5640
rect 9950 5630 9990 5640
rect 750 5620 800 5630
rect 1900 5620 1950 5630
rect 2200 5620 2250 5630
rect 2500 5620 2550 5630
rect 2600 5620 2700 5630
rect 3250 5620 3300 5630
rect 3700 5620 3800 5630
rect 7700 5620 7800 5630
rect 7950 5620 8000 5630
rect 8500 5620 8550 5630
rect 9000 5620 9050 5630
rect 9950 5620 9990 5630
rect 750 5610 800 5620
rect 1900 5610 1950 5620
rect 2200 5610 2250 5620
rect 2500 5610 2550 5620
rect 2600 5610 2700 5620
rect 3250 5610 3300 5620
rect 3700 5610 3800 5620
rect 7700 5610 7800 5620
rect 7950 5610 8000 5620
rect 8500 5610 8550 5620
rect 9000 5610 9050 5620
rect 9950 5610 9990 5620
rect 750 5600 800 5610
rect 1900 5600 1950 5610
rect 2200 5600 2250 5610
rect 2500 5600 2550 5610
rect 2600 5600 2700 5610
rect 3250 5600 3300 5610
rect 3700 5600 3800 5610
rect 7700 5600 7800 5610
rect 7950 5600 8000 5610
rect 8500 5600 8550 5610
rect 9000 5600 9050 5610
rect 9950 5600 9990 5610
rect 1900 5590 1950 5600
rect 2200 5590 2250 5600
rect 2450 5590 2500 5600
rect 2600 5590 2650 5600
rect 3250 5590 3300 5600
rect 3450 5590 3500 5600
rect 3650 5590 3750 5600
rect 5100 5590 5150 5600
rect 5600 5590 5650 5600
rect 5800 5590 5850 5600
rect 6300 5590 6450 5600
rect 6900 5590 6950 5600
rect 7450 5590 7600 5600
rect 7950 5590 8000 5600
rect 8850 5590 8950 5600
rect 1900 5580 1950 5590
rect 2200 5580 2250 5590
rect 2450 5580 2500 5590
rect 2600 5580 2650 5590
rect 3250 5580 3300 5590
rect 3450 5580 3500 5590
rect 3650 5580 3750 5590
rect 5100 5580 5150 5590
rect 5600 5580 5650 5590
rect 5800 5580 5850 5590
rect 6300 5580 6450 5590
rect 6900 5580 6950 5590
rect 7450 5580 7600 5590
rect 7950 5580 8000 5590
rect 8850 5580 8950 5590
rect 1900 5570 1950 5580
rect 2200 5570 2250 5580
rect 2450 5570 2500 5580
rect 2600 5570 2650 5580
rect 3250 5570 3300 5580
rect 3450 5570 3500 5580
rect 3650 5570 3750 5580
rect 5100 5570 5150 5580
rect 5600 5570 5650 5580
rect 5800 5570 5850 5580
rect 6300 5570 6450 5580
rect 6900 5570 6950 5580
rect 7450 5570 7600 5580
rect 7950 5570 8000 5580
rect 8850 5570 8950 5580
rect 1900 5560 1950 5570
rect 2200 5560 2250 5570
rect 2450 5560 2500 5570
rect 2600 5560 2650 5570
rect 3250 5560 3300 5570
rect 3450 5560 3500 5570
rect 3650 5560 3750 5570
rect 5100 5560 5150 5570
rect 5600 5560 5650 5570
rect 5800 5560 5850 5570
rect 6300 5560 6450 5570
rect 6900 5560 6950 5570
rect 7450 5560 7600 5570
rect 7950 5560 8000 5570
rect 8850 5560 8950 5570
rect 1900 5550 1950 5560
rect 2200 5550 2250 5560
rect 2450 5550 2500 5560
rect 2600 5550 2650 5560
rect 3250 5550 3300 5560
rect 3450 5550 3500 5560
rect 3650 5550 3750 5560
rect 5100 5550 5150 5560
rect 5600 5550 5650 5560
rect 5800 5550 5850 5560
rect 6300 5550 6450 5560
rect 6900 5550 6950 5560
rect 7450 5550 7600 5560
rect 7950 5550 8000 5560
rect 8850 5550 8950 5560
rect 1900 5540 1950 5550
rect 2200 5540 2250 5550
rect 2400 5540 2450 5550
rect 2550 5540 2600 5550
rect 3250 5540 3300 5550
rect 3450 5540 3500 5550
rect 5650 5540 5750 5550
rect 5900 5540 5950 5550
rect 6200 5540 6250 5550
rect 6500 5540 6550 5550
rect 6900 5540 6950 5550
rect 7450 5540 7500 5550
rect 7750 5540 7800 5550
rect 7950 5540 8050 5550
rect 8100 5540 8250 5550
rect 8700 5540 8750 5550
rect 9000 5540 9050 5550
rect 9100 5540 9150 5550
rect 1900 5530 1950 5540
rect 2200 5530 2250 5540
rect 2400 5530 2450 5540
rect 2550 5530 2600 5540
rect 3250 5530 3300 5540
rect 3450 5530 3500 5540
rect 5650 5530 5750 5540
rect 5900 5530 5950 5540
rect 6200 5530 6250 5540
rect 6500 5530 6550 5540
rect 6900 5530 6950 5540
rect 7450 5530 7500 5540
rect 7750 5530 7800 5540
rect 7950 5530 8050 5540
rect 8100 5530 8250 5540
rect 8700 5530 8750 5540
rect 9000 5530 9050 5540
rect 9100 5530 9150 5540
rect 1900 5520 1950 5530
rect 2200 5520 2250 5530
rect 2400 5520 2450 5530
rect 2550 5520 2600 5530
rect 3250 5520 3300 5530
rect 3450 5520 3500 5530
rect 5650 5520 5750 5530
rect 5900 5520 5950 5530
rect 6200 5520 6250 5530
rect 6500 5520 6550 5530
rect 6900 5520 6950 5530
rect 7450 5520 7500 5530
rect 7750 5520 7800 5530
rect 7950 5520 8050 5530
rect 8100 5520 8250 5530
rect 8700 5520 8750 5530
rect 9000 5520 9050 5530
rect 9100 5520 9150 5530
rect 1900 5510 1950 5520
rect 2200 5510 2250 5520
rect 2400 5510 2450 5520
rect 2550 5510 2600 5520
rect 3250 5510 3300 5520
rect 3450 5510 3500 5520
rect 5650 5510 5750 5520
rect 5900 5510 5950 5520
rect 6200 5510 6250 5520
rect 6500 5510 6550 5520
rect 6900 5510 6950 5520
rect 7450 5510 7500 5520
rect 7750 5510 7800 5520
rect 7950 5510 8050 5520
rect 8100 5510 8250 5520
rect 8700 5510 8750 5520
rect 9000 5510 9050 5520
rect 9100 5510 9150 5520
rect 1900 5500 1950 5510
rect 2200 5500 2250 5510
rect 2400 5500 2450 5510
rect 2550 5500 2600 5510
rect 3250 5500 3300 5510
rect 3450 5500 3500 5510
rect 5650 5500 5750 5510
rect 5900 5500 5950 5510
rect 6200 5500 6250 5510
rect 6500 5500 6550 5510
rect 6900 5500 6950 5510
rect 7450 5500 7500 5510
rect 7750 5500 7800 5510
rect 7950 5500 8050 5510
rect 8100 5500 8250 5510
rect 8700 5500 8750 5510
rect 9000 5500 9050 5510
rect 9100 5500 9150 5510
rect 450 5490 600 5500
rect 2200 5490 2250 5500
rect 2400 5490 2450 5500
rect 2550 5490 2600 5500
rect 2850 5490 2950 5500
rect 3200 5490 3300 5500
rect 3550 5490 3600 5500
rect 5100 5490 5150 5500
rect 5200 5490 5250 5500
rect 5550 5490 5600 5500
rect 5650 5490 5700 5500
rect 5900 5490 5950 5500
rect 6450 5490 6500 5500
rect 7400 5490 7500 5500
rect 7750 5490 7800 5500
rect 7950 5490 8000 5500
rect 8050 5490 8100 5500
rect 8500 5490 8600 5500
rect 450 5480 600 5490
rect 2200 5480 2250 5490
rect 2400 5480 2450 5490
rect 2550 5480 2600 5490
rect 2850 5480 2950 5490
rect 3200 5480 3300 5490
rect 3550 5480 3600 5490
rect 5100 5480 5150 5490
rect 5200 5480 5250 5490
rect 5550 5480 5600 5490
rect 5650 5480 5700 5490
rect 5900 5480 5950 5490
rect 6450 5480 6500 5490
rect 7400 5480 7500 5490
rect 7750 5480 7800 5490
rect 7950 5480 8000 5490
rect 8050 5480 8100 5490
rect 8500 5480 8600 5490
rect 450 5470 600 5480
rect 2200 5470 2250 5480
rect 2400 5470 2450 5480
rect 2550 5470 2600 5480
rect 2850 5470 2950 5480
rect 3200 5470 3300 5480
rect 3550 5470 3600 5480
rect 5100 5470 5150 5480
rect 5200 5470 5250 5480
rect 5550 5470 5600 5480
rect 5650 5470 5700 5480
rect 5900 5470 5950 5480
rect 6450 5470 6500 5480
rect 7400 5470 7500 5480
rect 7750 5470 7800 5480
rect 7950 5470 8000 5480
rect 8050 5470 8100 5480
rect 8500 5470 8600 5480
rect 450 5460 600 5470
rect 2200 5460 2250 5470
rect 2400 5460 2450 5470
rect 2550 5460 2600 5470
rect 2850 5460 2950 5470
rect 3200 5460 3300 5470
rect 3550 5460 3600 5470
rect 5100 5460 5150 5470
rect 5200 5460 5250 5470
rect 5550 5460 5600 5470
rect 5650 5460 5700 5470
rect 5900 5460 5950 5470
rect 6450 5460 6500 5470
rect 7400 5460 7500 5470
rect 7750 5460 7800 5470
rect 7950 5460 8000 5470
rect 8050 5460 8100 5470
rect 8500 5460 8600 5470
rect 450 5450 600 5460
rect 2200 5450 2250 5460
rect 2400 5450 2450 5460
rect 2550 5450 2600 5460
rect 2850 5450 2950 5460
rect 3200 5450 3300 5460
rect 3550 5450 3600 5460
rect 5100 5450 5150 5460
rect 5200 5450 5250 5460
rect 5550 5450 5600 5460
rect 5650 5450 5700 5460
rect 5900 5450 5950 5460
rect 6450 5450 6500 5460
rect 7400 5450 7500 5460
rect 7750 5450 7800 5460
rect 7950 5450 8000 5460
rect 8050 5450 8100 5460
rect 8500 5450 8600 5460
rect 450 5440 500 5450
rect 1950 5440 2000 5450
rect 2600 5440 2650 5450
rect 2850 5440 2900 5450
rect 2950 5440 3050 5450
rect 3150 5440 3250 5450
rect 5100 5440 5150 5450
rect 5450 5440 5500 5450
rect 5600 5440 5650 5450
rect 5900 5440 5950 5450
rect 6500 5440 6600 5450
rect 7350 5440 7400 5450
rect 7450 5440 7500 5450
rect 7950 5440 8000 5450
rect 9100 5440 9150 5450
rect 9450 5440 9550 5450
rect 450 5430 500 5440
rect 1950 5430 2000 5440
rect 2600 5430 2650 5440
rect 2850 5430 2900 5440
rect 2950 5430 3050 5440
rect 3150 5430 3250 5440
rect 5100 5430 5150 5440
rect 5450 5430 5500 5440
rect 5600 5430 5650 5440
rect 5900 5430 5950 5440
rect 6500 5430 6600 5440
rect 7350 5430 7400 5440
rect 7450 5430 7500 5440
rect 7950 5430 8000 5440
rect 9100 5430 9150 5440
rect 9450 5430 9550 5440
rect 450 5420 500 5430
rect 1950 5420 2000 5430
rect 2600 5420 2650 5430
rect 2850 5420 2900 5430
rect 2950 5420 3050 5430
rect 3150 5420 3250 5430
rect 5100 5420 5150 5430
rect 5450 5420 5500 5430
rect 5600 5420 5650 5430
rect 5900 5420 5950 5430
rect 6500 5420 6600 5430
rect 7350 5420 7400 5430
rect 7450 5420 7500 5430
rect 7950 5420 8000 5430
rect 9100 5420 9150 5430
rect 9450 5420 9550 5430
rect 450 5410 500 5420
rect 1950 5410 2000 5420
rect 2600 5410 2650 5420
rect 2850 5410 2900 5420
rect 2950 5410 3050 5420
rect 3150 5410 3250 5420
rect 5100 5410 5150 5420
rect 5450 5410 5500 5420
rect 5600 5410 5650 5420
rect 5900 5410 5950 5420
rect 6500 5410 6600 5420
rect 7350 5410 7400 5420
rect 7450 5410 7500 5420
rect 7950 5410 8000 5420
rect 9100 5410 9150 5420
rect 9450 5410 9550 5420
rect 450 5400 500 5410
rect 1950 5400 2000 5410
rect 2600 5400 2650 5410
rect 2850 5400 2900 5410
rect 2950 5400 3050 5410
rect 3150 5400 3250 5410
rect 5100 5400 5150 5410
rect 5450 5400 5500 5410
rect 5600 5400 5650 5410
rect 5900 5400 5950 5410
rect 6500 5400 6600 5410
rect 7350 5400 7400 5410
rect 7450 5400 7500 5410
rect 7950 5400 8000 5410
rect 9100 5400 9150 5410
rect 9450 5400 9550 5410
rect 400 5390 450 5400
rect 550 5390 600 5400
rect 1950 5390 2000 5400
rect 2600 5390 2900 5400
rect 5450 5390 5600 5400
rect 5850 5390 5900 5400
rect 6650 5390 6700 5400
rect 7350 5390 7450 5400
rect 7750 5390 7800 5400
rect 7850 5390 8000 5400
rect 8100 5390 8150 5400
rect 8200 5390 8250 5400
rect 8300 5390 8350 5400
rect 9000 5390 9050 5400
rect 9250 5390 9400 5400
rect 9450 5390 9500 5400
rect 400 5380 450 5390
rect 550 5380 600 5390
rect 1950 5380 2000 5390
rect 2600 5380 2900 5390
rect 5450 5380 5600 5390
rect 5850 5380 5900 5390
rect 6650 5380 6700 5390
rect 7350 5380 7450 5390
rect 7750 5380 7800 5390
rect 7850 5380 8000 5390
rect 8100 5380 8150 5390
rect 8200 5380 8250 5390
rect 8300 5380 8350 5390
rect 9000 5380 9050 5390
rect 9250 5380 9400 5390
rect 9450 5380 9500 5390
rect 400 5370 450 5380
rect 550 5370 600 5380
rect 1950 5370 2000 5380
rect 2600 5370 2900 5380
rect 5450 5370 5600 5380
rect 5850 5370 5900 5380
rect 6650 5370 6700 5380
rect 7350 5370 7450 5380
rect 7750 5370 7800 5380
rect 7850 5370 8000 5380
rect 8100 5370 8150 5380
rect 8200 5370 8250 5380
rect 8300 5370 8350 5380
rect 9000 5370 9050 5380
rect 9250 5370 9400 5380
rect 9450 5370 9500 5380
rect 400 5360 450 5370
rect 550 5360 600 5370
rect 1950 5360 2000 5370
rect 2600 5360 2900 5370
rect 5450 5360 5600 5370
rect 5850 5360 5900 5370
rect 6650 5360 6700 5370
rect 7350 5360 7450 5370
rect 7750 5360 7800 5370
rect 7850 5360 8000 5370
rect 8100 5360 8150 5370
rect 8200 5360 8250 5370
rect 8300 5360 8350 5370
rect 9000 5360 9050 5370
rect 9250 5360 9400 5370
rect 9450 5360 9500 5370
rect 400 5350 450 5360
rect 550 5350 600 5360
rect 1950 5350 2000 5360
rect 2600 5350 2900 5360
rect 5450 5350 5600 5360
rect 5850 5350 5900 5360
rect 6650 5350 6700 5360
rect 7350 5350 7450 5360
rect 7750 5350 7800 5360
rect 7850 5350 8000 5360
rect 8100 5350 8150 5360
rect 8200 5350 8250 5360
rect 8300 5350 8350 5360
rect 9000 5350 9050 5360
rect 9250 5350 9400 5360
rect 9450 5350 9500 5360
rect 550 5340 600 5350
rect 2000 5340 2050 5350
rect 2450 5340 2550 5350
rect 2600 5340 2750 5350
rect 3500 5340 3550 5350
rect 5700 5340 5850 5350
rect 6500 5340 6750 5350
rect 7350 5340 7400 5350
rect 7500 5340 7600 5350
rect 7900 5340 8050 5350
rect 8800 5340 8850 5350
rect 9100 5340 9150 5350
rect 9350 5340 9400 5350
rect 9450 5340 9500 5350
rect 9600 5340 9650 5350
rect 550 5330 600 5340
rect 2000 5330 2050 5340
rect 2450 5330 2550 5340
rect 2600 5330 2750 5340
rect 3500 5330 3550 5340
rect 5700 5330 5850 5340
rect 6500 5330 6750 5340
rect 7350 5330 7400 5340
rect 7500 5330 7600 5340
rect 7900 5330 8050 5340
rect 8800 5330 8850 5340
rect 9100 5330 9150 5340
rect 9350 5330 9400 5340
rect 9450 5330 9500 5340
rect 9600 5330 9650 5340
rect 550 5320 600 5330
rect 2000 5320 2050 5330
rect 2450 5320 2550 5330
rect 2600 5320 2750 5330
rect 3500 5320 3550 5330
rect 5700 5320 5850 5330
rect 6500 5320 6750 5330
rect 7350 5320 7400 5330
rect 7500 5320 7600 5330
rect 7900 5320 8050 5330
rect 8800 5320 8850 5330
rect 9100 5320 9150 5330
rect 9350 5320 9400 5330
rect 9450 5320 9500 5330
rect 9600 5320 9650 5330
rect 550 5310 600 5320
rect 2000 5310 2050 5320
rect 2450 5310 2550 5320
rect 2600 5310 2750 5320
rect 3500 5310 3550 5320
rect 5700 5310 5850 5320
rect 6500 5310 6750 5320
rect 7350 5310 7400 5320
rect 7500 5310 7600 5320
rect 7900 5310 8050 5320
rect 8800 5310 8850 5320
rect 9100 5310 9150 5320
rect 9350 5310 9400 5320
rect 9450 5310 9500 5320
rect 9600 5310 9650 5320
rect 550 5300 600 5310
rect 2000 5300 2050 5310
rect 2450 5300 2550 5310
rect 2600 5300 2750 5310
rect 3500 5300 3550 5310
rect 5700 5300 5850 5310
rect 6500 5300 6750 5310
rect 7350 5300 7400 5310
rect 7500 5300 7600 5310
rect 7900 5300 8050 5310
rect 8800 5300 8850 5310
rect 9100 5300 9150 5310
rect 9350 5300 9400 5310
rect 9450 5300 9500 5310
rect 9600 5300 9650 5310
rect 600 5290 650 5300
rect 2000 5290 2050 5300
rect 2400 5290 2450 5300
rect 2600 5290 2650 5300
rect 2750 5290 2900 5300
rect 5150 5290 5200 5300
rect 6250 5290 6450 5300
rect 7300 5290 7350 5300
rect 7900 5290 7950 5300
rect 8500 5290 8550 5300
rect 8650 5290 8700 5300
rect 8950 5290 9050 5300
rect 9600 5290 9650 5300
rect 9750 5290 9850 5300
rect 9900 5290 9950 5300
rect 600 5280 650 5290
rect 2000 5280 2050 5290
rect 2400 5280 2450 5290
rect 2600 5280 2650 5290
rect 2750 5280 2900 5290
rect 5150 5280 5200 5290
rect 6250 5280 6450 5290
rect 7300 5280 7350 5290
rect 7900 5280 7950 5290
rect 8500 5280 8550 5290
rect 8650 5280 8700 5290
rect 8950 5280 9050 5290
rect 9600 5280 9650 5290
rect 9750 5280 9850 5290
rect 9900 5280 9950 5290
rect 600 5270 650 5280
rect 2000 5270 2050 5280
rect 2400 5270 2450 5280
rect 2600 5270 2650 5280
rect 2750 5270 2900 5280
rect 5150 5270 5200 5280
rect 6250 5270 6450 5280
rect 7300 5270 7350 5280
rect 7900 5270 7950 5280
rect 8500 5270 8550 5280
rect 8650 5270 8700 5280
rect 8950 5270 9050 5280
rect 9600 5270 9650 5280
rect 9750 5270 9850 5280
rect 9900 5270 9950 5280
rect 600 5260 650 5270
rect 2000 5260 2050 5270
rect 2400 5260 2450 5270
rect 2600 5260 2650 5270
rect 2750 5260 2900 5270
rect 5150 5260 5200 5270
rect 6250 5260 6450 5270
rect 7300 5260 7350 5270
rect 7900 5260 7950 5270
rect 8500 5260 8550 5270
rect 8650 5260 8700 5270
rect 8950 5260 9050 5270
rect 9600 5260 9650 5270
rect 9750 5260 9850 5270
rect 9900 5260 9950 5270
rect 600 5250 650 5260
rect 2000 5250 2050 5260
rect 2400 5250 2450 5260
rect 2600 5250 2650 5260
rect 2750 5250 2900 5260
rect 5150 5250 5200 5260
rect 6250 5250 6450 5260
rect 7300 5250 7350 5260
rect 7900 5250 7950 5260
rect 8500 5250 8550 5260
rect 8650 5250 8700 5260
rect 8950 5250 9050 5260
rect 9600 5250 9650 5260
rect 9750 5250 9850 5260
rect 9900 5250 9950 5260
rect 600 5240 650 5250
rect 2000 5240 2050 5250
rect 3450 5240 3500 5250
rect 5100 5240 5150 5250
rect 7300 5240 7350 5250
rect 7900 5240 7950 5250
rect 8400 5240 8500 5250
rect 8750 5240 8850 5250
rect 9000 5240 9050 5250
rect 9250 5240 9300 5250
rect 9400 5240 9500 5250
rect 600 5230 650 5240
rect 2000 5230 2050 5240
rect 3450 5230 3500 5240
rect 5100 5230 5150 5240
rect 7300 5230 7350 5240
rect 7900 5230 7950 5240
rect 8400 5230 8500 5240
rect 8750 5230 8850 5240
rect 9000 5230 9050 5240
rect 9250 5230 9300 5240
rect 9400 5230 9500 5240
rect 600 5220 650 5230
rect 2000 5220 2050 5230
rect 3450 5220 3500 5230
rect 5100 5220 5150 5230
rect 7300 5220 7350 5230
rect 7900 5220 7950 5230
rect 8400 5220 8500 5230
rect 8750 5220 8850 5230
rect 9000 5220 9050 5230
rect 9250 5220 9300 5230
rect 9400 5220 9500 5230
rect 600 5210 650 5220
rect 2000 5210 2050 5220
rect 3450 5210 3500 5220
rect 5100 5210 5150 5220
rect 7300 5210 7350 5220
rect 7900 5210 7950 5220
rect 8400 5210 8500 5220
rect 8750 5210 8850 5220
rect 9000 5210 9050 5220
rect 9250 5210 9300 5220
rect 9400 5210 9500 5220
rect 600 5200 650 5210
rect 2000 5200 2050 5210
rect 3450 5200 3500 5210
rect 5100 5200 5150 5210
rect 7300 5200 7350 5210
rect 7900 5200 7950 5210
rect 8400 5200 8500 5210
rect 8750 5200 8850 5210
rect 9000 5200 9050 5210
rect 9250 5200 9300 5210
rect 9400 5200 9500 5210
rect 600 5190 700 5200
rect 2000 5190 2050 5200
rect 2700 5190 2800 5200
rect 2900 5190 3000 5200
rect 5100 5190 5200 5200
rect 7950 5190 8000 5200
rect 8250 5190 8300 5200
rect 9350 5190 9500 5200
rect 9600 5190 9650 5200
rect 9750 5190 9800 5200
rect 600 5180 700 5190
rect 2000 5180 2050 5190
rect 2700 5180 2800 5190
rect 2900 5180 3000 5190
rect 5100 5180 5200 5190
rect 7950 5180 8000 5190
rect 8250 5180 8300 5190
rect 9350 5180 9500 5190
rect 9600 5180 9650 5190
rect 9750 5180 9800 5190
rect 600 5170 700 5180
rect 2000 5170 2050 5180
rect 2700 5170 2800 5180
rect 2900 5170 3000 5180
rect 5100 5170 5200 5180
rect 7950 5170 8000 5180
rect 8250 5170 8300 5180
rect 9350 5170 9500 5180
rect 9600 5170 9650 5180
rect 9750 5170 9800 5180
rect 600 5160 700 5170
rect 2000 5160 2050 5170
rect 2700 5160 2800 5170
rect 2900 5160 3000 5170
rect 5100 5160 5200 5170
rect 7950 5160 8000 5170
rect 8250 5160 8300 5170
rect 9350 5160 9500 5170
rect 9600 5160 9650 5170
rect 9750 5160 9800 5170
rect 600 5150 700 5160
rect 2000 5150 2050 5160
rect 2700 5150 2800 5160
rect 2900 5150 3000 5160
rect 5100 5150 5200 5160
rect 7950 5150 8000 5160
rect 8250 5150 8300 5160
rect 9350 5150 9500 5160
rect 9600 5150 9650 5160
rect 9750 5150 9800 5160
rect 2050 5140 2100 5150
rect 2750 5140 3000 5150
rect 3400 5140 3450 5150
rect 5150 5140 5200 5150
rect 7950 5140 8050 5150
rect 8100 5140 8200 5150
rect 8400 5140 8450 5150
rect 8500 5140 8550 5150
rect 8600 5140 8650 5150
rect 8700 5140 8750 5150
rect 9050 5140 9100 5150
rect 9450 5140 9500 5150
rect 9850 5140 9950 5150
rect 2050 5130 2100 5140
rect 2750 5130 3000 5140
rect 3400 5130 3450 5140
rect 5150 5130 5200 5140
rect 7950 5130 8050 5140
rect 8100 5130 8200 5140
rect 8400 5130 8450 5140
rect 8500 5130 8550 5140
rect 8600 5130 8650 5140
rect 8700 5130 8750 5140
rect 9050 5130 9100 5140
rect 9450 5130 9500 5140
rect 9850 5130 9950 5140
rect 2050 5120 2100 5130
rect 2750 5120 3000 5130
rect 3400 5120 3450 5130
rect 5150 5120 5200 5130
rect 7950 5120 8050 5130
rect 8100 5120 8200 5130
rect 8400 5120 8450 5130
rect 8500 5120 8550 5130
rect 8600 5120 8650 5130
rect 8700 5120 8750 5130
rect 9050 5120 9100 5130
rect 9450 5120 9500 5130
rect 9850 5120 9950 5130
rect 2050 5110 2100 5120
rect 2750 5110 3000 5120
rect 3400 5110 3450 5120
rect 5150 5110 5200 5120
rect 7950 5110 8050 5120
rect 8100 5110 8200 5120
rect 8400 5110 8450 5120
rect 8500 5110 8550 5120
rect 8600 5110 8650 5120
rect 8700 5110 8750 5120
rect 9050 5110 9100 5120
rect 9450 5110 9500 5120
rect 9850 5110 9950 5120
rect 2050 5100 2100 5110
rect 2750 5100 3000 5110
rect 3400 5100 3450 5110
rect 5150 5100 5200 5110
rect 7950 5100 8050 5110
rect 8100 5100 8200 5110
rect 8400 5100 8450 5110
rect 8500 5100 8550 5110
rect 8600 5100 8650 5110
rect 8700 5100 8750 5110
rect 9050 5100 9100 5110
rect 9450 5100 9500 5110
rect 9850 5100 9950 5110
rect 500 5090 600 5100
rect 2050 5090 2150 5100
rect 2800 5090 2850 5100
rect 7300 5090 7350 5100
rect 7950 5090 8050 5100
rect 8150 5090 8300 5100
rect 8500 5090 8550 5100
rect 8700 5090 8900 5100
rect 9050 5090 9100 5100
rect 9200 5090 9250 5100
rect 9750 5090 9850 5100
rect 500 5080 600 5090
rect 2050 5080 2150 5090
rect 2800 5080 2850 5090
rect 7300 5080 7350 5090
rect 7950 5080 8050 5090
rect 8150 5080 8300 5090
rect 8500 5080 8550 5090
rect 8700 5080 8900 5090
rect 9050 5080 9100 5090
rect 9200 5080 9250 5090
rect 9750 5080 9850 5090
rect 500 5070 600 5080
rect 2050 5070 2150 5080
rect 2800 5070 2850 5080
rect 7300 5070 7350 5080
rect 7950 5070 8050 5080
rect 8150 5070 8300 5080
rect 8500 5070 8550 5080
rect 8700 5070 8900 5080
rect 9050 5070 9100 5080
rect 9200 5070 9250 5080
rect 9750 5070 9850 5080
rect 500 5060 600 5070
rect 2050 5060 2150 5070
rect 2800 5060 2850 5070
rect 7300 5060 7350 5070
rect 7950 5060 8050 5070
rect 8150 5060 8300 5070
rect 8500 5060 8550 5070
rect 8700 5060 8900 5070
rect 9050 5060 9100 5070
rect 9200 5060 9250 5070
rect 9750 5060 9850 5070
rect 500 5050 600 5060
rect 2050 5050 2150 5060
rect 2800 5050 2850 5060
rect 7300 5050 7350 5060
rect 7950 5050 8050 5060
rect 8150 5050 8300 5060
rect 8500 5050 8550 5060
rect 8700 5050 8900 5060
rect 9050 5050 9100 5060
rect 9200 5050 9250 5060
rect 9750 5050 9850 5060
rect 400 5040 450 5050
rect 2100 5040 2200 5050
rect 2750 5040 2900 5050
rect 3350 5040 3400 5050
rect 7950 5040 8000 5050
rect 8050 5040 8100 5050
rect 8650 5040 8700 5050
rect 8850 5040 8950 5050
rect 9350 5040 9400 5050
rect 9500 5040 9550 5050
rect 9600 5040 9650 5050
rect 400 5030 450 5040
rect 2100 5030 2200 5040
rect 2750 5030 2900 5040
rect 3350 5030 3400 5040
rect 7950 5030 8000 5040
rect 8050 5030 8100 5040
rect 8650 5030 8700 5040
rect 8850 5030 8950 5040
rect 9350 5030 9400 5040
rect 9500 5030 9550 5040
rect 9600 5030 9650 5040
rect 400 5020 450 5030
rect 2100 5020 2200 5030
rect 2750 5020 2900 5030
rect 3350 5020 3400 5030
rect 7950 5020 8000 5030
rect 8050 5020 8100 5030
rect 8650 5020 8700 5030
rect 8850 5020 8950 5030
rect 9350 5020 9400 5030
rect 9500 5020 9550 5030
rect 9600 5020 9650 5030
rect 400 5010 450 5020
rect 2100 5010 2200 5020
rect 2750 5010 2900 5020
rect 3350 5010 3400 5020
rect 7950 5010 8000 5020
rect 8050 5010 8100 5020
rect 8650 5010 8700 5020
rect 8850 5010 8950 5020
rect 9350 5010 9400 5020
rect 9500 5010 9550 5020
rect 9600 5010 9650 5020
rect 400 5000 450 5010
rect 2100 5000 2200 5010
rect 2750 5000 2900 5010
rect 3350 5000 3400 5010
rect 7950 5000 8000 5010
rect 8050 5000 8100 5010
rect 8650 5000 8700 5010
rect 8850 5000 8950 5010
rect 9350 5000 9400 5010
rect 9500 5000 9550 5010
rect 9600 5000 9650 5010
rect 400 4990 450 5000
rect 2100 4990 2300 5000
rect 2600 4990 2800 5000
rect 5700 4990 5750 5000
rect 7950 4990 8000 5000
rect 8400 4990 8450 5000
rect 8500 4990 8550 5000
rect 8650 4990 8750 5000
rect 9100 4990 9150 5000
rect 9200 4990 9350 5000
rect 9400 4990 9500 5000
rect 9600 4990 9650 5000
rect 9700 4990 9750 5000
rect 400 4980 450 4990
rect 2100 4980 2300 4990
rect 2600 4980 2800 4990
rect 5700 4980 5750 4990
rect 7950 4980 8000 4990
rect 8400 4980 8450 4990
rect 8500 4980 8550 4990
rect 8650 4980 8750 4990
rect 9100 4980 9150 4990
rect 9200 4980 9350 4990
rect 9400 4980 9500 4990
rect 9600 4980 9650 4990
rect 9700 4980 9750 4990
rect 400 4970 450 4980
rect 2100 4970 2300 4980
rect 2600 4970 2800 4980
rect 5700 4970 5750 4980
rect 7950 4970 8000 4980
rect 8400 4970 8450 4980
rect 8500 4970 8550 4980
rect 8650 4970 8750 4980
rect 9100 4970 9150 4980
rect 9200 4970 9350 4980
rect 9400 4970 9500 4980
rect 9600 4970 9650 4980
rect 9700 4970 9750 4980
rect 400 4960 450 4970
rect 2100 4960 2300 4970
rect 2600 4960 2800 4970
rect 5700 4960 5750 4970
rect 7950 4960 8000 4970
rect 8400 4960 8450 4970
rect 8500 4960 8550 4970
rect 8650 4960 8750 4970
rect 9100 4960 9150 4970
rect 9200 4960 9350 4970
rect 9400 4960 9500 4970
rect 9600 4960 9650 4970
rect 9700 4960 9750 4970
rect 400 4950 450 4960
rect 2100 4950 2300 4960
rect 2600 4950 2800 4960
rect 5700 4950 5750 4960
rect 7950 4950 8000 4960
rect 8400 4950 8450 4960
rect 8500 4950 8550 4960
rect 8650 4950 8750 4960
rect 9100 4950 9150 4960
rect 9200 4950 9350 4960
rect 9400 4950 9500 4960
rect 9600 4950 9650 4960
rect 9700 4950 9750 4960
rect 200 4940 450 4950
rect 2200 4940 2350 4950
rect 2600 4940 2700 4950
rect 3300 4940 3350 4950
rect 4000 4940 4050 4950
rect 4350 4940 4450 4950
rect 5600 4940 5700 4950
rect 5850 4940 5900 4950
rect 6300 4940 6450 4950
rect 7700 4940 7750 4950
rect 7950 4940 8000 4950
rect 8300 4940 8350 4950
rect 8450 4940 8500 4950
rect 8550 4940 8600 4950
rect 8700 4940 8750 4950
rect 9300 4940 9350 4950
rect 9450 4940 9500 4950
rect 9700 4940 9750 4950
rect 200 4930 450 4940
rect 2200 4930 2350 4940
rect 2600 4930 2700 4940
rect 3300 4930 3350 4940
rect 4000 4930 4050 4940
rect 4350 4930 4450 4940
rect 5600 4930 5700 4940
rect 5850 4930 5900 4940
rect 6300 4930 6450 4940
rect 7700 4930 7750 4940
rect 7950 4930 8000 4940
rect 8300 4930 8350 4940
rect 8450 4930 8500 4940
rect 8550 4930 8600 4940
rect 8700 4930 8750 4940
rect 9300 4930 9350 4940
rect 9450 4930 9500 4940
rect 9700 4930 9750 4940
rect 200 4920 450 4930
rect 2200 4920 2350 4930
rect 2600 4920 2700 4930
rect 3300 4920 3350 4930
rect 4000 4920 4050 4930
rect 4350 4920 4450 4930
rect 5600 4920 5700 4930
rect 5850 4920 5900 4930
rect 6300 4920 6450 4930
rect 7700 4920 7750 4930
rect 7950 4920 8000 4930
rect 8300 4920 8350 4930
rect 8450 4920 8500 4930
rect 8550 4920 8600 4930
rect 8700 4920 8750 4930
rect 9300 4920 9350 4930
rect 9450 4920 9500 4930
rect 9700 4920 9750 4930
rect 200 4910 450 4920
rect 2200 4910 2350 4920
rect 2600 4910 2700 4920
rect 3300 4910 3350 4920
rect 4000 4910 4050 4920
rect 4350 4910 4450 4920
rect 5600 4910 5700 4920
rect 5850 4910 5900 4920
rect 6300 4910 6450 4920
rect 7700 4910 7750 4920
rect 7950 4910 8000 4920
rect 8300 4910 8350 4920
rect 8450 4910 8500 4920
rect 8550 4910 8600 4920
rect 8700 4910 8750 4920
rect 9300 4910 9350 4920
rect 9450 4910 9500 4920
rect 9700 4910 9750 4920
rect 200 4900 450 4910
rect 2200 4900 2350 4910
rect 2600 4900 2700 4910
rect 3300 4900 3350 4910
rect 4000 4900 4050 4910
rect 4350 4900 4450 4910
rect 5600 4900 5700 4910
rect 5850 4900 5900 4910
rect 6300 4900 6450 4910
rect 7700 4900 7750 4910
rect 7950 4900 8000 4910
rect 8300 4900 8350 4910
rect 8450 4900 8500 4910
rect 8550 4900 8600 4910
rect 8700 4900 8750 4910
rect 9300 4900 9350 4910
rect 9450 4900 9500 4910
rect 9700 4900 9750 4910
rect 50 4890 150 4900
rect 2650 4890 2700 4900
rect 3300 4890 3350 4900
rect 3900 4890 4000 4900
rect 4050 4890 4100 4900
rect 4550 4890 4600 4900
rect 4700 4890 4800 4900
rect 5550 4890 5600 4900
rect 5650 4890 5700 4900
rect 5850 4890 6150 4900
rect 6400 4890 6450 4900
rect 7650 4890 7700 4900
rect 7950 4890 8000 4900
rect 8100 4890 8150 4900
rect 8200 4890 8400 4900
rect 8700 4890 8750 4900
rect 8850 4890 8900 4900
rect 8950 4890 9050 4900
rect 9700 4890 9750 4900
rect 50 4880 150 4890
rect 2650 4880 2700 4890
rect 3300 4880 3350 4890
rect 3900 4880 4000 4890
rect 4050 4880 4100 4890
rect 4550 4880 4600 4890
rect 4700 4880 4800 4890
rect 5550 4880 5600 4890
rect 5650 4880 5700 4890
rect 5850 4880 6150 4890
rect 6400 4880 6450 4890
rect 7650 4880 7700 4890
rect 7950 4880 8000 4890
rect 8100 4880 8150 4890
rect 8200 4880 8400 4890
rect 8700 4880 8750 4890
rect 8850 4880 8900 4890
rect 8950 4880 9050 4890
rect 9700 4880 9750 4890
rect 50 4870 150 4880
rect 2650 4870 2700 4880
rect 3300 4870 3350 4880
rect 3900 4870 4000 4880
rect 4050 4870 4100 4880
rect 4550 4870 4600 4880
rect 4700 4870 4800 4880
rect 5550 4870 5600 4880
rect 5650 4870 5700 4880
rect 5850 4870 6150 4880
rect 6400 4870 6450 4880
rect 7650 4870 7700 4880
rect 7950 4870 8000 4880
rect 8100 4870 8150 4880
rect 8200 4870 8400 4880
rect 8700 4870 8750 4880
rect 8850 4870 8900 4880
rect 8950 4870 9050 4880
rect 9700 4870 9750 4880
rect 50 4860 150 4870
rect 2650 4860 2700 4870
rect 3300 4860 3350 4870
rect 3900 4860 4000 4870
rect 4050 4860 4100 4870
rect 4550 4860 4600 4870
rect 4700 4860 4800 4870
rect 5550 4860 5600 4870
rect 5650 4860 5700 4870
rect 5850 4860 6150 4870
rect 6400 4860 6450 4870
rect 7650 4860 7700 4870
rect 7950 4860 8000 4870
rect 8100 4860 8150 4870
rect 8200 4860 8400 4870
rect 8700 4860 8750 4870
rect 8850 4860 8900 4870
rect 8950 4860 9050 4870
rect 9700 4860 9750 4870
rect 50 4850 150 4860
rect 2650 4850 2700 4860
rect 3300 4850 3350 4860
rect 3900 4850 4000 4860
rect 4050 4850 4100 4860
rect 4550 4850 4600 4860
rect 4700 4850 4800 4860
rect 5550 4850 5600 4860
rect 5650 4850 5700 4860
rect 5850 4850 6150 4860
rect 6400 4850 6450 4860
rect 7650 4850 7700 4860
rect 7950 4850 8000 4860
rect 8100 4850 8150 4860
rect 8200 4850 8400 4860
rect 8700 4850 8750 4860
rect 8850 4850 8900 4860
rect 8950 4850 9050 4860
rect 9700 4850 9750 4860
rect 0 4840 250 4850
rect 2700 4840 2750 4850
rect 3650 4840 3850 4850
rect 3950 4840 4000 4850
rect 4900 4840 4950 4850
rect 5500 4840 5550 4850
rect 5650 4840 5700 4850
rect 5950 4840 6000 4850
rect 6300 4840 6400 4850
rect 6450 4840 6500 4850
rect 7350 4840 7400 4850
rect 7950 4840 8200 4850
rect 8350 4840 8400 4850
rect 8750 4840 8800 4850
rect 9000 4840 9050 4850
rect 9350 4840 9400 4850
rect 0 4830 250 4840
rect 2700 4830 2750 4840
rect 3650 4830 3850 4840
rect 3950 4830 4000 4840
rect 4900 4830 4950 4840
rect 5500 4830 5550 4840
rect 5650 4830 5700 4840
rect 5950 4830 6000 4840
rect 6300 4830 6400 4840
rect 6450 4830 6500 4840
rect 7350 4830 7400 4840
rect 7950 4830 8200 4840
rect 8350 4830 8400 4840
rect 8750 4830 8800 4840
rect 9000 4830 9050 4840
rect 9350 4830 9400 4840
rect 0 4820 250 4830
rect 2700 4820 2750 4830
rect 3650 4820 3850 4830
rect 3950 4820 4000 4830
rect 4900 4820 4950 4830
rect 5500 4820 5550 4830
rect 5650 4820 5700 4830
rect 5950 4820 6000 4830
rect 6300 4820 6400 4830
rect 6450 4820 6500 4830
rect 7350 4820 7400 4830
rect 7950 4820 8200 4830
rect 8350 4820 8400 4830
rect 8750 4820 8800 4830
rect 9000 4820 9050 4830
rect 9350 4820 9400 4830
rect 0 4810 250 4820
rect 2700 4810 2750 4820
rect 3650 4810 3850 4820
rect 3950 4810 4000 4820
rect 4900 4810 4950 4820
rect 5500 4810 5550 4820
rect 5650 4810 5700 4820
rect 5950 4810 6000 4820
rect 6300 4810 6400 4820
rect 6450 4810 6500 4820
rect 7350 4810 7400 4820
rect 7950 4810 8200 4820
rect 8350 4810 8400 4820
rect 8750 4810 8800 4820
rect 9000 4810 9050 4820
rect 9350 4810 9400 4820
rect 0 4800 250 4810
rect 2700 4800 2750 4810
rect 3650 4800 3850 4810
rect 3950 4800 4000 4810
rect 4900 4800 4950 4810
rect 5500 4800 5550 4810
rect 5650 4800 5700 4810
rect 5950 4800 6000 4810
rect 6300 4800 6400 4810
rect 6450 4800 6500 4810
rect 7350 4800 7400 4810
rect 7950 4800 8200 4810
rect 8350 4800 8400 4810
rect 8750 4800 8800 4810
rect 9000 4800 9050 4810
rect 9350 4800 9400 4810
rect 0 4790 200 4800
rect 2400 4790 2450 4800
rect 2750 4790 2850 4800
rect 3250 4790 3350 4800
rect 3600 4790 3650 4800
rect 5000 4790 5050 4800
rect 5450 4790 5500 4800
rect 5600 4790 5650 4800
rect 6000 4790 6450 4800
rect 6500 4790 6550 4800
rect 7350 4790 7400 4800
rect 7700 4790 7800 4800
rect 7850 4790 8000 4800
rect 8450 4790 8500 4800
rect 8650 4790 8700 4800
rect 8800 4790 8900 4800
rect 9350 4790 9400 4800
rect 9500 4790 9600 4800
rect 9900 4790 9990 4800
rect 0 4780 200 4790
rect 2400 4780 2450 4790
rect 2750 4780 2850 4790
rect 3250 4780 3350 4790
rect 3600 4780 3650 4790
rect 5000 4780 5050 4790
rect 5450 4780 5500 4790
rect 5600 4780 5650 4790
rect 6000 4780 6450 4790
rect 6500 4780 6550 4790
rect 7350 4780 7400 4790
rect 7700 4780 7800 4790
rect 7850 4780 8000 4790
rect 8450 4780 8500 4790
rect 8650 4780 8700 4790
rect 8800 4780 8900 4790
rect 9350 4780 9400 4790
rect 9500 4780 9600 4790
rect 9900 4780 9990 4790
rect 0 4770 200 4780
rect 2400 4770 2450 4780
rect 2750 4770 2850 4780
rect 3250 4770 3350 4780
rect 3600 4770 3650 4780
rect 5000 4770 5050 4780
rect 5450 4770 5500 4780
rect 5600 4770 5650 4780
rect 6000 4770 6450 4780
rect 6500 4770 6550 4780
rect 7350 4770 7400 4780
rect 7700 4770 7800 4780
rect 7850 4770 8000 4780
rect 8450 4770 8500 4780
rect 8650 4770 8700 4780
rect 8800 4770 8900 4780
rect 9350 4770 9400 4780
rect 9500 4770 9600 4780
rect 9900 4770 9990 4780
rect 0 4760 200 4770
rect 2400 4760 2450 4770
rect 2750 4760 2850 4770
rect 3250 4760 3350 4770
rect 3600 4760 3650 4770
rect 5000 4760 5050 4770
rect 5450 4760 5500 4770
rect 5600 4760 5650 4770
rect 6000 4760 6450 4770
rect 6500 4760 6550 4770
rect 7350 4760 7400 4770
rect 7700 4760 7800 4770
rect 7850 4760 8000 4770
rect 8450 4760 8500 4770
rect 8650 4760 8700 4770
rect 8800 4760 8900 4770
rect 9350 4760 9400 4770
rect 9500 4760 9600 4770
rect 9900 4760 9990 4770
rect 0 4750 200 4760
rect 2400 4750 2450 4760
rect 2750 4750 2850 4760
rect 3250 4750 3350 4760
rect 3600 4750 3650 4760
rect 5000 4750 5050 4760
rect 5450 4750 5500 4760
rect 5600 4750 5650 4760
rect 6000 4750 6450 4760
rect 6500 4750 6550 4760
rect 7350 4750 7400 4760
rect 7700 4750 7800 4760
rect 7850 4750 8000 4760
rect 8450 4750 8500 4760
rect 8650 4750 8700 4760
rect 8800 4750 8900 4760
rect 9350 4750 9400 4760
rect 9500 4750 9600 4760
rect 9900 4750 9990 4760
rect 50 4740 200 4750
rect 2450 4740 2500 4750
rect 2750 4740 2900 4750
rect 2950 4740 3000 4750
rect 3300 4740 3350 4750
rect 3550 4740 3600 4750
rect 5050 4740 5100 4750
rect 5450 4740 5500 4750
rect 5600 4740 5650 4750
rect 6350 4740 6450 4750
rect 6550 4740 6600 4750
rect 7700 4740 7750 4750
rect 7800 4740 7850 4750
rect 8600 4740 8700 4750
rect 8750 4740 8800 4750
rect 9800 4740 9850 4750
rect 50 4730 200 4740
rect 2450 4730 2500 4740
rect 2750 4730 2900 4740
rect 2950 4730 3000 4740
rect 3300 4730 3350 4740
rect 3550 4730 3600 4740
rect 5050 4730 5100 4740
rect 5450 4730 5500 4740
rect 5600 4730 5650 4740
rect 6350 4730 6450 4740
rect 6550 4730 6600 4740
rect 7700 4730 7750 4740
rect 7800 4730 7850 4740
rect 8600 4730 8700 4740
rect 8750 4730 8800 4740
rect 9800 4730 9850 4740
rect 50 4720 200 4730
rect 2450 4720 2500 4730
rect 2750 4720 2900 4730
rect 2950 4720 3000 4730
rect 3300 4720 3350 4730
rect 3550 4720 3600 4730
rect 5050 4720 5100 4730
rect 5450 4720 5500 4730
rect 5600 4720 5650 4730
rect 6350 4720 6450 4730
rect 6550 4720 6600 4730
rect 7700 4720 7750 4730
rect 7800 4720 7850 4730
rect 8600 4720 8700 4730
rect 8750 4720 8800 4730
rect 9800 4720 9850 4730
rect 50 4710 200 4720
rect 2450 4710 2500 4720
rect 2750 4710 2900 4720
rect 2950 4710 3000 4720
rect 3300 4710 3350 4720
rect 3550 4710 3600 4720
rect 5050 4710 5100 4720
rect 5450 4710 5500 4720
rect 5600 4710 5650 4720
rect 6350 4710 6450 4720
rect 6550 4710 6600 4720
rect 7700 4710 7750 4720
rect 7800 4710 7850 4720
rect 8600 4710 8700 4720
rect 8750 4710 8800 4720
rect 9800 4710 9850 4720
rect 50 4700 200 4710
rect 2450 4700 2500 4710
rect 2750 4700 2900 4710
rect 2950 4700 3000 4710
rect 3300 4700 3350 4710
rect 3550 4700 3600 4710
rect 5050 4700 5100 4710
rect 5450 4700 5500 4710
rect 5600 4700 5650 4710
rect 6350 4700 6450 4710
rect 6550 4700 6600 4710
rect 7700 4700 7750 4710
rect 7800 4700 7850 4710
rect 8600 4700 8700 4710
rect 8750 4700 8800 4710
rect 9800 4700 9850 4710
rect 0 4690 150 4700
rect 2550 4690 2750 4700
rect 2800 4690 2850 4700
rect 2950 4690 3000 4700
rect 3150 4690 3200 4700
rect 3250 4690 3350 4700
rect 5100 4690 5150 4700
rect 5450 4690 5500 4700
rect 5600 4690 5700 4700
rect 6350 4690 6450 4700
rect 6550 4690 6600 4700
rect 7500 4690 7600 4700
rect 8200 4690 8350 4700
rect 8650 4690 8700 4700
rect 8750 4690 8800 4700
rect 9750 4690 9800 4700
rect 0 4680 150 4690
rect 2550 4680 2750 4690
rect 2800 4680 2850 4690
rect 2950 4680 3000 4690
rect 3150 4680 3200 4690
rect 3250 4680 3350 4690
rect 5100 4680 5150 4690
rect 5450 4680 5500 4690
rect 5600 4680 5700 4690
rect 6350 4680 6450 4690
rect 6550 4680 6600 4690
rect 7500 4680 7600 4690
rect 8200 4680 8350 4690
rect 8650 4680 8700 4690
rect 8750 4680 8800 4690
rect 9750 4680 9800 4690
rect 0 4670 150 4680
rect 2550 4670 2750 4680
rect 2800 4670 2850 4680
rect 2950 4670 3000 4680
rect 3150 4670 3200 4680
rect 3250 4670 3350 4680
rect 5100 4670 5150 4680
rect 5450 4670 5500 4680
rect 5600 4670 5700 4680
rect 6350 4670 6450 4680
rect 6550 4670 6600 4680
rect 7500 4670 7600 4680
rect 8200 4670 8350 4680
rect 8650 4670 8700 4680
rect 8750 4670 8800 4680
rect 9750 4670 9800 4680
rect 0 4660 150 4670
rect 2550 4660 2750 4670
rect 2800 4660 2850 4670
rect 2950 4660 3000 4670
rect 3150 4660 3200 4670
rect 3250 4660 3350 4670
rect 5100 4660 5150 4670
rect 5450 4660 5500 4670
rect 5600 4660 5700 4670
rect 6350 4660 6450 4670
rect 6550 4660 6600 4670
rect 7500 4660 7600 4670
rect 8200 4660 8350 4670
rect 8650 4660 8700 4670
rect 8750 4660 8800 4670
rect 9750 4660 9800 4670
rect 0 4650 150 4660
rect 2550 4650 2750 4660
rect 2800 4650 2850 4660
rect 2950 4650 3000 4660
rect 3150 4650 3200 4660
rect 3250 4650 3350 4660
rect 5100 4650 5150 4660
rect 5450 4650 5500 4660
rect 5600 4650 5700 4660
rect 6350 4650 6450 4660
rect 6550 4650 6600 4660
rect 7500 4650 7600 4660
rect 8200 4650 8350 4660
rect 8650 4650 8700 4660
rect 8750 4650 8800 4660
rect 9750 4650 9800 4660
rect 0 4640 50 4650
rect 3250 4640 3300 4650
rect 5150 4640 5200 4650
rect 5450 4640 5550 4650
rect 5750 4640 5950 4650
rect 6000 4640 6400 4650
rect 6550 4640 6600 4650
rect 7850 4640 7900 4650
rect 8000 4640 8050 4650
rect 8150 4640 8250 4650
rect 8450 4640 8500 4650
rect 8650 4640 8700 4650
rect 8900 4640 8950 4650
rect 9250 4640 9300 4650
rect 9700 4640 9750 4650
rect 0 4630 50 4640
rect 3250 4630 3300 4640
rect 5150 4630 5200 4640
rect 5450 4630 5550 4640
rect 5750 4630 5950 4640
rect 6000 4630 6400 4640
rect 6550 4630 6600 4640
rect 7850 4630 7900 4640
rect 8000 4630 8050 4640
rect 8150 4630 8250 4640
rect 8450 4630 8500 4640
rect 8650 4630 8700 4640
rect 8900 4630 8950 4640
rect 9250 4630 9300 4640
rect 9700 4630 9750 4640
rect 0 4620 50 4630
rect 3250 4620 3300 4630
rect 5150 4620 5200 4630
rect 5450 4620 5550 4630
rect 5750 4620 5950 4630
rect 6000 4620 6400 4630
rect 6550 4620 6600 4630
rect 7850 4620 7900 4630
rect 8000 4620 8050 4630
rect 8150 4620 8250 4630
rect 8450 4620 8500 4630
rect 8650 4620 8700 4630
rect 8900 4620 8950 4630
rect 9250 4620 9300 4630
rect 9700 4620 9750 4630
rect 0 4610 50 4620
rect 3250 4610 3300 4620
rect 5150 4610 5200 4620
rect 5450 4610 5550 4620
rect 5750 4610 5950 4620
rect 6000 4610 6400 4620
rect 6550 4610 6600 4620
rect 7850 4610 7900 4620
rect 8000 4610 8050 4620
rect 8150 4610 8250 4620
rect 8450 4610 8500 4620
rect 8650 4610 8700 4620
rect 8900 4610 8950 4620
rect 9250 4610 9300 4620
rect 9700 4610 9750 4620
rect 0 4600 50 4610
rect 3250 4600 3300 4610
rect 5150 4600 5200 4610
rect 5450 4600 5550 4610
rect 5750 4600 5950 4610
rect 6000 4600 6400 4610
rect 6550 4600 6600 4610
rect 7850 4600 7900 4610
rect 8000 4600 8050 4610
rect 8150 4600 8250 4610
rect 8450 4600 8500 4610
rect 8650 4600 8700 4610
rect 8900 4600 8950 4610
rect 9250 4600 9300 4610
rect 9700 4600 9750 4610
rect 3450 4590 3500 4600
rect 5500 4590 5600 4600
rect 5650 4590 5700 4600
rect 5750 4590 5800 4600
rect 6150 4590 6250 4600
rect 6500 4590 6550 4600
rect 7900 4590 7950 4600
rect 8000 4590 8100 4600
rect 8450 4590 8500 4600
rect 8650 4590 8700 4600
rect 9650 4590 9700 4600
rect 3450 4580 3500 4590
rect 5500 4580 5600 4590
rect 5650 4580 5700 4590
rect 5750 4580 5800 4590
rect 6150 4580 6250 4590
rect 6500 4580 6550 4590
rect 7900 4580 7950 4590
rect 8000 4580 8100 4590
rect 8450 4580 8500 4590
rect 8650 4580 8700 4590
rect 9650 4580 9700 4590
rect 3450 4570 3500 4580
rect 5500 4570 5600 4580
rect 5650 4570 5700 4580
rect 5750 4570 5800 4580
rect 6150 4570 6250 4580
rect 6500 4570 6550 4580
rect 7900 4570 7950 4580
rect 8000 4570 8100 4580
rect 8450 4570 8500 4580
rect 8650 4570 8700 4580
rect 9650 4570 9700 4580
rect 3450 4560 3500 4570
rect 5500 4560 5600 4570
rect 5650 4560 5700 4570
rect 5750 4560 5800 4570
rect 6150 4560 6250 4570
rect 6500 4560 6550 4570
rect 7900 4560 7950 4570
rect 8000 4560 8100 4570
rect 8450 4560 8500 4570
rect 8650 4560 8700 4570
rect 9650 4560 9700 4570
rect 3450 4550 3500 4560
rect 5500 4550 5600 4560
rect 5650 4550 5700 4560
rect 5750 4550 5800 4560
rect 6150 4550 6250 4560
rect 6500 4550 6550 4560
rect 7900 4550 7950 4560
rect 8000 4550 8100 4560
rect 8450 4550 8500 4560
rect 8650 4550 8700 4560
rect 9650 4550 9700 4560
rect 3000 4540 3050 4550
rect 3200 4540 3250 4550
rect 5500 4540 5600 4550
rect 6250 4540 6300 4550
rect 7400 4540 7500 4550
rect 7600 4540 7650 4550
rect 7700 4540 7900 4550
rect 8450 4540 8500 4550
rect 8550 4540 8600 4550
rect 8900 4540 8950 4550
rect 9600 4540 9650 4550
rect 3000 4530 3050 4540
rect 3200 4530 3250 4540
rect 5500 4530 5600 4540
rect 6250 4530 6300 4540
rect 7400 4530 7500 4540
rect 7600 4530 7650 4540
rect 7700 4530 7900 4540
rect 8450 4530 8500 4540
rect 8550 4530 8600 4540
rect 8900 4530 8950 4540
rect 9600 4530 9650 4540
rect 3000 4520 3050 4530
rect 3200 4520 3250 4530
rect 5500 4520 5600 4530
rect 6250 4520 6300 4530
rect 7400 4520 7500 4530
rect 7600 4520 7650 4530
rect 7700 4520 7900 4530
rect 8450 4520 8500 4530
rect 8550 4520 8600 4530
rect 8900 4520 8950 4530
rect 9600 4520 9650 4530
rect 3000 4510 3050 4520
rect 3200 4510 3250 4520
rect 5500 4510 5600 4520
rect 6250 4510 6300 4520
rect 7400 4510 7500 4520
rect 7600 4510 7650 4520
rect 7700 4510 7900 4520
rect 8450 4510 8500 4520
rect 8550 4510 8600 4520
rect 8900 4510 8950 4520
rect 9600 4510 9650 4520
rect 3000 4500 3050 4510
rect 3200 4500 3250 4510
rect 5500 4500 5600 4510
rect 6250 4500 6300 4510
rect 7400 4500 7500 4510
rect 7600 4500 7650 4510
rect 7700 4500 7900 4510
rect 8450 4500 8500 4510
rect 8550 4500 8600 4510
rect 8900 4500 8950 4510
rect 9600 4500 9650 4510
rect 2950 4490 3000 4500
rect 3050 4490 3150 4500
rect 3400 4490 3450 4500
rect 5250 4490 5300 4500
rect 5750 4490 5800 4500
rect 6200 4490 6250 4500
rect 6400 4490 6500 4500
rect 8350 4490 8400 4500
rect 9550 4490 9600 4500
rect 9950 4490 9990 4500
rect 2950 4480 3000 4490
rect 3050 4480 3150 4490
rect 3400 4480 3450 4490
rect 5250 4480 5300 4490
rect 5750 4480 5800 4490
rect 6200 4480 6250 4490
rect 6400 4480 6500 4490
rect 8350 4480 8400 4490
rect 9550 4480 9600 4490
rect 9950 4480 9990 4490
rect 2950 4470 3000 4480
rect 3050 4470 3150 4480
rect 3400 4470 3450 4480
rect 5250 4470 5300 4480
rect 5750 4470 5800 4480
rect 6200 4470 6250 4480
rect 6400 4470 6500 4480
rect 8350 4470 8400 4480
rect 9550 4470 9600 4480
rect 9950 4470 9990 4480
rect 2950 4460 3000 4470
rect 3050 4460 3150 4470
rect 3400 4460 3450 4470
rect 5250 4460 5300 4470
rect 5750 4460 5800 4470
rect 6200 4460 6250 4470
rect 6400 4460 6500 4470
rect 8350 4460 8400 4470
rect 9550 4460 9600 4470
rect 9950 4460 9990 4470
rect 2950 4450 3000 4460
rect 3050 4450 3150 4460
rect 3400 4450 3450 4460
rect 5250 4450 5300 4460
rect 5750 4450 5800 4460
rect 6200 4450 6250 4460
rect 6400 4450 6500 4460
rect 8350 4450 8400 4460
rect 9550 4450 9600 4460
rect 9950 4450 9990 4460
rect 2950 4440 3000 4450
rect 3050 4440 3150 4450
rect 3200 4440 3250 4450
rect 4600 4440 4700 4450
rect 6150 4440 6200 4450
rect 6350 4440 6500 4450
rect 7750 4440 7800 4450
rect 8150 4440 8250 4450
rect 9200 4440 9250 4450
rect 9500 4440 9550 4450
rect 9900 4440 9950 4450
rect 2950 4430 3000 4440
rect 3050 4430 3150 4440
rect 3200 4430 3250 4440
rect 4600 4430 4700 4440
rect 6150 4430 6200 4440
rect 6350 4430 6500 4440
rect 7750 4430 7800 4440
rect 8150 4430 8250 4440
rect 9200 4430 9250 4440
rect 9500 4430 9550 4440
rect 9900 4430 9950 4440
rect 2950 4420 3000 4430
rect 3050 4420 3150 4430
rect 3200 4420 3250 4430
rect 4600 4420 4700 4430
rect 6150 4420 6200 4430
rect 6350 4420 6500 4430
rect 7750 4420 7800 4430
rect 8150 4420 8250 4430
rect 9200 4420 9250 4430
rect 9500 4420 9550 4430
rect 9900 4420 9950 4430
rect 2950 4410 3000 4420
rect 3050 4410 3150 4420
rect 3200 4410 3250 4420
rect 4600 4410 4700 4420
rect 6150 4410 6200 4420
rect 6350 4410 6500 4420
rect 7750 4410 7800 4420
rect 8150 4410 8250 4420
rect 9200 4410 9250 4420
rect 9500 4410 9550 4420
rect 9900 4410 9950 4420
rect 2950 4400 3000 4410
rect 3050 4400 3150 4410
rect 3200 4400 3250 4410
rect 4600 4400 4700 4410
rect 6150 4400 6200 4410
rect 6350 4400 6500 4410
rect 7750 4400 7800 4410
rect 8150 4400 8250 4410
rect 9200 4400 9250 4410
rect 9500 4400 9550 4410
rect 9900 4400 9950 4410
rect 3050 4390 3100 4400
rect 3200 4390 3250 4400
rect 3350 4390 3400 4400
rect 4550 4390 4600 4400
rect 4750 4390 4850 4400
rect 6050 4390 6450 4400
rect 7850 4390 7900 4400
rect 8550 4390 8650 4400
rect 8700 4390 8750 4400
rect 9450 4390 9500 4400
rect 9850 4390 9990 4400
rect 3050 4380 3100 4390
rect 3200 4380 3250 4390
rect 3350 4380 3400 4390
rect 4550 4380 4600 4390
rect 4750 4380 4850 4390
rect 6050 4380 6450 4390
rect 7850 4380 7900 4390
rect 8550 4380 8650 4390
rect 8700 4380 8750 4390
rect 9450 4380 9500 4390
rect 9850 4380 9990 4390
rect 3050 4370 3100 4380
rect 3200 4370 3250 4380
rect 3350 4370 3400 4380
rect 4550 4370 4600 4380
rect 4750 4370 4850 4380
rect 6050 4370 6450 4380
rect 7850 4370 7900 4380
rect 8550 4370 8650 4380
rect 8700 4370 8750 4380
rect 9450 4370 9500 4380
rect 9850 4370 9990 4380
rect 3050 4360 3100 4370
rect 3200 4360 3250 4370
rect 3350 4360 3400 4370
rect 4550 4360 4600 4370
rect 4750 4360 4850 4370
rect 6050 4360 6450 4370
rect 7850 4360 7900 4370
rect 8550 4360 8650 4370
rect 8700 4360 8750 4370
rect 9450 4360 9500 4370
rect 9850 4360 9990 4370
rect 3050 4350 3100 4360
rect 3200 4350 3250 4360
rect 3350 4350 3400 4360
rect 4550 4350 4600 4360
rect 4750 4350 4850 4360
rect 6050 4350 6450 4360
rect 7850 4350 7900 4360
rect 8550 4350 8650 4360
rect 8700 4350 8750 4360
rect 9450 4350 9500 4360
rect 9850 4350 9990 4360
rect 2900 4340 2950 4350
rect 3150 4340 3300 4350
rect 4200 4340 4250 4350
rect 4900 4340 4950 4350
rect 5300 4340 5350 4350
rect 6200 4340 6300 4350
rect 7350 4340 7400 4350
rect 8400 4340 8450 4350
rect 9400 4340 9450 4350
rect 2900 4330 2950 4340
rect 3150 4330 3300 4340
rect 4200 4330 4250 4340
rect 4900 4330 4950 4340
rect 5300 4330 5350 4340
rect 6200 4330 6300 4340
rect 7350 4330 7400 4340
rect 8400 4330 8450 4340
rect 9400 4330 9450 4340
rect 2900 4320 2950 4330
rect 3150 4320 3300 4330
rect 4200 4320 4250 4330
rect 4900 4320 4950 4330
rect 5300 4320 5350 4330
rect 6200 4320 6300 4330
rect 7350 4320 7400 4330
rect 8400 4320 8450 4330
rect 9400 4320 9450 4330
rect 2900 4310 2950 4320
rect 3150 4310 3300 4320
rect 4200 4310 4250 4320
rect 4900 4310 4950 4320
rect 5300 4310 5350 4320
rect 6200 4310 6300 4320
rect 7350 4310 7400 4320
rect 8400 4310 8450 4320
rect 9400 4310 9450 4320
rect 2900 4300 2950 4310
rect 3150 4300 3300 4310
rect 4200 4300 4250 4310
rect 4900 4300 4950 4310
rect 5300 4300 5350 4310
rect 6200 4300 6300 4310
rect 7350 4300 7400 4310
rect 8400 4300 8450 4310
rect 9400 4300 9450 4310
rect 2900 4290 3200 4300
rect 4150 4290 4200 4300
rect 4300 4290 4350 4300
rect 4500 4290 4550 4300
rect 6100 4290 6200 4300
rect 7200 4290 7300 4300
rect 8400 4290 8450 4300
rect 8550 4290 8750 4300
rect 8800 4290 8850 4300
rect 2900 4280 3200 4290
rect 4150 4280 4200 4290
rect 4300 4280 4350 4290
rect 4500 4280 4550 4290
rect 6100 4280 6200 4290
rect 7200 4280 7300 4290
rect 8400 4280 8450 4290
rect 8550 4280 8750 4290
rect 8800 4280 8850 4290
rect 2900 4270 3200 4280
rect 4150 4270 4200 4280
rect 4300 4270 4350 4280
rect 4500 4270 4550 4280
rect 6100 4270 6200 4280
rect 7200 4270 7300 4280
rect 8400 4270 8450 4280
rect 8550 4270 8750 4280
rect 8800 4270 8850 4280
rect 2900 4260 3200 4270
rect 4150 4260 4200 4270
rect 4300 4260 4350 4270
rect 4500 4260 4550 4270
rect 6100 4260 6200 4270
rect 7200 4260 7300 4270
rect 8400 4260 8450 4270
rect 8550 4260 8750 4270
rect 8800 4260 8850 4270
rect 2900 4250 3200 4260
rect 4150 4250 4200 4260
rect 4300 4250 4350 4260
rect 4500 4250 4550 4260
rect 6100 4250 6200 4260
rect 7200 4250 7300 4260
rect 8400 4250 8450 4260
rect 8550 4250 8750 4260
rect 8800 4250 8850 4260
rect 2900 4240 2950 4250
rect 3000 4240 3200 4250
rect 4100 4240 4150 4250
rect 4350 4240 4400 4250
rect 4450 4240 4500 4250
rect 4950 4240 5000 4250
rect 7450 4240 7500 4250
rect 8450 4240 8500 4250
rect 9200 4240 9350 4250
rect 9750 4240 9800 4250
rect 2900 4230 2950 4240
rect 3000 4230 3200 4240
rect 4100 4230 4150 4240
rect 4350 4230 4400 4240
rect 4450 4230 4500 4240
rect 4950 4230 5000 4240
rect 7450 4230 7500 4240
rect 8450 4230 8500 4240
rect 9200 4230 9350 4240
rect 9750 4230 9800 4240
rect 2900 4220 2950 4230
rect 3000 4220 3200 4230
rect 4100 4220 4150 4230
rect 4350 4220 4400 4230
rect 4450 4220 4500 4230
rect 4950 4220 5000 4230
rect 7450 4220 7500 4230
rect 8450 4220 8500 4230
rect 9200 4220 9350 4230
rect 9750 4220 9800 4230
rect 2900 4210 2950 4220
rect 3000 4210 3200 4220
rect 4100 4210 4150 4220
rect 4350 4210 4400 4220
rect 4450 4210 4500 4220
rect 4950 4210 5000 4220
rect 7450 4210 7500 4220
rect 8450 4210 8500 4220
rect 9200 4210 9350 4220
rect 9750 4210 9800 4220
rect 2900 4200 2950 4210
rect 3000 4200 3200 4210
rect 4100 4200 4150 4210
rect 4350 4200 4400 4210
rect 4450 4200 4500 4210
rect 4950 4200 5000 4210
rect 7450 4200 7500 4210
rect 8450 4200 8500 4210
rect 9200 4200 9350 4210
rect 9750 4200 9800 4210
rect 2850 4190 2950 4200
rect 3000 4190 3250 4200
rect 5000 4190 5050 4200
rect 5500 4190 5600 4200
rect 7250 4190 7300 4200
rect 2850 4180 2950 4190
rect 3000 4180 3250 4190
rect 5000 4180 5050 4190
rect 5500 4180 5600 4190
rect 7250 4180 7300 4190
rect 2850 4170 2950 4180
rect 3000 4170 3250 4180
rect 5000 4170 5050 4180
rect 5500 4170 5600 4180
rect 7250 4170 7300 4180
rect 2850 4160 2950 4170
rect 3000 4160 3250 4170
rect 5000 4160 5050 4170
rect 5500 4160 5600 4170
rect 7250 4160 7300 4170
rect 2850 4150 2950 4160
rect 3000 4150 3250 4160
rect 5000 4150 5050 4160
rect 5500 4150 5600 4160
rect 7250 4150 7300 4160
rect 2850 4140 3200 4150
rect 4050 4140 4100 4150
rect 4650 4140 4900 4150
rect 5050 4140 5100 4150
rect 5400 4140 5450 4150
rect 5500 4140 5550 4150
rect 5600 4140 5650 4150
rect 7350 4140 7500 4150
rect 2850 4130 3200 4140
rect 4050 4130 4100 4140
rect 4650 4130 4900 4140
rect 5050 4130 5100 4140
rect 5400 4130 5450 4140
rect 5500 4130 5550 4140
rect 5600 4130 5650 4140
rect 7350 4130 7500 4140
rect 2850 4120 3200 4130
rect 4050 4120 4100 4130
rect 4650 4120 4900 4130
rect 5050 4120 5100 4130
rect 5400 4120 5450 4130
rect 5500 4120 5550 4130
rect 5600 4120 5650 4130
rect 7350 4120 7500 4130
rect 2850 4110 3200 4120
rect 4050 4110 4100 4120
rect 4650 4110 4900 4120
rect 5050 4110 5100 4120
rect 5400 4110 5450 4120
rect 5500 4110 5550 4120
rect 5600 4110 5650 4120
rect 7350 4110 7500 4120
rect 2850 4100 3200 4110
rect 4050 4100 4100 4110
rect 4650 4100 4900 4110
rect 5050 4100 5100 4110
rect 5400 4100 5450 4110
rect 5500 4100 5550 4110
rect 5600 4100 5650 4110
rect 7350 4100 7500 4110
rect 2850 4090 2900 4100
rect 2950 4090 3100 4100
rect 4600 4090 4650 4100
rect 5500 4090 5550 4100
rect 5650 4090 5700 4100
rect 7600 4090 7650 4100
rect 8750 4090 8800 4100
rect 2850 4080 2900 4090
rect 2950 4080 3100 4090
rect 4600 4080 4650 4090
rect 5500 4080 5550 4090
rect 5650 4080 5700 4090
rect 7600 4080 7650 4090
rect 8750 4080 8800 4090
rect 2850 4070 2900 4080
rect 2950 4070 3100 4080
rect 4600 4070 4650 4080
rect 5500 4070 5550 4080
rect 5650 4070 5700 4080
rect 7600 4070 7650 4080
rect 8750 4070 8800 4080
rect 2850 4060 2900 4070
rect 2950 4060 3100 4070
rect 4600 4060 4650 4070
rect 5500 4060 5550 4070
rect 5650 4060 5700 4070
rect 7600 4060 7650 4070
rect 8750 4060 8800 4070
rect 2850 4050 2900 4060
rect 2950 4050 3100 4060
rect 4600 4050 4650 4060
rect 5500 4050 5550 4060
rect 5650 4050 5700 4060
rect 7600 4050 7650 4060
rect 8750 4050 8800 4060
rect 2750 4040 2800 4050
rect 2950 4040 3100 4050
rect 4000 4040 4050 4050
rect 4600 4040 4650 4050
rect 4700 4040 4750 4050
rect 5100 4040 5150 4050
rect 5500 4040 5550 4050
rect 5700 4040 5750 4050
rect 7200 4040 7250 4050
rect 8350 4040 8550 4050
rect 8650 4040 8700 4050
rect 2750 4030 2800 4040
rect 2950 4030 3100 4040
rect 4000 4030 4050 4040
rect 4600 4030 4650 4040
rect 4700 4030 4750 4040
rect 5100 4030 5150 4040
rect 5500 4030 5550 4040
rect 5700 4030 5750 4040
rect 7200 4030 7250 4040
rect 8350 4030 8550 4040
rect 8650 4030 8700 4040
rect 2750 4020 2800 4030
rect 2950 4020 3100 4030
rect 4000 4020 4050 4030
rect 4600 4020 4650 4030
rect 4700 4020 4750 4030
rect 5100 4020 5150 4030
rect 5500 4020 5550 4030
rect 5700 4020 5750 4030
rect 7200 4020 7250 4030
rect 8350 4020 8550 4030
rect 8650 4020 8700 4030
rect 2750 4010 2800 4020
rect 2950 4010 3100 4020
rect 4000 4010 4050 4020
rect 4600 4010 4650 4020
rect 4700 4010 4750 4020
rect 5100 4010 5150 4020
rect 5500 4010 5550 4020
rect 5700 4010 5750 4020
rect 7200 4010 7250 4020
rect 8350 4010 8550 4020
rect 8650 4010 8700 4020
rect 2750 4000 2800 4010
rect 2950 4000 3100 4010
rect 4000 4000 4050 4010
rect 4600 4000 4650 4010
rect 4700 4000 4750 4010
rect 5100 4000 5150 4010
rect 5500 4000 5550 4010
rect 5700 4000 5750 4010
rect 7200 4000 7250 4010
rect 8350 4000 8550 4010
rect 8650 4000 8700 4010
rect 2900 3990 3000 4000
rect 3050 3990 3100 4000
rect 3250 3990 3300 4000
rect 3950 3990 4000 4000
rect 5150 3990 5200 4000
rect 5800 3990 6100 4000
rect 6150 3990 6350 4000
rect 7150 3990 7200 4000
rect 7850 3990 7900 4000
rect 8200 3990 8250 4000
rect 2900 3980 3000 3990
rect 3050 3980 3100 3990
rect 3250 3980 3300 3990
rect 3950 3980 4000 3990
rect 5150 3980 5200 3990
rect 5800 3980 6100 3990
rect 6150 3980 6350 3990
rect 7150 3980 7200 3990
rect 7850 3980 7900 3990
rect 8200 3980 8250 3990
rect 2900 3970 3000 3980
rect 3050 3970 3100 3980
rect 3250 3970 3300 3980
rect 3950 3970 4000 3980
rect 5150 3970 5200 3980
rect 5800 3970 6100 3980
rect 6150 3970 6350 3980
rect 7150 3970 7200 3980
rect 7850 3970 7900 3980
rect 8200 3970 8250 3980
rect 2900 3960 3000 3970
rect 3050 3960 3100 3970
rect 3250 3960 3300 3970
rect 3950 3960 4000 3970
rect 5150 3960 5200 3970
rect 5800 3960 6100 3970
rect 6150 3960 6350 3970
rect 7150 3960 7200 3970
rect 7850 3960 7900 3970
rect 8200 3960 8250 3970
rect 2900 3950 3000 3960
rect 3050 3950 3100 3960
rect 3250 3950 3300 3960
rect 3950 3950 4000 3960
rect 5150 3950 5200 3960
rect 5800 3950 6100 3960
rect 6150 3950 6350 3960
rect 7150 3950 7200 3960
rect 7850 3950 7900 3960
rect 8200 3950 8250 3960
rect 2850 3940 3150 3950
rect 3250 3940 3300 3950
rect 3900 3940 3950 3950
rect 4150 3940 4300 3950
rect 6300 3940 6350 3950
rect 7150 3940 7200 3950
rect 7950 3940 8000 3950
rect 8050 3940 8150 3950
rect 2850 3930 3150 3940
rect 3250 3930 3300 3940
rect 3900 3930 3950 3940
rect 4150 3930 4300 3940
rect 6300 3930 6350 3940
rect 7150 3930 7200 3940
rect 7950 3930 8000 3940
rect 8050 3930 8150 3940
rect 2850 3920 3150 3930
rect 3250 3920 3300 3930
rect 3900 3920 3950 3930
rect 4150 3920 4300 3930
rect 6300 3920 6350 3930
rect 7150 3920 7200 3930
rect 7950 3920 8000 3930
rect 8050 3920 8150 3930
rect 2850 3910 3150 3920
rect 3250 3910 3300 3920
rect 3900 3910 3950 3920
rect 4150 3910 4300 3920
rect 6300 3910 6350 3920
rect 7150 3910 7200 3920
rect 7950 3910 8000 3920
rect 8050 3910 8150 3920
rect 2850 3900 3150 3910
rect 3250 3900 3300 3910
rect 3900 3900 3950 3910
rect 4150 3900 4300 3910
rect 6300 3900 6350 3910
rect 7150 3900 7200 3910
rect 7950 3900 8000 3910
rect 8050 3900 8150 3910
rect 2850 3890 3100 3900
rect 3850 3890 3900 3900
rect 4100 3890 4150 3900
rect 4250 3890 4300 3900
rect 5200 3890 5250 3900
rect 6300 3890 6400 3900
rect 8050 3890 8100 3900
rect 9600 3890 9700 3900
rect 2850 3880 3100 3890
rect 3850 3880 3900 3890
rect 4100 3880 4150 3890
rect 4250 3880 4300 3890
rect 5200 3880 5250 3890
rect 6300 3880 6400 3890
rect 8050 3880 8100 3890
rect 9600 3880 9700 3890
rect 2850 3870 3100 3880
rect 3850 3870 3900 3880
rect 4100 3870 4150 3880
rect 4250 3870 4300 3880
rect 5200 3870 5250 3880
rect 6300 3870 6400 3880
rect 8050 3870 8100 3880
rect 9600 3870 9700 3880
rect 2850 3860 3100 3870
rect 3850 3860 3900 3870
rect 4100 3860 4150 3870
rect 4250 3860 4300 3870
rect 5200 3860 5250 3870
rect 6300 3860 6400 3870
rect 8050 3860 8100 3870
rect 9600 3860 9700 3870
rect 2850 3850 3100 3860
rect 3850 3850 3900 3860
rect 4100 3850 4150 3860
rect 4250 3850 4300 3860
rect 5200 3850 5250 3860
rect 6300 3850 6400 3860
rect 8050 3850 8100 3860
rect 9600 3850 9700 3860
rect 2850 3840 3000 3850
rect 3850 3840 3900 3850
rect 4050 3840 4100 3850
rect 4250 3840 4300 3850
rect 6300 3840 6400 3850
rect 7100 3840 7150 3850
rect 8200 3840 8250 3850
rect 9600 3840 9650 3850
rect 9700 3840 9750 3850
rect 2850 3830 3000 3840
rect 3850 3830 3900 3840
rect 4050 3830 4100 3840
rect 4250 3830 4300 3840
rect 6300 3830 6400 3840
rect 7100 3830 7150 3840
rect 8200 3830 8250 3840
rect 9600 3830 9650 3840
rect 9700 3830 9750 3840
rect 2850 3820 3000 3830
rect 3850 3820 3900 3830
rect 4050 3820 4100 3830
rect 4250 3820 4300 3830
rect 6300 3820 6400 3830
rect 7100 3820 7150 3830
rect 8200 3820 8250 3830
rect 9600 3820 9650 3830
rect 9700 3820 9750 3830
rect 2850 3810 3000 3820
rect 3850 3810 3900 3820
rect 4050 3810 4100 3820
rect 4250 3810 4300 3820
rect 6300 3810 6400 3820
rect 7100 3810 7150 3820
rect 8200 3810 8250 3820
rect 9600 3810 9650 3820
rect 9700 3810 9750 3820
rect 2850 3800 3000 3810
rect 3850 3800 3900 3810
rect 4050 3800 4100 3810
rect 4250 3800 4300 3810
rect 6300 3800 6400 3810
rect 7100 3800 7150 3810
rect 8200 3800 8250 3810
rect 9600 3800 9650 3810
rect 9700 3800 9750 3810
rect 2900 3790 2950 3800
rect 3100 3790 3200 3800
rect 3850 3790 3900 3800
rect 4000 3790 4050 3800
rect 4100 3790 4200 3800
rect 5250 3790 5300 3800
rect 6300 3790 6450 3800
rect 8100 3790 8250 3800
rect 9650 3790 9750 3800
rect 2900 3780 2950 3790
rect 3100 3780 3200 3790
rect 3850 3780 3900 3790
rect 4000 3780 4050 3790
rect 4100 3780 4200 3790
rect 5250 3780 5300 3790
rect 6300 3780 6450 3790
rect 8100 3780 8250 3790
rect 9650 3780 9750 3790
rect 2900 3770 2950 3780
rect 3100 3770 3200 3780
rect 3850 3770 3900 3780
rect 4000 3770 4050 3780
rect 4100 3770 4200 3780
rect 5250 3770 5300 3780
rect 6300 3770 6450 3780
rect 8100 3770 8250 3780
rect 9650 3770 9750 3780
rect 2900 3760 2950 3770
rect 3100 3760 3200 3770
rect 3850 3760 3900 3770
rect 4000 3760 4050 3770
rect 4100 3760 4200 3770
rect 5250 3760 5300 3770
rect 6300 3760 6450 3770
rect 8100 3760 8250 3770
rect 9650 3760 9750 3770
rect 2900 3750 2950 3760
rect 3100 3750 3200 3760
rect 3850 3750 3900 3760
rect 4000 3750 4050 3760
rect 4100 3750 4200 3760
rect 5250 3750 5300 3760
rect 6300 3750 6450 3760
rect 8100 3750 8250 3760
rect 9650 3750 9750 3760
rect 2850 3740 2950 3750
rect 3850 3740 3900 3750
rect 3950 3740 4050 3750
rect 6400 3740 6500 3750
rect 8150 3740 8200 3750
rect 2850 3730 2950 3740
rect 3850 3730 3900 3740
rect 3950 3730 4050 3740
rect 6400 3730 6500 3740
rect 8150 3730 8200 3740
rect 2850 3720 2950 3730
rect 3850 3720 3900 3730
rect 3950 3720 4050 3730
rect 6400 3720 6500 3730
rect 8150 3720 8200 3730
rect 2850 3710 2950 3720
rect 3850 3710 3900 3720
rect 3950 3710 4050 3720
rect 6400 3710 6500 3720
rect 8150 3710 8200 3720
rect 2850 3700 2950 3710
rect 3850 3700 3900 3710
rect 3950 3700 4050 3710
rect 6400 3700 6500 3710
rect 8150 3700 8200 3710
rect 3050 3690 3100 3700
rect 3300 3690 3350 3700
rect 3900 3690 4000 3700
rect 6450 3690 6500 3700
rect 7000 3690 7050 3700
rect 8400 3690 8500 3700
rect 3050 3680 3100 3690
rect 3300 3680 3350 3690
rect 3900 3680 4000 3690
rect 6450 3680 6500 3690
rect 7000 3680 7050 3690
rect 8400 3680 8500 3690
rect 3050 3670 3100 3680
rect 3300 3670 3350 3680
rect 3900 3670 4000 3680
rect 6450 3670 6500 3680
rect 7000 3670 7050 3680
rect 8400 3670 8500 3680
rect 3050 3660 3100 3670
rect 3300 3660 3350 3670
rect 3900 3660 4000 3670
rect 6450 3660 6500 3670
rect 7000 3660 7050 3670
rect 8400 3660 8500 3670
rect 3050 3650 3100 3660
rect 3300 3650 3350 3660
rect 3900 3650 4000 3660
rect 6450 3650 6500 3660
rect 7000 3650 7050 3660
rect 8400 3650 8500 3660
rect 3150 3640 3200 3650
rect 3300 3640 3350 3650
rect 3900 3640 3950 3650
rect 5300 3640 5350 3650
rect 6400 3640 6500 3650
rect 6950 3640 7000 3650
rect 8200 3640 8250 3650
rect 3150 3630 3200 3640
rect 3300 3630 3350 3640
rect 3900 3630 3950 3640
rect 5300 3630 5350 3640
rect 6400 3630 6500 3640
rect 6950 3630 7000 3640
rect 8200 3630 8250 3640
rect 3150 3620 3200 3630
rect 3300 3620 3350 3630
rect 3900 3620 3950 3630
rect 5300 3620 5350 3630
rect 6400 3620 6500 3630
rect 6950 3620 7000 3630
rect 8200 3620 8250 3630
rect 3150 3610 3200 3620
rect 3300 3610 3350 3620
rect 3900 3610 3950 3620
rect 5300 3610 5350 3620
rect 6400 3610 6500 3620
rect 6950 3610 7000 3620
rect 8200 3610 8250 3620
rect 3150 3600 3200 3610
rect 3300 3600 3350 3610
rect 3900 3600 3950 3610
rect 5300 3600 5350 3610
rect 6400 3600 6500 3610
rect 6950 3600 7000 3610
rect 8200 3600 8250 3610
rect 3350 3590 3400 3600
rect 3900 3590 3950 3600
rect 5300 3590 5350 3600
rect 6350 3590 6450 3600
rect 8250 3590 8300 3600
rect 8400 3590 8500 3600
rect 3350 3580 3400 3590
rect 3900 3580 3950 3590
rect 5300 3580 5350 3590
rect 6350 3580 6450 3590
rect 8250 3580 8300 3590
rect 8400 3580 8500 3590
rect 3350 3570 3400 3580
rect 3900 3570 3950 3580
rect 5300 3570 5350 3580
rect 6350 3570 6450 3580
rect 8250 3570 8300 3580
rect 8400 3570 8500 3580
rect 3350 3560 3400 3570
rect 3900 3560 3950 3570
rect 5300 3560 5350 3570
rect 6350 3560 6450 3570
rect 8250 3560 8300 3570
rect 8400 3560 8500 3570
rect 3350 3550 3400 3560
rect 3900 3550 3950 3560
rect 5300 3550 5350 3560
rect 6350 3550 6450 3560
rect 8250 3550 8300 3560
rect 8400 3550 8500 3560
rect 2500 3540 2600 3550
rect 3250 3540 3300 3550
rect 3400 3540 3450 3550
rect 3900 3540 3950 3550
rect 4700 3540 4750 3550
rect 5300 3540 5350 3550
rect 6350 3540 6400 3550
rect 8300 3540 8350 3550
rect 8450 3540 8500 3550
rect 9300 3540 9400 3550
rect 2500 3530 2600 3540
rect 3250 3530 3300 3540
rect 3400 3530 3450 3540
rect 3900 3530 3950 3540
rect 4700 3530 4750 3540
rect 5300 3530 5350 3540
rect 6350 3530 6400 3540
rect 8300 3530 8350 3540
rect 8450 3530 8500 3540
rect 9300 3530 9400 3540
rect 2500 3520 2600 3530
rect 3250 3520 3300 3530
rect 3400 3520 3450 3530
rect 3900 3520 3950 3530
rect 4700 3520 4750 3530
rect 5300 3520 5350 3530
rect 6350 3520 6400 3530
rect 8300 3520 8350 3530
rect 8450 3520 8500 3530
rect 9300 3520 9400 3530
rect 2500 3510 2600 3520
rect 3250 3510 3300 3520
rect 3400 3510 3450 3520
rect 3900 3510 3950 3520
rect 4700 3510 4750 3520
rect 5300 3510 5350 3520
rect 6350 3510 6400 3520
rect 8300 3510 8350 3520
rect 8450 3510 8500 3520
rect 9300 3510 9400 3520
rect 2500 3500 2600 3510
rect 3250 3500 3300 3510
rect 3400 3500 3450 3510
rect 3900 3500 3950 3510
rect 4700 3500 4750 3510
rect 5300 3500 5350 3510
rect 6350 3500 6400 3510
rect 8300 3500 8350 3510
rect 8450 3500 8500 3510
rect 9300 3500 9400 3510
rect 2300 3490 2350 3500
rect 2800 3490 2850 3500
rect 3400 3490 3450 3500
rect 4300 3490 4350 3500
rect 4500 3490 4700 3500
rect 4950 3490 5050 3500
rect 5300 3490 5350 3500
rect 6300 3490 6400 3500
rect 8450 3490 8500 3500
rect 9200 3490 9300 3500
rect 2300 3480 2350 3490
rect 2800 3480 2850 3490
rect 3400 3480 3450 3490
rect 4300 3480 4350 3490
rect 4500 3480 4700 3490
rect 4950 3480 5050 3490
rect 5300 3480 5350 3490
rect 6300 3480 6400 3490
rect 8450 3480 8500 3490
rect 9200 3480 9300 3490
rect 2300 3470 2350 3480
rect 2800 3470 2850 3480
rect 3400 3470 3450 3480
rect 4300 3470 4350 3480
rect 4500 3470 4700 3480
rect 4950 3470 5050 3480
rect 5300 3470 5350 3480
rect 6300 3470 6400 3480
rect 8450 3470 8500 3480
rect 9200 3470 9300 3480
rect 2300 3460 2350 3470
rect 2800 3460 2850 3470
rect 3400 3460 3450 3470
rect 4300 3460 4350 3470
rect 4500 3460 4700 3470
rect 4950 3460 5050 3470
rect 5300 3460 5350 3470
rect 6300 3460 6400 3470
rect 8450 3460 8500 3470
rect 9200 3460 9300 3470
rect 2300 3450 2350 3460
rect 2800 3450 2850 3460
rect 3400 3450 3450 3460
rect 4300 3450 4350 3460
rect 4500 3450 4700 3460
rect 4950 3450 5050 3460
rect 5300 3450 5350 3460
rect 6300 3450 6400 3460
rect 8450 3450 8500 3460
rect 9200 3450 9300 3460
rect 2200 3440 2250 3450
rect 2950 3440 3000 3450
rect 3950 3440 4000 3450
rect 4300 3440 4350 3450
rect 4450 3440 4500 3450
rect 4600 3440 4700 3450
rect 4900 3440 5000 3450
rect 5300 3440 5350 3450
rect 6200 3440 6350 3450
rect 9150 3440 9200 3450
rect 2200 3430 2250 3440
rect 2950 3430 3000 3440
rect 3950 3430 4000 3440
rect 4300 3430 4350 3440
rect 4450 3430 4500 3440
rect 4600 3430 4700 3440
rect 4900 3430 5000 3440
rect 5300 3430 5350 3440
rect 6200 3430 6350 3440
rect 9150 3430 9200 3440
rect 2200 3420 2250 3430
rect 2950 3420 3000 3430
rect 3950 3420 4000 3430
rect 4300 3420 4350 3430
rect 4450 3420 4500 3430
rect 4600 3420 4700 3430
rect 4900 3420 5000 3430
rect 5300 3420 5350 3430
rect 6200 3420 6350 3430
rect 9150 3420 9200 3430
rect 2200 3410 2250 3420
rect 2950 3410 3000 3420
rect 3950 3410 4000 3420
rect 4300 3410 4350 3420
rect 4450 3410 4500 3420
rect 4600 3410 4700 3420
rect 4900 3410 5000 3420
rect 5300 3410 5350 3420
rect 6200 3410 6350 3420
rect 9150 3410 9200 3420
rect 2200 3400 2250 3410
rect 2950 3400 3000 3410
rect 3950 3400 4000 3410
rect 4300 3400 4350 3410
rect 4450 3400 4500 3410
rect 4600 3400 4700 3410
rect 4900 3400 5000 3410
rect 5300 3400 5350 3410
rect 6200 3400 6350 3410
rect 9150 3400 9200 3410
rect 2150 3390 2200 3400
rect 3050 3390 3100 3400
rect 3500 3390 3600 3400
rect 3950 3390 4000 3400
rect 4250 3390 4350 3400
rect 4700 3390 4800 3400
rect 4850 3390 4900 3400
rect 5300 3390 5350 3400
rect 6150 3390 6250 3400
rect 9100 3390 9150 3400
rect 2150 3380 2200 3390
rect 3050 3380 3100 3390
rect 3500 3380 3600 3390
rect 3950 3380 4000 3390
rect 4250 3380 4350 3390
rect 4700 3380 4800 3390
rect 4850 3380 4900 3390
rect 5300 3380 5350 3390
rect 6150 3380 6250 3390
rect 9100 3380 9150 3390
rect 2150 3370 2200 3380
rect 3050 3370 3100 3380
rect 3500 3370 3600 3380
rect 3950 3370 4000 3380
rect 4250 3370 4350 3380
rect 4700 3370 4800 3380
rect 4850 3370 4900 3380
rect 5300 3370 5350 3380
rect 6150 3370 6250 3380
rect 9100 3370 9150 3380
rect 2150 3360 2200 3370
rect 3050 3360 3100 3370
rect 3500 3360 3600 3370
rect 3950 3360 4000 3370
rect 4250 3360 4350 3370
rect 4700 3360 4800 3370
rect 4850 3360 4900 3370
rect 5300 3360 5350 3370
rect 6150 3360 6250 3370
rect 9100 3360 9150 3370
rect 2150 3350 2200 3360
rect 3050 3350 3100 3360
rect 3500 3350 3600 3360
rect 3950 3350 4000 3360
rect 4250 3350 4350 3360
rect 4700 3350 4800 3360
rect 4850 3350 4900 3360
rect 5300 3350 5350 3360
rect 6150 3350 6250 3360
rect 9100 3350 9150 3360
rect 2100 3340 2150 3350
rect 3100 3340 3150 3350
rect 4000 3340 4050 3350
rect 4300 3340 4350 3350
rect 4600 3340 4700 3350
rect 4750 3340 4850 3350
rect 5300 3340 5350 3350
rect 6150 3340 6200 3350
rect 8450 3340 8500 3350
rect 9050 3340 9100 3350
rect 2100 3330 2150 3340
rect 3100 3330 3150 3340
rect 4000 3330 4050 3340
rect 4300 3330 4350 3340
rect 4600 3330 4700 3340
rect 4750 3330 4850 3340
rect 5300 3330 5350 3340
rect 6150 3330 6200 3340
rect 8450 3330 8500 3340
rect 9050 3330 9100 3340
rect 2100 3320 2150 3330
rect 3100 3320 3150 3330
rect 4000 3320 4050 3330
rect 4300 3320 4350 3330
rect 4600 3320 4700 3330
rect 4750 3320 4850 3330
rect 5300 3320 5350 3330
rect 6150 3320 6200 3330
rect 8450 3320 8500 3330
rect 9050 3320 9100 3330
rect 2100 3310 2150 3320
rect 3100 3310 3150 3320
rect 4000 3310 4050 3320
rect 4300 3310 4350 3320
rect 4600 3310 4700 3320
rect 4750 3310 4850 3320
rect 5300 3310 5350 3320
rect 6150 3310 6200 3320
rect 8450 3310 8500 3320
rect 9050 3310 9100 3320
rect 2100 3300 2150 3310
rect 3100 3300 3150 3310
rect 4000 3300 4050 3310
rect 4300 3300 4350 3310
rect 4600 3300 4700 3310
rect 4750 3300 4850 3310
rect 5300 3300 5350 3310
rect 6150 3300 6200 3310
rect 8450 3300 8500 3310
rect 9050 3300 9100 3310
rect 3550 3290 3600 3300
rect 4050 3290 4150 3300
rect 4200 3290 4250 3300
rect 4300 3290 4350 3300
rect 4500 3290 4550 3300
rect 4650 3290 4750 3300
rect 6150 3290 6200 3300
rect 9350 3290 9400 3300
rect 9650 3290 9700 3300
rect 3550 3280 3600 3290
rect 4050 3280 4150 3290
rect 4200 3280 4250 3290
rect 4300 3280 4350 3290
rect 4500 3280 4550 3290
rect 4650 3280 4750 3290
rect 6150 3280 6200 3290
rect 9350 3280 9400 3290
rect 9650 3280 9700 3290
rect 3550 3270 3600 3280
rect 4050 3270 4150 3280
rect 4200 3270 4250 3280
rect 4300 3270 4350 3280
rect 4500 3270 4550 3280
rect 4650 3270 4750 3280
rect 6150 3270 6200 3280
rect 9350 3270 9400 3280
rect 9650 3270 9700 3280
rect 3550 3260 3600 3270
rect 4050 3260 4150 3270
rect 4200 3260 4250 3270
rect 4300 3260 4350 3270
rect 4500 3260 4550 3270
rect 4650 3260 4750 3270
rect 6150 3260 6200 3270
rect 9350 3260 9400 3270
rect 9650 3260 9700 3270
rect 3550 3250 3600 3260
rect 4050 3250 4150 3260
rect 4200 3250 4250 3260
rect 4300 3250 4350 3260
rect 4500 3250 4550 3260
rect 4650 3250 4750 3260
rect 6150 3250 6200 3260
rect 9350 3250 9400 3260
rect 9650 3250 9700 3260
rect 2050 3240 2100 3250
rect 3150 3240 3200 3250
rect 3550 3240 3650 3250
rect 4100 3240 4350 3250
rect 4600 3240 4650 3250
rect 6200 3240 6250 3250
rect 6500 3240 6550 3250
rect 6600 3240 6650 3250
rect 8400 3240 8450 3250
rect 9100 3240 9150 3250
rect 9350 3240 9400 3250
rect 9550 3240 9600 3250
rect 2050 3230 2100 3240
rect 3150 3230 3200 3240
rect 3550 3230 3650 3240
rect 4100 3230 4350 3240
rect 4600 3230 4650 3240
rect 6200 3230 6250 3240
rect 6500 3230 6550 3240
rect 6600 3230 6650 3240
rect 8400 3230 8450 3240
rect 9100 3230 9150 3240
rect 9350 3230 9400 3240
rect 9550 3230 9600 3240
rect 2050 3220 2100 3230
rect 3150 3220 3200 3230
rect 3550 3220 3650 3230
rect 4100 3220 4350 3230
rect 4600 3220 4650 3230
rect 6200 3220 6250 3230
rect 6500 3220 6550 3230
rect 6600 3220 6650 3230
rect 8400 3220 8450 3230
rect 9100 3220 9150 3230
rect 9350 3220 9400 3230
rect 9550 3220 9600 3230
rect 2050 3210 2100 3220
rect 3150 3210 3200 3220
rect 3550 3210 3650 3220
rect 4100 3210 4350 3220
rect 4600 3210 4650 3220
rect 6200 3210 6250 3220
rect 6500 3210 6550 3220
rect 6600 3210 6650 3220
rect 8400 3210 8450 3220
rect 9100 3210 9150 3220
rect 9350 3210 9400 3220
rect 9550 3210 9600 3220
rect 2050 3200 2100 3210
rect 3150 3200 3200 3210
rect 3550 3200 3650 3210
rect 4100 3200 4350 3210
rect 4600 3200 4650 3210
rect 6200 3200 6250 3210
rect 6500 3200 6550 3210
rect 6600 3200 6650 3210
rect 8400 3200 8450 3210
rect 9100 3200 9150 3210
rect 9350 3200 9400 3210
rect 9550 3200 9600 3210
rect 4150 3190 4200 3200
rect 4300 3190 4400 3200
rect 4500 3190 4550 3200
rect 4900 3190 4950 3200
rect 5250 3190 5300 3200
rect 6200 3190 6300 3200
rect 6350 3190 6400 3200
rect 6600 3190 6650 3200
rect 9050 3190 9100 3200
rect 9200 3190 9400 3200
rect 9450 3190 9550 3200
rect 4150 3180 4200 3190
rect 4300 3180 4400 3190
rect 4500 3180 4550 3190
rect 4900 3180 4950 3190
rect 5250 3180 5300 3190
rect 6200 3180 6300 3190
rect 6350 3180 6400 3190
rect 6600 3180 6650 3190
rect 9050 3180 9100 3190
rect 9200 3180 9400 3190
rect 9450 3180 9550 3190
rect 4150 3170 4200 3180
rect 4300 3170 4400 3180
rect 4500 3170 4550 3180
rect 4900 3170 4950 3180
rect 5250 3170 5300 3180
rect 6200 3170 6300 3180
rect 6350 3170 6400 3180
rect 6600 3170 6650 3180
rect 9050 3170 9100 3180
rect 9200 3170 9400 3180
rect 9450 3170 9550 3180
rect 4150 3160 4200 3170
rect 4300 3160 4400 3170
rect 4500 3160 4550 3170
rect 4900 3160 4950 3170
rect 5250 3160 5300 3170
rect 6200 3160 6300 3170
rect 6350 3160 6400 3170
rect 6600 3160 6650 3170
rect 9050 3160 9100 3170
rect 9200 3160 9400 3170
rect 9450 3160 9550 3170
rect 4150 3150 4200 3160
rect 4300 3150 4400 3160
rect 4500 3150 4550 3160
rect 4900 3150 4950 3160
rect 5250 3150 5300 3160
rect 6200 3150 6300 3160
rect 6350 3150 6400 3160
rect 6600 3150 6650 3160
rect 9050 3150 9100 3160
rect 9200 3150 9400 3160
rect 9450 3150 9550 3160
rect 4150 3140 4200 3150
rect 4500 3140 4550 3150
rect 4850 3140 4900 3150
rect 5250 3140 5300 3150
rect 8350 3140 8400 3150
rect 9050 3140 9100 3150
rect 9200 3140 9550 3150
rect 4150 3130 4200 3140
rect 4500 3130 4550 3140
rect 4850 3130 4900 3140
rect 5250 3130 5300 3140
rect 8350 3130 8400 3140
rect 9050 3130 9100 3140
rect 9200 3130 9550 3140
rect 4150 3120 4200 3130
rect 4500 3120 4550 3130
rect 4850 3120 4900 3130
rect 5250 3120 5300 3130
rect 8350 3120 8400 3130
rect 9050 3120 9100 3130
rect 9200 3120 9550 3130
rect 4150 3110 4200 3120
rect 4500 3110 4550 3120
rect 4850 3110 4900 3120
rect 5250 3110 5300 3120
rect 8350 3110 8400 3120
rect 9050 3110 9100 3120
rect 9200 3110 9550 3120
rect 4150 3100 4200 3110
rect 4500 3100 4550 3110
rect 4850 3100 4900 3110
rect 5250 3100 5300 3110
rect 8350 3100 8400 3110
rect 9050 3100 9100 3110
rect 9200 3100 9550 3110
rect 2000 3090 2050 3100
rect 3800 3090 3900 3100
rect 4000 3090 4050 3100
rect 4150 3090 4250 3100
rect 4500 3090 4550 3100
rect 4600 3090 4800 3100
rect 4850 3090 4900 3100
rect 6550 3090 6600 3100
rect 9250 3090 9400 3100
rect 9450 3090 9500 3100
rect 2000 3080 2050 3090
rect 3800 3080 3900 3090
rect 4000 3080 4050 3090
rect 4150 3080 4250 3090
rect 4500 3080 4550 3090
rect 4600 3080 4800 3090
rect 4850 3080 4900 3090
rect 6550 3080 6600 3090
rect 9250 3080 9400 3090
rect 9450 3080 9500 3090
rect 2000 3070 2050 3080
rect 3800 3070 3900 3080
rect 4000 3070 4050 3080
rect 4150 3070 4250 3080
rect 4500 3070 4550 3080
rect 4600 3070 4800 3080
rect 4850 3070 4900 3080
rect 6550 3070 6600 3080
rect 9250 3070 9400 3080
rect 9450 3070 9500 3080
rect 2000 3060 2050 3070
rect 3800 3060 3900 3070
rect 4000 3060 4050 3070
rect 4150 3060 4250 3070
rect 4500 3060 4550 3070
rect 4600 3060 4800 3070
rect 4850 3060 4900 3070
rect 6550 3060 6600 3070
rect 9250 3060 9400 3070
rect 9450 3060 9500 3070
rect 2000 3050 2050 3060
rect 3800 3050 3900 3060
rect 4000 3050 4050 3060
rect 4150 3050 4250 3060
rect 4500 3050 4550 3060
rect 4600 3050 4800 3060
rect 4850 3050 4900 3060
rect 6550 3050 6600 3060
rect 9250 3050 9400 3060
rect 9450 3050 9500 3060
rect 2000 3040 2050 3050
rect 3150 3040 3200 3050
rect 3750 3040 3850 3050
rect 4200 3040 4300 3050
rect 4550 3040 4650 3050
rect 4750 3040 4850 3050
rect 5200 3040 5250 3050
rect 6550 3040 6600 3050
rect 8300 3040 8350 3050
rect 9000 3040 9050 3050
rect 9400 3040 9450 3050
rect 2000 3030 2050 3040
rect 3150 3030 3200 3040
rect 3750 3030 3850 3040
rect 4200 3030 4300 3040
rect 4550 3030 4650 3040
rect 4750 3030 4850 3040
rect 5200 3030 5250 3040
rect 6550 3030 6600 3040
rect 8300 3030 8350 3040
rect 9000 3030 9050 3040
rect 9400 3030 9450 3040
rect 2000 3020 2050 3030
rect 3150 3020 3200 3030
rect 3750 3020 3850 3030
rect 4200 3020 4300 3030
rect 4550 3020 4650 3030
rect 4750 3020 4850 3030
rect 5200 3020 5250 3030
rect 6550 3020 6600 3030
rect 8300 3020 8350 3030
rect 9000 3020 9050 3030
rect 9400 3020 9450 3030
rect 2000 3010 2050 3020
rect 3150 3010 3200 3020
rect 3750 3010 3850 3020
rect 4200 3010 4300 3020
rect 4550 3010 4650 3020
rect 4750 3010 4850 3020
rect 5200 3010 5250 3020
rect 6550 3010 6600 3020
rect 8300 3010 8350 3020
rect 9000 3010 9050 3020
rect 9400 3010 9450 3020
rect 2000 3000 2050 3010
rect 3150 3000 3200 3010
rect 3750 3000 3850 3010
rect 4200 3000 4300 3010
rect 4550 3000 4650 3010
rect 4750 3000 4850 3010
rect 5200 3000 5250 3010
rect 6550 3000 6600 3010
rect 8300 3000 8350 3010
rect 9000 3000 9050 3010
rect 9400 3000 9450 3010
rect 2000 2990 2050 3000
rect 3150 2990 3200 3000
rect 3850 2990 3900 3000
rect 4150 2990 4200 3000
rect 4300 2990 4350 3000
rect 4550 2990 4850 3000
rect 8950 2990 9050 3000
rect 9150 2990 9200 3000
rect 9250 2990 9400 3000
rect 2000 2980 2050 2990
rect 3150 2980 3200 2990
rect 3850 2980 3900 2990
rect 4150 2980 4200 2990
rect 4300 2980 4350 2990
rect 4550 2980 4850 2990
rect 8950 2980 9050 2990
rect 9150 2980 9200 2990
rect 9250 2980 9400 2990
rect 2000 2970 2050 2980
rect 3150 2970 3200 2980
rect 3850 2970 3900 2980
rect 4150 2970 4200 2980
rect 4300 2970 4350 2980
rect 4550 2970 4850 2980
rect 8950 2970 9050 2980
rect 9150 2970 9200 2980
rect 9250 2970 9400 2980
rect 2000 2960 2050 2970
rect 3150 2960 3200 2970
rect 3850 2960 3900 2970
rect 4150 2960 4200 2970
rect 4300 2960 4350 2970
rect 4550 2960 4850 2970
rect 8950 2960 9050 2970
rect 9150 2960 9200 2970
rect 9250 2960 9400 2970
rect 2000 2950 2050 2960
rect 3150 2950 3200 2960
rect 3850 2950 3900 2960
rect 4150 2950 4200 2960
rect 4300 2950 4350 2960
rect 4550 2950 4850 2960
rect 8950 2950 9050 2960
rect 9150 2950 9200 2960
rect 9250 2950 9400 2960
rect 3850 2940 3900 2950
rect 4350 2940 4400 2950
rect 4550 2940 4600 2950
rect 5150 2940 5200 2950
rect 8900 2940 9000 2950
rect 9100 2940 9150 2950
rect 9200 2940 9400 2950
rect 3850 2930 3900 2940
rect 4350 2930 4400 2940
rect 4550 2930 4600 2940
rect 5150 2930 5200 2940
rect 8900 2930 9000 2940
rect 9100 2930 9150 2940
rect 9200 2930 9400 2940
rect 3850 2920 3900 2930
rect 4350 2920 4400 2930
rect 4550 2920 4600 2930
rect 5150 2920 5200 2930
rect 8900 2920 9000 2930
rect 9100 2920 9150 2930
rect 9200 2920 9400 2930
rect 3850 2910 3900 2920
rect 4350 2910 4400 2920
rect 4550 2910 4600 2920
rect 5150 2910 5200 2920
rect 8900 2910 9000 2920
rect 9100 2910 9150 2920
rect 9200 2910 9400 2920
rect 3850 2900 3900 2910
rect 4350 2900 4400 2910
rect 4550 2900 4600 2910
rect 5150 2900 5200 2910
rect 8900 2900 9000 2910
rect 9100 2900 9150 2910
rect 9200 2900 9400 2910
rect 3950 2890 4000 2900
rect 4450 2890 4500 2900
rect 4600 2890 4750 2900
rect 5100 2890 5150 2900
rect 7250 2890 7300 2900
rect 7350 2890 7400 2900
rect 7500 2890 7550 2900
rect 8200 2890 8250 2900
rect 8900 2890 9100 2900
rect 9200 2890 9300 2900
rect 3950 2880 4000 2890
rect 4450 2880 4500 2890
rect 4600 2880 4750 2890
rect 5100 2880 5150 2890
rect 7250 2880 7300 2890
rect 7350 2880 7400 2890
rect 7500 2880 7550 2890
rect 8200 2880 8250 2890
rect 8900 2880 9100 2890
rect 9200 2880 9300 2890
rect 3950 2870 4000 2880
rect 4450 2870 4500 2880
rect 4600 2870 4750 2880
rect 5100 2870 5150 2880
rect 7250 2870 7300 2880
rect 7350 2870 7400 2880
rect 7500 2870 7550 2880
rect 8200 2870 8250 2880
rect 8900 2870 9100 2880
rect 9200 2870 9300 2880
rect 3950 2860 4000 2870
rect 4450 2860 4500 2870
rect 4600 2860 4750 2870
rect 5100 2860 5150 2870
rect 7250 2860 7300 2870
rect 7350 2860 7400 2870
rect 7500 2860 7550 2870
rect 8200 2860 8250 2870
rect 8900 2860 9100 2870
rect 9200 2860 9300 2870
rect 3950 2850 4000 2860
rect 4450 2850 4500 2860
rect 4600 2850 4750 2860
rect 5100 2850 5150 2860
rect 7250 2850 7300 2860
rect 7350 2850 7400 2860
rect 7500 2850 7550 2860
rect 8200 2850 8250 2860
rect 8900 2850 9100 2860
rect 9200 2850 9300 2860
rect 4250 2840 4300 2850
rect 4500 2840 4850 2850
rect 4900 2840 5100 2850
rect 7150 2840 7200 2850
rect 7550 2840 7600 2850
rect 8900 2840 9050 2850
rect 4250 2830 4300 2840
rect 4500 2830 4850 2840
rect 4900 2830 5100 2840
rect 7150 2830 7200 2840
rect 7550 2830 7600 2840
rect 8900 2830 9050 2840
rect 4250 2820 4300 2830
rect 4500 2820 4850 2830
rect 4900 2820 5100 2830
rect 7150 2820 7200 2830
rect 7550 2820 7600 2830
rect 8900 2820 9050 2830
rect 4250 2810 4300 2820
rect 4500 2810 4850 2820
rect 4900 2810 5100 2820
rect 7150 2810 7200 2820
rect 7550 2810 7600 2820
rect 8900 2810 9050 2820
rect 4250 2800 4300 2810
rect 4500 2800 4850 2810
rect 4900 2800 5100 2810
rect 7150 2800 7200 2810
rect 7550 2800 7600 2810
rect 8900 2800 9050 2810
rect 3900 2790 3950 2800
rect 4750 2790 5150 2800
rect 6000 2790 6100 2800
rect 7050 2790 7100 2800
rect 8750 2790 9000 2800
rect 3900 2780 3950 2790
rect 4750 2780 5150 2790
rect 6000 2780 6100 2790
rect 7050 2780 7100 2790
rect 8750 2780 9000 2790
rect 3900 2770 3950 2780
rect 4750 2770 5150 2780
rect 6000 2770 6100 2780
rect 7050 2770 7100 2780
rect 8750 2770 9000 2780
rect 3900 2760 3950 2770
rect 4750 2760 5150 2770
rect 6000 2760 6100 2770
rect 7050 2760 7100 2770
rect 8750 2760 9000 2770
rect 3900 2750 3950 2760
rect 4750 2750 5150 2760
rect 6000 2750 6100 2760
rect 7050 2750 7100 2760
rect 8750 2750 9000 2760
rect 5000 2740 5150 2750
rect 5900 2740 6150 2750
rect 6950 2740 7000 2750
rect 7650 2740 7700 2750
rect 8700 2740 8750 2750
rect 8800 2740 8950 2750
rect 9050 2740 9150 2750
rect 9950 2740 9990 2750
rect 5000 2730 5150 2740
rect 5900 2730 6150 2740
rect 6950 2730 7000 2740
rect 7650 2730 7700 2740
rect 8700 2730 8750 2740
rect 8800 2730 8950 2740
rect 9050 2730 9150 2740
rect 9950 2730 9990 2740
rect 5000 2720 5150 2730
rect 5900 2720 6150 2730
rect 6950 2720 7000 2730
rect 7650 2720 7700 2730
rect 8700 2720 8750 2730
rect 8800 2720 8950 2730
rect 9050 2720 9150 2730
rect 9950 2720 9990 2730
rect 5000 2710 5150 2720
rect 5900 2710 6150 2720
rect 6950 2710 7000 2720
rect 7650 2710 7700 2720
rect 8700 2710 8750 2720
rect 8800 2710 8950 2720
rect 9050 2710 9150 2720
rect 9950 2710 9990 2720
rect 5000 2700 5150 2710
rect 5900 2700 6150 2710
rect 6950 2700 7000 2710
rect 7650 2700 7700 2710
rect 8700 2700 8750 2710
rect 8800 2700 8950 2710
rect 9050 2700 9150 2710
rect 9950 2700 9990 2710
rect 1950 2690 2000 2700
rect 4950 2690 5100 2700
rect 5850 2690 6000 2700
rect 6100 2690 6200 2700
rect 6900 2690 6950 2700
rect 8900 2690 9200 2700
rect 9950 2690 9990 2700
rect 1950 2680 2000 2690
rect 4950 2680 5100 2690
rect 5850 2680 6000 2690
rect 6100 2680 6200 2690
rect 6900 2680 6950 2690
rect 8900 2680 9200 2690
rect 9950 2680 9990 2690
rect 1950 2670 2000 2680
rect 4950 2670 5100 2680
rect 5850 2670 6000 2680
rect 6100 2670 6200 2680
rect 6900 2670 6950 2680
rect 8900 2670 9200 2680
rect 9950 2670 9990 2680
rect 1950 2660 2000 2670
rect 4950 2660 5100 2670
rect 5850 2660 6000 2670
rect 6100 2660 6200 2670
rect 6900 2660 6950 2670
rect 8900 2660 9200 2670
rect 9950 2660 9990 2670
rect 1950 2650 2000 2660
rect 4950 2650 5100 2660
rect 5850 2650 6000 2660
rect 6100 2650 6200 2660
rect 6900 2650 6950 2660
rect 8900 2650 9200 2660
rect 9950 2650 9990 2660
rect 2100 2640 2250 2650
rect 2800 2640 2850 2650
rect 2900 2640 3000 2650
rect 3050 2640 3100 2650
rect 4950 2640 5050 2650
rect 5800 2640 5950 2650
rect 6150 2640 6250 2650
rect 6850 2640 6900 2650
rect 8000 2640 8050 2650
rect 9000 2640 9050 2650
rect 9150 2640 9200 2650
rect 9950 2640 9990 2650
rect 2100 2630 2250 2640
rect 2800 2630 2850 2640
rect 2900 2630 3000 2640
rect 3050 2630 3100 2640
rect 4950 2630 5050 2640
rect 5800 2630 5950 2640
rect 6150 2630 6250 2640
rect 6850 2630 6900 2640
rect 8000 2630 8050 2640
rect 9000 2630 9050 2640
rect 9150 2630 9200 2640
rect 9950 2630 9990 2640
rect 2100 2620 2250 2630
rect 2800 2620 2850 2630
rect 2900 2620 3000 2630
rect 3050 2620 3100 2630
rect 4950 2620 5050 2630
rect 5800 2620 5950 2630
rect 6150 2620 6250 2630
rect 6850 2620 6900 2630
rect 8000 2620 8050 2630
rect 9000 2620 9050 2630
rect 9150 2620 9200 2630
rect 9950 2620 9990 2630
rect 2100 2610 2250 2620
rect 2800 2610 2850 2620
rect 2900 2610 3000 2620
rect 3050 2610 3100 2620
rect 4950 2610 5050 2620
rect 5800 2610 5950 2620
rect 6150 2610 6250 2620
rect 6850 2610 6900 2620
rect 8000 2610 8050 2620
rect 9000 2610 9050 2620
rect 9150 2610 9200 2620
rect 9950 2610 9990 2620
rect 2100 2600 2250 2610
rect 2800 2600 2850 2610
rect 2900 2600 3000 2610
rect 3050 2600 3100 2610
rect 4950 2600 5050 2610
rect 5800 2600 5950 2610
rect 6150 2600 6250 2610
rect 6850 2600 6900 2610
rect 8000 2600 8050 2610
rect 9000 2600 9050 2610
rect 9150 2600 9200 2610
rect 9950 2600 9990 2610
rect 1900 2590 1950 2600
rect 4250 2590 4300 2600
rect 5750 2590 5950 2600
rect 6200 2590 6250 2600
rect 6800 2590 6850 2600
rect 7750 2590 7800 2600
rect 9000 2590 9050 2600
rect 9900 2590 9990 2600
rect 1900 2580 1950 2590
rect 4250 2580 4300 2590
rect 5750 2580 5950 2590
rect 6200 2580 6250 2590
rect 6800 2580 6850 2590
rect 7750 2580 7800 2590
rect 9000 2580 9050 2590
rect 9900 2580 9990 2590
rect 1900 2570 1950 2580
rect 4250 2570 4300 2580
rect 5750 2570 5950 2580
rect 6200 2570 6250 2580
rect 6800 2570 6850 2580
rect 7750 2570 7800 2580
rect 9000 2570 9050 2580
rect 9900 2570 9990 2580
rect 1900 2560 1950 2570
rect 4250 2560 4300 2570
rect 5750 2560 5950 2570
rect 6200 2560 6250 2570
rect 6800 2560 6850 2570
rect 7750 2560 7800 2570
rect 9000 2560 9050 2570
rect 9900 2560 9990 2570
rect 1900 2550 1950 2560
rect 4250 2550 4300 2560
rect 5750 2550 5950 2560
rect 6200 2550 6250 2560
rect 6800 2550 6850 2560
rect 7750 2550 7800 2560
rect 9000 2550 9050 2560
rect 9900 2550 9990 2560
rect 1900 2540 1950 2550
rect 2050 2540 2100 2550
rect 2200 2540 2350 2550
rect 4150 2540 4200 2550
rect 5750 2540 5850 2550
rect 6200 2540 6300 2550
rect 6750 2540 6800 2550
rect 7250 2540 7300 2550
rect 7850 2540 7900 2550
rect 9050 2540 9150 2550
rect 9450 2540 9550 2550
rect 1900 2530 1950 2540
rect 2050 2530 2100 2540
rect 2200 2530 2350 2540
rect 4150 2530 4200 2540
rect 5750 2530 5850 2540
rect 6200 2530 6300 2540
rect 6750 2530 6800 2540
rect 7250 2530 7300 2540
rect 7850 2530 7900 2540
rect 9050 2530 9150 2540
rect 9450 2530 9550 2540
rect 1900 2520 1950 2530
rect 2050 2520 2100 2530
rect 2200 2520 2350 2530
rect 4150 2520 4200 2530
rect 5750 2520 5850 2530
rect 6200 2520 6300 2530
rect 6750 2520 6800 2530
rect 7250 2520 7300 2530
rect 7850 2520 7900 2530
rect 9050 2520 9150 2530
rect 9450 2520 9550 2530
rect 1900 2510 1950 2520
rect 2050 2510 2100 2520
rect 2200 2510 2350 2520
rect 4150 2510 4200 2520
rect 5750 2510 5850 2520
rect 6200 2510 6300 2520
rect 6750 2510 6800 2520
rect 7250 2510 7300 2520
rect 7850 2510 7900 2520
rect 9050 2510 9150 2520
rect 9450 2510 9550 2520
rect 1900 2500 1950 2510
rect 2050 2500 2100 2510
rect 2200 2500 2350 2510
rect 4150 2500 4200 2510
rect 5750 2500 5850 2510
rect 6200 2500 6300 2510
rect 6750 2500 6800 2510
rect 7250 2500 7300 2510
rect 7850 2500 7900 2510
rect 9050 2500 9150 2510
rect 9450 2500 9550 2510
rect 1900 2490 1950 2500
rect 4000 2490 4050 2500
rect 5550 2490 5800 2500
rect 6250 2490 6350 2500
rect 7300 2490 7350 2500
rect 9300 2490 9400 2500
rect 9450 2490 9650 2500
rect 1900 2480 1950 2490
rect 4000 2480 4050 2490
rect 5550 2480 5800 2490
rect 6250 2480 6350 2490
rect 7300 2480 7350 2490
rect 9300 2480 9400 2490
rect 9450 2480 9650 2490
rect 1900 2470 1950 2480
rect 4000 2470 4050 2480
rect 5550 2470 5800 2480
rect 6250 2470 6350 2480
rect 7300 2470 7350 2480
rect 9300 2470 9400 2480
rect 9450 2470 9650 2480
rect 1900 2460 1950 2470
rect 4000 2460 4050 2470
rect 5550 2460 5800 2470
rect 6250 2460 6350 2470
rect 7300 2460 7350 2470
rect 9300 2460 9400 2470
rect 9450 2460 9650 2470
rect 1900 2450 1950 2460
rect 4000 2450 4050 2460
rect 5550 2450 5800 2460
rect 6250 2450 6350 2460
rect 7300 2450 7350 2460
rect 9300 2450 9400 2460
rect 9450 2450 9650 2460
rect 5550 2440 5800 2450
rect 6300 2440 6350 2450
rect 9350 2440 9500 2450
rect 9550 2440 9700 2450
rect 5550 2430 5800 2440
rect 6300 2430 6350 2440
rect 9350 2430 9500 2440
rect 9550 2430 9700 2440
rect 5550 2420 5800 2430
rect 6300 2420 6350 2430
rect 9350 2420 9500 2430
rect 9550 2420 9700 2430
rect 5550 2410 5800 2420
rect 6300 2410 6350 2420
rect 9350 2410 9500 2420
rect 9550 2410 9700 2420
rect 5550 2400 5800 2410
rect 6300 2400 6350 2410
rect 9350 2400 9500 2410
rect 9550 2400 9700 2410
rect 3250 2390 3300 2400
rect 5650 2390 5750 2400
rect 6300 2390 6400 2400
rect 6750 2390 6850 2400
rect 9400 2390 9450 2400
rect 9600 2390 9800 2400
rect 3250 2380 3300 2390
rect 5650 2380 5750 2390
rect 6300 2380 6400 2390
rect 6750 2380 6850 2390
rect 9400 2380 9450 2390
rect 9600 2380 9800 2390
rect 3250 2370 3300 2380
rect 5650 2370 5750 2380
rect 6300 2370 6400 2380
rect 6750 2370 6850 2380
rect 9400 2370 9450 2380
rect 9600 2370 9800 2380
rect 3250 2360 3300 2370
rect 5650 2360 5750 2370
rect 6300 2360 6400 2370
rect 6750 2360 6850 2370
rect 9400 2360 9450 2370
rect 9600 2360 9800 2370
rect 3250 2350 3300 2360
rect 5650 2350 5750 2360
rect 6300 2350 6400 2360
rect 6750 2350 6850 2360
rect 9400 2350 9450 2360
rect 9600 2350 9800 2360
rect 1850 2340 1900 2350
rect 5650 2340 5750 2350
rect 5900 2340 6000 2350
rect 6350 2340 6400 2350
rect 6750 2340 6950 2350
rect 8400 2340 8550 2350
rect 9150 2340 9450 2350
rect 9600 2340 9650 2350
rect 9750 2340 9800 2350
rect 1850 2330 1900 2340
rect 5650 2330 5750 2340
rect 5900 2330 6000 2340
rect 6350 2330 6400 2340
rect 6750 2330 6950 2340
rect 8400 2330 8550 2340
rect 9150 2330 9450 2340
rect 9600 2330 9650 2340
rect 9750 2330 9800 2340
rect 1850 2320 1900 2330
rect 5650 2320 5750 2330
rect 5900 2320 6000 2330
rect 6350 2320 6400 2330
rect 6750 2320 6950 2330
rect 8400 2320 8550 2330
rect 9150 2320 9450 2330
rect 9600 2320 9650 2330
rect 9750 2320 9800 2330
rect 1850 2310 1900 2320
rect 5650 2310 5750 2320
rect 5900 2310 6000 2320
rect 6350 2310 6400 2320
rect 6750 2310 6950 2320
rect 8400 2310 8550 2320
rect 9150 2310 9450 2320
rect 9600 2310 9650 2320
rect 9750 2310 9800 2320
rect 1850 2300 1900 2310
rect 5650 2300 5750 2310
rect 5900 2300 6000 2310
rect 6350 2300 6400 2310
rect 6750 2300 6950 2310
rect 8400 2300 8550 2310
rect 9150 2300 9450 2310
rect 9600 2300 9650 2310
rect 9750 2300 9800 2310
rect 5400 2290 5550 2300
rect 5600 2290 5700 2300
rect 5900 2290 6050 2300
rect 6400 2290 6450 2300
rect 6800 2290 6850 2300
rect 6950 2290 7200 2300
rect 7500 2290 7600 2300
rect 8550 2290 8600 2300
rect 9250 2290 9350 2300
rect 9450 2290 9500 2300
rect 9550 2290 9600 2300
rect 9750 2290 9800 2300
rect 5400 2280 5550 2290
rect 5600 2280 5700 2290
rect 5900 2280 6050 2290
rect 6400 2280 6450 2290
rect 6800 2280 6850 2290
rect 6950 2280 7200 2290
rect 7500 2280 7600 2290
rect 8550 2280 8600 2290
rect 9250 2280 9350 2290
rect 9450 2280 9500 2290
rect 9550 2280 9600 2290
rect 9750 2280 9800 2290
rect 5400 2270 5550 2280
rect 5600 2270 5700 2280
rect 5900 2270 6050 2280
rect 6400 2270 6450 2280
rect 6800 2270 6850 2280
rect 6950 2270 7200 2280
rect 7500 2270 7600 2280
rect 8550 2270 8600 2280
rect 9250 2270 9350 2280
rect 9450 2270 9500 2280
rect 9550 2270 9600 2280
rect 9750 2270 9800 2280
rect 5400 2260 5550 2270
rect 5600 2260 5700 2270
rect 5900 2260 6050 2270
rect 6400 2260 6450 2270
rect 6800 2260 6850 2270
rect 6950 2260 7200 2270
rect 7500 2260 7600 2270
rect 8550 2260 8600 2270
rect 9250 2260 9350 2270
rect 9450 2260 9500 2270
rect 9550 2260 9600 2270
rect 9750 2260 9800 2270
rect 5400 2250 5550 2260
rect 5600 2250 5700 2260
rect 5900 2250 6050 2260
rect 6400 2250 6450 2260
rect 6800 2250 6850 2260
rect 6950 2250 7200 2260
rect 7500 2250 7600 2260
rect 8550 2250 8600 2260
rect 9250 2250 9350 2260
rect 9450 2250 9500 2260
rect 9550 2250 9600 2260
rect 9750 2250 9800 2260
rect 5350 2240 5700 2250
rect 6450 2240 6500 2250
rect 6800 2240 6900 2250
rect 7250 2240 7350 2250
rect 7500 2240 7550 2250
rect 7600 2240 7650 2250
rect 8650 2240 8800 2250
rect 9050 2240 9100 2250
rect 9200 2240 9250 2250
rect 9400 2240 9450 2250
rect 9500 2240 9550 2250
rect 5350 2230 5700 2240
rect 6450 2230 6500 2240
rect 6800 2230 6900 2240
rect 7250 2230 7350 2240
rect 7500 2230 7550 2240
rect 7600 2230 7650 2240
rect 8650 2230 8800 2240
rect 9050 2230 9100 2240
rect 9200 2230 9250 2240
rect 9400 2230 9450 2240
rect 9500 2230 9550 2240
rect 5350 2220 5700 2230
rect 6450 2220 6500 2230
rect 6800 2220 6900 2230
rect 7250 2220 7350 2230
rect 7500 2220 7550 2230
rect 7600 2220 7650 2230
rect 8650 2220 8800 2230
rect 9050 2220 9100 2230
rect 9200 2220 9250 2230
rect 9400 2220 9450 2230
rect 9500 2220 9550 2230
rect 5350 2210 5700 2220
rect 6450 2210 6500 2220
rect 6800 2210 6900 2220
rect 7250 2210 7350 2220
rect 7500 2210 7550 2220
rect 7600 2210 7650 2220
rect 8650 2210 8800 2220
rect 9050 2210 9100 2220
rect 9200 2210 9250 2220
rect 9400 2210 9450 2220
rect 9500 2210 9550 2220
rect 5350 2200 5700 2210
rect 6450 2200 6500 2210
rect 6800 2200 6900 2210
rect 7250 2200 7350 2210
rect 7500 2200 7550 2210
rect 7600 2200 7650 2210
rect 8650 2200 8800 2210
rect 9050 2200 9100 2210
rect 9200 2200 9250 2210
rect 9400 2200 9450 2210
rect 9500 2200 9550 2210
rect 2650 2190 2750 2200
rect 5300 2190 5650 2200
rect 6900 2190 7000 2200
rect 7350 2190 7400 2200
rect 7650 2190 7700 2200
rect 9200 2190 9250 2200
rect 9500 2190 9600 2200
rect 9650 2190 9750 2200
rect 2650 2180 2750 2190
rect 5300 2180 5650 2190
rect 6900 2180 7000 2190
rect 7350 2180 7400 2190
rect 7650 2180 7700 2190
rect 9200 2180 9250 2190
rect 9500 2180 9600 2190
rect 9650 2180 9750 2190
rect 2650 2170 2750 2180
rect 5300 2170 5650 2180
rect 6900 2170 7000 2180
rect 7350 2170 7400 2180
rect 7650 2170 7700 2180
rect 9200 2170 9250 2180
rect 9500 2170 9600 2180
rect 9650 2170 9750 2180
rect 2650 2160 2750 2170
rect 5300 2160 5650 2170
rect 6900 2160 7000 2170
rect 7350 2160 7400 2170
rect 7650 2160 7700 2170
rect 9200 2160 9250 2170
rect 9500 2160 9600 2170
rect 9650 2160 9750 2170
rect 2650 2150 2750 2160
rect 5300 2150 5650 2160
rect 6900 2150 7000 2160
rect 7350 2150 7400 2160
rect 7650 2150 7700 2160
rect 9200 2150 9250 2160
rect 9500 2150 9600 2160
rect 9650 2150 9750 2160
rect 5250 2140 5550 2150
rect 6100 2140 6200 2150
rect 6950 2140 7050 2150
rect 7250 2140 7350 2150
rect 7750 2140 7800 2150
rect 9200 2140 9250 2150
rect 9650 2140 9700 2150
rect 5250 2130 5550 2140
rect 6100 2130 6200 2140
rect 6950 2130 7050 2140
rect 7250 2130 7350 2140
rect 7750 2130 7800 2140
rect 9200 2130 9250 2140
rect 9650 2130 9700 2140
rect 5250 2120 5550 2130
rect 6100 2120 6200 2130
rect 6950 2120 7050 2130
rect 7250 2120 7350 2130
rect 7750 2120 7800 2130
rect 9200 2120 9250 2130
rect 9650 2120 9700 2130
rect 5250 2110 5550 2120
rect 6100 2110 6200 2120
rect 6950 2110 7050 2120
rect 7250 2110 7350 2120
rect 7750 2110 7800 2120
rect 9200 2110 9250 2120
rect 9650 2110 9700 2120
rect 5250 2100 5550 2110
rect 6100 2100 6200 2110
rect 6950 2100 7050 2110
rect 7250 2100 7350 2110
rect 7750 2100 7800 2110
rect 9200 2100 9250 2110
rect 9650 2100 9700 2110
rect 5100 2090 5150 2100
rect 5250 2090 5350 2100
rect 6100 2090 6200 2100
rect 6500 2090 6550 2100
rect 6750 2090 6800 2100
rect 7000 2090 7350 2100
rect 8400 2090 8450 2100
rect 9150 2090 9200 2100
rect 9250 2090 9300 2100
rect 9600 2090 9650 2100
rect 5100 2080 5150 2090
rect 5250 2080 5350 2090
rect 6100 2080 6200 2090
rect 6500 2080 6550 2090
rect 6750 2080 6800 2090
rect 7000 2080 7350 2090
rect 8400 2080 8450 2090
rect 9150 2080 9200 2090
rect 9250 2080 9300 2090
rect 9600 2080 9650 2090
rect 5100 2070 5150 2080
rect 5250 2070 5350 2080
rect 6100 2070 6200 2080
rect 6500 2070 6550 2080
rect 6750 2070 6800 2080
rect 7000 2070 7350 2080
rect 8400 2070 8450 2080
rect 9150 2070 9200 2080
rect 9250 2070 9300 2080
rect 9600 2070 9650 2080
rect 5100 2060 5150 2070
rect 5250 2060 5350 2070
rect 6100 2060 6200 2070
rect 6500 2060 6550 2070
rect 6750 2060 6800 2070
rect 7000 2060 7350 2070
rect 8400 2060 8450 2070
rect 9150 2060 9200 2070
rect 9250 2060 9300 2070
rect 9600 2060 9650 2070
rect 5100 2050 5150 2060
rect 5250 2050 5350 2060
rect 6100 2050 6200 2060
rect 6500 2050 6550 2060
rect 6750 2050 6800 2060
rect 7000 2050 7350 2060
rect 8400 2050 8450 2060
rect 9150 2050 9200 2060
rect 9250 2050 9300 2060
rect 9600 2050 9650 2060
rect 3250 2040 3300 2050
rect 5100 2040 5300 2050
rect 6100 2040 6300 2050
rect 6500 2040 6550 2050
rect 6750 2040 6800 2050
rect 7050 2040 7250 2050
rect 7900 2040 7950 2050
rect 9050 2040 9100 2050
rect 3250 2030 3300 2040
rect 5100 2030 5300 2040
rect 6100 2030 6300 2040
rect 6500 2030 6550 2040
rect 6750 2030 6800 2040
rect 7050 2030 7250 2040
rect 7900 2030 7950 2040
rect 9050 2030 9100 2040
rect 3250 2020 3300 2030
rect 5100 2020 5300 2030
rect 6100 2020 6300 2030
rect 6500 2020 6550 2030
rect 6750 2020 6800 2030
rect 7050 2020 7250 2030
rect 7900 2020 7950 2030
rect 9050 2020 9100 2030
rect 3250 2010 3300 2020
rect 5100 2010 5300 2020
rect 6100 2010 6300 2020
rect 6500 2010 6550 2020
rect 6750 2010 6800 2020
rect 7050 2010 7250 2020
rect 7900 2010 7950 2020
rect 9050 2010 9100 2020
rect 3250 2000 3300 2010
rect 5100 2000 5300 2010
rect 6100 2000 6300 2010
rect 6500 2000 6550 2010
rect 6750 2000 6800 2010
rect 7050 2000 7250 2010
rect 7900 2000 7950 2010
rect 9050 2000 9100 2010
rect 3250 1990 3350 2000
rect 4800 1990 4850 2000
rect 5000 1990 5250 2000
rect 6100 1990 6350 2000
rect 6500 1990 6550 2000
rect 7750 1990 7950 2000
rect 8600 1990 9050 2000
rect 3250 1980 3350 1990
rect 4800 1980 4850 1990
rect 5000 1980 5250 1990
rect 6100 1980 6350 1990
rect 6500 1980 6550 1990
rect 7750 1980 7950 1990
rect 8600 1980 9050 1990
rect 3250 1970 3350 1980
rect 4800 1970 4850 1980
rect 5000 1970 5250 1980
rect 6100 1970 6350 1980
rect 6500 1970 6550 1980
rect 7750 1970 7950 1980
rect 8600 1970 9050 1980
rect 3250 1960 3350 1970
rect 4800 1960 4850 1970
rect 5000 1960 5250 1970
rect 6100 1960 6350 1970
rect 6500 1960 6550 1970
rect 7750 1960 7950 1970
rect 8600 1960 9050 1970
rect 3250 1950 3350 1960
rect 4800 1950 4850 1960
rect 5000 1950 5250 1960
rect 6100 1950 6350 1960
rect 6500 1950 6550 1960
rect 7750 1950 7950 1960
rect 8600 1950 9050 1960
rect 3300 1940 3350 1950
rect 4450 1940 4500 1950
rect 4550 1940 4700 1950
rect 4850 1940 4900 1950
rect 4950 1940 5000 1950
rect 6100 1940 6200 1950
rect 6300 1940 6350 1950
rect 6500 1940 6550 1950
rect 7750 1940 7800 1950
rect 3300 1930 3350 1940
rect 4450 1930 4500 1940
rect 4550 1930 4700 1940
rect 4850 1930 4900 1940
rect 4950 1930 5000 1940
rect 6100 1930 6200 1940
rect 6300 1930 6350 1940
rect 6500 1930 6550 1940
rect 7750 1930 7800 1940
rect 3300 1920 3350 1930
rect 4450 1920 4500 1930
rect 4550 1920 4700 1930
rect 4850 1920 4900 1930
rect 4950 1920 5000 1930
rect 6100 1920 6200 1930
rect 6300 1920 6350 1930
rect 6500 1920 6550 1930
rect 7750 1920 7800 1930
rect 3300 1910 3350 1920
rect 4450 1910 4500 1920
rect 4550 1910 4700 1920
rect 4850 1910 4900 1920
rect 4950 1910 5000 1920
rect 6100 1910 6200 1920
rect 6300 1910 6350 1920
rect 6500 1910 6550 1920
rect 7750 1910 7800 1920
rect 3300 1900 3350 1910
rect 4450 1900 4500 1910
rect 4550 1900 4700 1910
rect 4850 1900 4900 1910
rect 4950 1900 5000 1910
rect 6100 1900 6200 1910
rect 6300 1900 6350 1910
rect 6500 1900 6550 1910
rect 7750 1900 7800 1910
rect 2500 1890 2750 1900
rect 3300 1890 3350 1900
rect 4350 1890 4450 1900
rect 4500 1890 4750 1900
rect 4800 1890 4850 1900
rect 4900 1890 4950 1900
rect 6050 1890 6200 1900
rect 6300 1890 6400 1900
rect 6450 1890 6550 1900
rect 7750 1890 7800 1900
rect 2500 1880 2750 1890
rect 3300 1880 3350 1890
rect 4350 1880 4450 1890
rect 4500 1880 4750 1890
rect 4800 1880 4850 1890
rect 4900 1880 4950 1890
rect 6050 1880 6200 1890
rect 6300 1880 6400 1890
rect 6450 1880 6550 1890
rect 7750 1880 7800 1890
rect 2500 1870 2750 1880
rect 3300 1870 3350 1880
rect 4350 1870 4450 1880
rect 4500 1870 4750 1880
rect 4800 1870 4850 1880
rect 4900 1870 4950 1880
rect 6050 1870 6200 1880
rect 6300 1870 6400 1880
rect 6450 1870 6550 1880
rect 7750 1870 7800 1880
rect 2500 1860 2750 1870
rect 3300 1860 3350 1870
rect 4350 1860 4450 1870
rect 4500 1860 4750 1870
rect 4800 1860 4850 1870
rect 4900 1860 4950 1870
rect 6050 1860 6200 1870
rect 6300 1860 6400 1870
rect 6450 1860 6550 1870
rect 7750 1860 7800 1870
rect 2500 1850 2750 1860
rect 3300 1850 3350 1860
rect 4350 1850 4450 1860
rect 4500 1850 4750 1860
rect 4800 1850 4850 1860
rect 4900 1850 4950 1860
rect 6050 1850 6200 1860
rect 6300 1850 6400 1860
rect 6450 1850 6550 1860
rect 7750 1850 7800 1860
rect 2350 1840 2450 1850
rect 2750 1840 2850 1850
rect 4100 1840 4200 1850
rect 4500 1840 4550 1850
rect 4650 1840 4750 1850
rect 4900 1840 4950 1850
rect 6000 1840 6150 1850
rect 6250 1840 6350 1850
rect 6450 1840 6500 1850
rect 7750 1840 7800 1850
rect 9150 1840 9200 1850
rect 2350 1830 2450 1840
rect 2750 1830 2850 1840
rect 4100 1830 4200 1840
rect 4500 1830 4550 1840
rect 4650 1830 4750 1840
rect 4900 1830 4950 1840
rect 6000 1830 6150 1840
rect 6250 1830 6350 1840
rect 6450 1830 6500 1840
rect 7750 1830 7800 1840
rect 9150 1830 9200 1840
rect 2350 1820 2450 1830
rect 2750 1820 2850 1830
rect 4100 1820 4200 1830
rect 4500 1820 4550 1830
rect 4650 1820 4750 1830
rect 4900 1820 4950 1830
rect 6000 1820 6150 1830
rect 6250 1820 6350 1830
rect 6450 1820 6500 1830
rect 7750 1820 7800 1830
rect 9150 1820 9200 1830
rect 2350 1810 2450 1820
rect 2750 1810 2850 1820
rect 4100 1810 4200 1820
rect 4500 1810 4550 1820
rect 4650 1810 4750 1820
rect 4900 1810 4950 1820
rect 6000 1810 6150 1820
rect 6250 1810 6350 1820
rect 6450 1810 6500 1820
rect 7750 1810 7800 1820
rect 9150 1810 9200 1820
rect 2350 1800 2450 1810
rect 2750 1800 2850 1810
rect 4100 1800 4200 1810
rect 4500 1800 4550 1810
rect 4650 1800 4750 1810
rect 4900 1800 4950 1810
rect 6000 1800 6150 1810
rect 6250 1800 6350 1810
rect 6450 1800 6500 1810
rect 7750 1800 7800 1810
rect 9150 1800 9200 1810
rect 1850 1790 1900 1800
rect 2450 1790 2500 1800
rect 4200 1790 4250 1800
rect 4350 1790 4400 1800
rect 4500 1790 4700 1800
rect 4900 1790 4950 1800
rect 5200 1790 5250 1800
rect 5950 1790 6100 1800
rect 6250 1790 6350 1800
rect 6450 1790 6550 1800
rect 7800 1790 7850 1800
rect 8400 1790 8450 1800
rect 9100 1790 9200 1800
rect 1850 1780 1900 1790
rect 2450 1780 2500 1790
rect 4200 1780 4250 1790
rect 4350 1780 4400 1790
rect 4500 1780 4700 1790
rect 4900 1780 4950 1790
rect 5200 1780 5250 1790
rect 5950 1780 6100 1790
rect 6250 1780 6350 1790
rect 6450 1780 6550 1790
rect 7800 1780 7850 1790
rect 8400 1780 8450 1790
rect 9100 1780 9200 1790
rect 1850 1770 1900 1780
rect 2450 1770 2500 1780
rect 4200 1770 4250 1780
rect 4350 1770 4400 1780
rect 4500 1770 4700 1780
rect 4900 1770 4950 1780
rect 5200 1770 5250 1780
rect 5950 1770 6100 1780
rect 6250 1770 6350 1780
rect 6450 1770 6550 1780
rect 7800 1770 7850 1780
rect 8400 1770 8450 1780
rect 9100 1770 9200 1780
rect 1850 1760 1900 1770
rect 2450 1760 2500 1770
rect 4200 1760 4250 1770
rect 4350 1760 4400 1770
rect 4500 1760 4700 1770
rect 4900 1760 4950 1770
rect 5200 1760 5250 1770
rect 5950 1760 6100 1770
rect 6250 1760 6350 1770
rect 6450 1760 6550 1770
rect 7800 1760 7850 1770
rect 8400 1760 8450 1770
rect 9100 1760 9200 1770
rect 1850 1750 1900 1760
rect 2450 1750 2500 1760
rect 4200 1750 4250 1760
rect 4350 1750 4400 1760
rect 4500 1750 4700 1760
rect 4900 1750 4950 1760
rect 5200 1750 5250 1760
rect 5950 1750 6100 1760
rect 6250 1750 6350 1760
rect 6450 1750 6550 1760
rect 7800 1750 7850 1760
rect 8400 1750 8450 1760
rect 9100 1750 9200 1760
rect 1850 1740 1900 1750
rect 3250 1740 3300 1750
rect 4250 1740 4300 1750
rect 4350 1740 4400 1750
rect 4650 1740 4700 1750
rect 5150 1740 5200 1750
rect 5950 1740 6050 1750
rect 6300 1740 6350 1750
rect 6450 1740 6550 1750
rect 6800 1740 6850 1750
rect 7800 1740 7850 1750
rect 8400 1740 8450 1750
rect 9150 1740 9200 1750
rect 1850 1730 1900 1740
rect 3250 1730 3300 1740
rect 4250 1730 4300 1740
rect 4350 1730 4400 1740
rect 4650 1730 4700 1740
rect 5150 1730 5200 1740
rect 5950 1730 6050 1740
rect 6300 1730 6350 1740
rect 6450 1730 6550 1740
rect 6800 1730 6850 1740
rect 7800 1730 7850 1740
rect 8400 1730 8450 1740
rect 9150 1730 9200 1740
rect 1850 1720 1900 1730
rect 3250 1720 3300 1730
rect 4250 1720 4300 1730
rect 4350 1720 4400 1730
rect 4650 1720 4700 1730
rect 5150 1720 5200 1730
rect 5950 1720 6050 1730
rect 6300 1720 6350 1730
rect 6450 1720 6550 1730
rect 6800 1720 6850 1730
rect 7800 1720 7850 1730
rect 8400 1720 8450 1730
rect 9150 1720 9200 1730
rect 1850 1710 1900 1720
rect 3250 1710 3300 1720
rect 4250 1710 4300 1720
rect 4350 1710 4400 1720
rect 4650 1710 4700 1720
rect 5150 1710 5200 1720
rect 5950 1710 6050 1720
rect 6300 1710 6350 1720
rect 6450 1710 6550 1720
rect 6800 1710 6850 1720
rect 7800 1710 7850 1720
rect 8400 1710 8450 1720
rect 9150 1710 9200 1720
rect 1850 1700 1900 1710
rect 3250 1700 3300 1710
rect 4250 1700 4300 1710
rect 4350 1700 4400 1710
rect 4650 1700 4700 1710
rect 5150 1700 5200 1710
rect 5950 1700 6050 1710
rect 6300 1700 6350 1710
rect 6450 1700 6550 1710
rect 6800 1700 6850 1710
rect 7800 1700 7850 1710
rect 8400 1700 8450 1710
rect 9150 1700 9200 1710
rect 4250 1690 4300 1700
rect 4350 1690 4450 1700
rect 4500 1690 4600 1700
rect 5900 1690 6050 1700
rect 6300 1690 6400 1700
rect 6450 1690 6550 1700
rect 6800 1690 6850 1700
rect 7350 1690 7400 1700
rect 7800 1690 7850 1700
rect 8350 1690 8450 1700
rect 9150 1690 9200 1700
rect 4250 1680 4300 1690
rect 4350 1680 4450 1690
rect 4500 1680 4600 1690
rect 5900 1680 6050 1690
rect 6300 1680 6400 1690
rect 6450 1680 6550 1690
rect 6800 1680 6850 1690
rect 7350 1680 7400 1690
rect 7800 1680 7850 1690
rect 8350 1680 8450 1690
rect 9150 1680 9200 1690
rect 4250 1670 4300 1680
rect 4350 1670 4450 1680
rect 4500 1670 4600 1680
rect 5900 1670 6050 1680
rect 6300 1670 6400 1680
rect 6450 1670 6550 1680
rect 6800 1670 6850 1680
rect 7350 1670 7400 1680
rect 7800 1670 7850 1680
rect 8350 1670 8450 1680
rect 9150 1670 9200 1680
rect 4250 1660 4300 1670
rect 4350 1660 4450 1670
rect 4500 1660 4600 1670
rect 5900 1660 6050 1670
rect 6300 1660 6400 1670
rect 6450 1660 6550 1670
rect 6800 1660 6850 1670
rect 7350 1660 7400 1670
rect 7800 1660 7850 1670
rect 8350 1660 8450 1670
rect 9150 1660 9200 1670
rect 4250 1650 4300 1660
rect 4350 1650 4450 1660
rect 4500 1650 4600 1660
rect 5900 1650 6050 1660
rect 6300 1650 6400 1660
rect 6450 1650 6550 1660
rect 6800 1650 6850 1660
rect 7350 1650 7400 1660
rect 7800 1650 7850 1660
rect 8350 1650 8450 1660
rect 9150 1650 9200 1660
rect 1900 1640 1950 1650
rect 3200 1640 3250 1650
rect 4100 1640 4150 1650
rect 4300 1640 4550 1650
rect 4600 1640 4950 1650
rect 5900 1640 6000 1650
rect 6300 1640 6500 1650
rect 7350 1640 7400 1650
rect 7800 1640 7850 1650
rect 8350 1640 8400 1650
rect 1900 1630 1950 1640
rect 3200 1630 3250 1640
rect 4100 1630 4150 1640
rect 4300 1630 4550 1640
rect 4600 1630 4950 1640
rect 5900 1630 6000 1640
rect 6300 1630 6500 1640
rect 7350 1630 7400 1640
rect 7800 1630 7850 1640
rect 8350 1630 8400 1640
rect 1900 1620 1950 1630
rect 3200 1620 3250 1630
rect 4100 1620 4150 1630
rect 4300 1620 4550 1630
rect 4600 1620 4950 1630
rect 5900 1620 6000 1630
rect 6300 1620 6500 1630
rect 7350 1620 7400 1630
rect 7800 1620 7850 1630
rect 8350 1620 8400 1630
rect 1900 1610 1950 1620
rect 3200 1610 3250 1620
rect 4100 1610 4150 1620
rect 4300 1610 4550 1620
rect 4600 1610 4950 1620
rect 5900 1610 6000 1620
rect 6300 1610 6500 1620
rect 7350 1610 7400 1620
rect 7800 1610 7850 1620
rect 8350 1610 8400 1620
rect 1900 1600 1950 1610
rect 3200 1600 3250 1610
rect 4100 1600 4150 1610
rect 4300 1600 4550 1610
rect 4600 1600 4950 1610
rect 5900 1600 6000 1610
rect 6300 1600 6500 1610
rect 7350 1600 7400 1610
rect 7800 1600 7850 1610
rect 8350 1600 8400 1610
rect 3150 1590 3200 1600
rect 4100 1590 4150 1600
rect 4800 1590 5100 1600
rect 5800 1590 5850 1600
rect 5900 1590 6000 1600
rect 6300 1590 6450 1600
rect 7350 1590 7400 1600
rect 7800 1590 7850 1600
rect 8350 1590 8400 1600
rect 3150 1580 3200 1590
rect 4100 1580 4150 1590
rect 4800 1580 5100 1590
rect 5800 1580 5850 1590
rect 5900 1580 6000 1590
rect 6300 1580 6450 1590
rect 7350 1580 7400 1590
rect 7800 1580 7850 1590
rect 8350 1580 8400 1590
rect 3150 1570 3200 1580
rect 4100 1570 4150 1580
rect 4800 1570 5100 1580
rect 5800 1570 5850 1580
rect 5900 1570 6000 1580
rect 6300 1570 6450 1580
rect 7350 1570 7400 1580
rect 7800 1570 7850 1580
rect 8350 1570 8400 1580
rect 3150 1560 3200 1570
rect 4100 1560 4150 1570
rect 4800 1560 5100 1570
rect 5800 1560 5850 1570
rect 5900 1560 6000 1570
rect 6300 1560 6450 1570
rect 7350 1560 7400 1570
rect 7800 1560 7850 1570
rect 8350 1560 8400 1570
rect 3150 1550 3200 1560
rect 4100 1550 4150 1560
rect 4800 1550 5100 1560
rect 5800 1550 5850 1560
rect 5900 1550 6000 1560
rect 6300 1550 6450 1560
rect 7350 1550 7400 1560
rect 7800 1550 7850 1560
rect 8350 1550 8400 1560
rect 1950 1540 2000 1550
rect 3100 1540 3150 1550
rect 4100 1540 4150 1550
rect 4850 1540 5250 1550
rect 5350 1540 5400 1550
rect 5800 1540 6000 1550
rect 6300 1540 6400 1550
rect 7350 1540 7400 1550
rect 7800 1540 7850 1550
rect 8300 1540 8400 1550
rect 9750 1540 9800 1550
rect 1950 1530 2000 1540
rect 3100 1530 3150 1540
rect 4100 1530 4150 1540
rect 4850 1530 5250 1540
rect 5350 1530 5400 1540
rect 5800 1530 6000 1540
rect 6300 1530 6400 1540
rect 7350 1530 7400 1540
rect 7800 1530 7850 1540
rect 8300 1530 8400 1540
rect 9750 1530 9800 1540
rect 1950 1520 2000 1530
rect 3100 1520 3150 1530
rect 4100 1520 4150 1530
rect 4850 1520 5250 1530
rect 5350 1520 5400 1530
rect 5800 1520 6000 1530
rect 6300 1520 6400 1530
rect 7350 1520 7400 1530
rect 7800 1520 7850 1530
rect 8300 1520 8400 1530
rect 9750 1520 9800 1530
rect 1950 1510 2000 1520
rect 3100 1510 3150 1520
rect 4100 1510 4150 1520
rect 4850 1510 5250 1520
rect 5350 1510 5400 1520
rect 5800 1510 6000 1520
rect 6300 1510 6400 1520
rect 7350 1510 7400 1520
rect 7800 1510 7850 1520
rect 8300 1510 8400 1520
rect 9750 1510 9800 1520
rect 1950 1500 2000 1510
rect 3100 1500 3150 1510
rect 4100 1500 4150 1510
rect 4850 1500 5250 1510
rect 5350 1500 5400 1510
rect 5800 1500 6000 1510
rect 6300 1500 6400 1510
rect 7350 1500 7400 1510
rect 7800 1500 7850 1510
rect 8300 1500 8400 1510
rect 9750 1500 9800 1510
rect 900 1490 950 1500
rect 2000 1490 2050 1500
rect 3050 1490 3100 1500
rect 4100 1490 4150 1500
rect 4950 1490 5400 1500
rect 5800 1490 5950 1500
rect 6350 1490 6400 1500
rect 7800 1490 7850 1500
rect 8300 1490 8400 1500
rect 9750 1490 9800 1500
rect 900 1480 950 1490
rect 2000 1480 2050 1490
rect 3050 1480 3100 1490
rect 4100 1480 4150 1490
rect 4950 1480 5400 1490
rect 5800 1480 5950 1490
rect 6350 1480 6400 1490
rect 7800 1480 7850 1490
rect 8300 1480 8400 1490
rect 9750 1480 9800 1490
rect 900 1470 950 1480
rect 2000 1470 2050 1480
rect 3050 1470 3100 1480
rect 4100 1470 4150 1480
rect 4950 1470 5400 1480
rect 5800 1470 5950 1480
rect 6350 1470 6400 1480
rect 7800 1470 7850 1480
rect 8300 1470 8400 1480
rect 9750 1470 9800 1480
rect 900 1460 950 1470
rect 2000 1460 2050 1470
rect 3050 1460 3100 1470
rect 4100 1460 4150 1470
rect 4950 1460 5400 1470
rect 5800 1460 5950 1470
rect 6350 1460 6400 1470
rect 7800 1460 7850 1470
rect 8300 1460 8400 1470
rect 9750 1460 9800 1470
rect 900 1450 950 1460
rect 2000 1450 2050 1460
rect 3050 1450 3100 1460
rect 4100 1450 4150 1460
rect 4950 1450 5400 1460
rect 5800 1450 5950 1460
rect 6350 1450 6400 1460
rect 7800 1450 7850 1460
rect 8300 1450 8400 1460
rect 9750 1450 9800 1460
rect 850 1440 900 1450
rect 950 1440 1000 1450
rect 2050 1440 2100 1450
rect 2950 1440 3050 1450
rect 4950 1440 5400 1450
rect 5850 1440 5950 1450
rect 7850 1440 7900 1450
rect 8300 1440 8400 1450
rect 9700 1440 9750 1450
rect 850 1430 900 1440
rect 950 1430 1000 1440
rect 2050 1430 2100 1440
rect 2950 1430 3050 1440
rect 4950 1430 5400 1440
rect 5850 1430 5950 1440
rect 7850 1430 7900 1440
rect 8300 1430 8400 1440
rect 9700 1430 9750 1440
rect 850 1420 900 1430
rect 950 1420 1000 1430
rect 2050 1420 2100 1430
rect 2950 1420 3050 1430
rect 4950 1420 5400 1430
rect 5850 1420 5950 1430
rect 7850 1420 7900 1430
rect 8300 1420 8400 1430
rect 9700 1420 9750 1430
rect 850 1410 900 1420
rect 950 1410 1000 1420
rect 2050 1410 2100 1420
rect 2950 1410 3050 1420
rect 4950 1410 5400 1420
rect 5850 1410 5950 1420
rect 7850 1410 7900 1420
rect 8300 1410 8400 1420
rect 9700 1410 9750 1420
rect 850 1400 900 1410
rect 950 1400 1000 1410
rect 2050 1400 2100 1410
rect 2950 1400 3050 1410
rect 4950 1400 5400 1410
rect 5850 1400 5950 1410
rect 7850 1400 7900 1410
rect 8300 1400 8400 1410
rect 9700 1400 9750 1410
rect 800 1390 1000 1400
rect 2100 1390 2150 1400
rect 2850 1390 3000 1400
rect 3550 1390 3650 1400
rect 4150 1390 4200 1400
rect 4400 1390 4450 1400
rect 5100 1390 5450 1400
rect 5850 1390 5950 1400
rect 7850 1390 7900 1400
rect 8250 1390 8400 1400
rect 9700 1390 9750 1400
rect 800 1380 1000 1390
rect 2100 1380 2150 1390
rect 2850 1380 3000 1390
rect 3550 1380 3650 1390
rect 4150 1380 4200 1390
rect 4400 1380 4450 1390
rect 5100 1380 5450 1390
rect 5850 1380 5950 1390
rect 7850 1380 7900 1390
rect 8250 1380 8400 1390
rect 9700 1380 9750 1390
rect 800 1370 1000 1380
rect 2100 1370 2150 1380
rect 2850 1370 3000 1380
rect 3550 1370 3650 1380
rect 4150 1370 4200 1380
rect 4400 1370 4450 1380
rect 5100 1370 5450 1380
rect 5850 1370 5950 1380
rect 7850 1370 7900 1380
rect 8250 1370 8400 1380
rect 9700 1370 9750 1380
rect 800 1360 1000 1370
rect 2100 1360 2150 1370
rect 2850 1360 3000 1370
rect 3550 1360 3650 1370
rect 4150 1360 4200 1370
rect 4400 1360 4450 1370
rect 5100 1360 5450 1370
rect 5850 1360 5950 1370
rect 7850 1360 7900 1370
rect 8250 1360 8400 1370
rect 9700 1360 9750 1370
rect 800 1350 1000 1360
rect 2100 1350 2150 1360
rect 2850 1350 3000 1360
rect 3550 1350 3650 1360
rect 4150 1350 4200 1360
rect 4400 1350 4450 1360
rect 5100 1350 5450 1360
rect 5850 1350 5950 1360
rect 7850 1350 7900 1360
rect 8250 1350 8400 1360
rect 9700 1350 9750 1360
rect 800 1340 950 1350
rect 2100 1340 2200 1350
rect 2800 1340 2850 1350
rect 4150 1340 4200 1350
rect 4950 1340 5700 1350
rect 5850 1340 5950 1350
rect 7850 1340 7900 1350
rect 8250 1340 8350 1350
rect 800 1330 950 1340
rect 2100 1330 2200 1340
rect 2800 1330 2850 1340
rect 4150 1330 4200 1340
rect 4950 1330 5700 1340
rect 5850 1330 5950 1340
rect 7850 1330 7900 1340
rect 8250 1330 8350 1340
rect 800 1320 950 1330
rect 2100 1320 2200 1330
rect 2800 1320 2850 1330
rect 4150 1320 4200 1330
rect 4950 1320 5700 1330
rect 5850 1320 5950 1330
rect 7850 1320 7900 1330
rect 8250 1320 8350 1330
rect 800 1310 950 1320
rect 2100 1310 2200 1320
rect 2800 1310 2850 1320
rect 4150 1310 4200 1320
rect 4950 1310 5700 1320
rect 5850 1310 5950 1320
rect 7850 1310 7900 1320
rect 8250 1310 8350 1320
rect 800 1300 950 1310
rect 2100 1300 2200 1310
rect 2800 1300 2850 1310
rect 4150 1300 4200 1310
rect 4950 1300 5700 1310
rect 5850 1300 5950 1310
rect 7850 1300 7900 1310
rect 8250 1300 8350 1310
rect 800 1290 950 1300
rect 2150 1290 2250 1300
rect 2700 1290 2800 1300
rect 4150 1290 4200 1300
rect 4950 1290 5250 1300
rect 5450 1290 5750 1300
rect 5850 1290 5950 1300
rect 7850 1290 7900 1300
rect 9150 1290 9250 1300
rect 800 1280 950 1290
rect 2150 1280 2250 1290
rect 2700 1280 2800 1290
rect 4150 1280 4200 1290
rect 4950 1280 5250 1290
rect 5450 1280 5750 1290
rect 5850 1280 5950 1290
rect 7850 1280 7900 1290
rect 9150 1280 9250 1290
rect 800 1270 950 1280
rect 2150 1270 2250 1280
rect 2700 1270 2800 1280
rect 4150 1270 4200 1280
rect 4950 1270 5250 1280
rect 5450 1270 5750 1280
rect 5850 1270 5950 1280
rect 7850 1270 7900 1280
rect 9150 1270 9250 1280
rect 800 1260 950 1270
rect 2150 1260 2250 1270
rect 2700 1260 2800 1270
rect 4150 1260 4200 1270
rect 4950 1260 5250 1270
rect 5450 1260 5750 1270
rect 5850 1260 5950 1270
rect 7850 1260 7900 1270
rect 9150 1260 9250 1270
rect 800 1250 950 1260
rect 2150 1250 2250 1260
rect 2700 1250 2800 1260
rect 4150 1250 4200 1260
rect 4950 1250 5250 1260
rect 5450 1250 5750 1260
rect 5850 1250 5950 1260
rect 7850 1250 7900 1260
rect 9150 1250 9250 1260
rect 800 1240 950 1250
rect 2100 1240 2700 1250
rect 3800 1240 3850 1250
rect 4450 1240 4500 1250
rect 4750 1240 5000 1250
rect 5600 1240 5750 1250
rect 5850 1240 5950 1250
rect 6700 1240 6800 1250
rect 7850 1240 7900 1250
rect 9150 1240 9250 1250
rect 9750 1240 9800 1250
rect 800 1230 950 1240
rect 2100 1230 2700 1240
rect 3800 1230 3850 1240
rect 4450 1230 4500 1240
rect 4750 1230 5000 1240
rect 5600 1230 5750 1240
rect 5850 1230 5950 1240
rect 6700 1230 6800 1240
rect 7850 1230 7900 1240
rect 9150 1230 9250 1240
rect 9750 1230 9800 1240
rect 800 1220 950 1230
rect 2100 1220 2700 1230
rect 3800 1220 3850 1230
rect 4450 1220 4500 1230
rect 4750 1220 5000 1230
rect 5600 1220 5750 1230
rect 5850 1220 5950 1230
rect 6700 1220 6800 1230
rect 7850 1220 7900 1230
rect 9150 1220 9250 1230
rect 9750 1220 9800 1230
rect 800 1210 950 1220
rect 2100 1210 2700 1220
rect 3800 1210 3850 1220
rect 4450 1210 4500 1220
rect 4750 1210 5000 1220
rect 5600 1210 5750 1220
rect 5850 1210 5950 1220
rect 6700 1210 6800 1220
rect 7850 1210 7900 1220
rect 9150 1210 9250 1220
rect 9750 1210 9800 1220
rect 800 1200 950 1210
rect 2100 1200 2700 1210
rect 3800 1200 3850 1210
rect 4450 1200 4500 1210
rect 4750 1200 5000 1210
rect 5600 1200 5750 1210
rect 5850 1200 5950 1210
rect 6700 1200 6800 1210
rect 7850 1200 7900 1210
rect 9150 1200 9250 1210
rect 9750 1200 9800 1210
rect 750 1190 800 1200
rect 850 1190 900 1200
rect 2050 1190 2600 1200
rect 3550 1190 3600 1200
rect 4450 1190 4500 1200
rect 4550 1190 4700 1200
rect 4900 1190 5000 1200
rect 5050 1190 5400 1200
rect 5600 1190 5950 1200
rect 6600 1190 6650 1200
rect 7900 1190 7950 1200
rect 9150 1190 9250 1200
rect 9750 1190 9800 1200
rect 750 1180 800 1190
rect 850 1180 900 1190
rect 2050 1180 2600 1190
rect 3550 1180 3600 1190
rect 4450 1180 4500 1190
rect 4550 1180 4700 1190
rect 4900 1180 5000 1190
rect 5050 1180 5400 1190
rect 5600 1180 5950 1190
rect 6600 1180 6650 1190
rect 7900 1180 7950 1190
rect 9150 1180 9250 1190
rect 9750 1180 9800 1190
rect 750 1170 800 1180
rect 850 1170 900 1180
rect 2050 1170 2600 1180
rect 3550 1170 3600 1180
rect 4450 1170 4500 1180
rect 4550 1170 4700 1180
rect 4900 1170 5000 1180
rect 5050 1170 5400 1180
rect 5600 1170 5950 1180
rect 6600 1170 6650 1180
rect 7900 1170 7950 1180
rect 9150 1170 9250 1180
rect 9750 1170 9800 1180
rect 750 1160 800 1170
rect 850 1160 900 1170
rect 2050 1160 2600 1170
rect 3550 1160 3600 1170
rect 4450 1160 4500 1170
rect 4550 1160 4700 1170
rect 4900 1160 5000 1170
rect 5050 1160 5400 1170
rect 5600 1160 5950 1170
rect 6600 1160 6650 1170
rect 7900 1160 7950 1170
rect 9150 1160 9250 1170
rect 9750 1160 9800 1170
rect 750 1150 800 1160
rect 850 1150 900 1160
rect 2050 1150 2600 1160
rect 3550 1150 3600 1160
rect 4450 1150 4500 1160
rect 4550 1150 4700 1160
rect 4900 1150 5000 1160
rect 5050 1150 5400 1160
rect 5600 1150 5950 1160
rect 6600 1150 6650 1160
rect 7900 1150 7950 1160
rect 9150 1150 9250 1160
rect 9750 1150 9800 1160
rect 850 1140 900 1150
rect 2000 1140 2100 1150
rect 2250 1140 2400 1150
rect 2550 1140 2800 1150
rect 3600 1140 3650 1150
rect 3950 1140 4000 1150
rect 4550 1140 4900 1150
rect 5350 1140 5950 1150
rect 6500 1140 6600 1150
rect 7400 1140 7450 1150
rect 7900 1140 7950 1150
rect 9750 1140 9800 1150
rect 850 1130 900 1140
rect 2000 1130 2100 1140
rect 2250 1130 2400 1140
rect 2550 1130 2800 1140
rect 3600 1130 3650 1140
rect 3950 1130 4000 1140
rect 4550 1130 4900 1140
rect 5350 1130 5950 1140
rect 6500 1130 6600 1140
rect 7400 1130 7450 1140
rect 7900 1130 7950 1140
rect 9750 1130 9800 1140
rect 850 1120 900 1130
rect 2000 1120 2100 1130
rect 2250 1120 2400 1130
rect 2550 1120 2800 1130
rect 3600 1120 3650 1130
rect 3950 1120 4000 1130
rect 4550 1120 4900 1130
rect 5350 1120 5950 1130
rect 6500 1120 6600 1130
rect 7400 1120 7450 1130
rect 7900 1120 7950 1130
rect 9750 1120 9800 1130
rect 850 1110 900 1120
rect 2000 1110 2100 1120
rect 2250 1110 2400 1120
rect 2550 1110 2800 1120
rect 3600 1110 3650 1120
rect 3950 1110 4000 1120
rect 4550 1110 4900 1120
rect 5350 1110 5950 1120
rect 6500 1110 6600 1120
rect 7400 1110 7450 1120
rect 7900 1110 7950 1120
rect 9750 1110 9800 1120
rect 850 1100 900 1110
rect 2000 1100 2100 1110
rect 2250 1100 2400 1110
rect 2550 1100 2800 1110
rect 3600 1100 3650 1110
rect 3950 1100 4000 1110
rect 4550 1100 4900 1110
rect 5350 1100 5950 1110
rect 6500 1100 6600 1110
rect 7400 1100 7450 1110
rect 7900 1100 7950 1110
rect 9750 1100 9800 1110
rect 850 1090 900 1100
rect 1600 1090 1650 1100
rect 2000 1090 2050 1100
rect 2300 1090 2850 1100
rect 4500 1090 4650 1100
rect 5450 1090 5700 1100
rect 5800 1090 6000 1100
rect 6450 1090 6500 1100
rect 7400 1090 7450 1100
rect 7900 1090 7950 1100
rect 9000 1090 9050 1100
rect 9750 1090 9800 1100
rect 850 1080 900 1090
rect 1600 1080 1650 1090
rect 2000 1080 2050 1090
rect 2300 1080 2850 1090
rect 4500 1080 4650 1090
rect 5450 1080 5700 1090
rect 5800 1080 6000 1090
rect 6450 1080 6500 1090
rect 7400 1080 7450 1090
rect 7900 1080 7950 1090
rect 9000 1080 9050 1090
rect 9750 1080 9800 1090
rect 850 1070 900 1080
rect 1600 1070 1650 1080
rect 2000 1070 2050 1080
rect 2300 1070 2850 1080
rect 4500 1070 4650 1080
rect 5450 1070 5700 1080
rect 5800 1070 6000 1080
rect 6450 1070 6500 1080
rect 7400 1070 7450 1080
rect 7900 1070 7950 1080
rect 9000 1070 9050 1080
rect 9750 1070 9800 1080
rect 850 1060 900 1070
rect 1600 1060 1650 1070
rect 2000 1060 2050 1070
rect 2300 1060 2850 1070
rect 4500 1060 4650 1070
rect 5450 1060 5700 1070
rect 5800 1060 6000 1070
rect 6450 1060 6500 1070
rect 7400 1060 7450 1070
rect 7900 1060 7950 1070
rect 9000 1060 9050 1070
rect 9750 1060 9800 1070
rect 850 1050 900 1060
rect 1600 1050 1650 1060
rect 2000 1050 2050 1060
rect 2300 1050 2850 1060
rect 4500 1050 4650 1060
rect 5450 1050 5700 1060
rect 5800 1050 6000 1060
rect 6450 1050 6500 1060
rect 7400 1050 7450 1060
rect 7900 1050 7950 1060
rect 9000 1050 9050 1060
rect 9750 1050 9800 1060
rect 700 1040 750 1050
rect 1550 1040 1650 1050
rect 2000 1040 2050 1050
rect 2800 1040 2850 1050
rect 4100 1040 4150 1050
rect 4700 1040 4750 1050
rect 5450 1040 5650 1050
rect 5800 1040 5950 1050
rect 6400 1040 6450 1050
rect 7400 1040 7450 1050
rect 7900 1040 7950 1050
rect 8150 1040 8250 1050
rect 8900 1040 9100 1050
rect 700 1030 750 1040
rect 1550 1030 1650 1040
rect 2000 1030 2050 1040
rect 2800 1030 2850 1040
rect 4100 1030 4150 1040
rect 4700 1030 4750 1040
rect 5450 1030 5650 1040
rect 5800 1030 5950 1040
rect 6400 1030 6450 1040
rect 7400 1030 7450 1040
rect 7900 1030 7950 1040
rect 8150 1030 8250 1040
rect 8900 1030 9100 1040
rect 700 1020 750 1030
rect 1550 1020 1650 1030
rect 2000 1020 2050 1030
rect 2800 1020 2850 1030
rect 4100 1020 4150 1030
rect 4700 1020 4750 1030
rect 5450 1020 5650 1030
rect 5800 1020 5950 1030
rect 6400 1020 6450 1030
rect 7400 1020 7450 1030
rect 7900 1020 7950 1030
rect 8150 1020 8250 1030
rect 8900 1020 9100 1030
rect 700 1010 750 1020
rect 1550 1010 1650 1020
rect 2000 1010 2050 1020
rect 2800 1010 2850 1020
rect 4100 1010 4150 1020
rect 4700 1010 4750 1020
rect 5450 1010 5650 1020
rect 5800 1010 5950 1020
rect 6400 1010 6450 1020
rect 7400 1010 7450 1020
rect 7900 1010 7950 1020
rect 8150 1010 8250 1020
rect 8900 1010 9100 1020
rect 700 1000 750 1010
rect 1550 1000 1650 1010
rect 2000 1000 2050 1010
rect 2800 1000 2850 1010
rect 4100 1000 4150 1010
rect 4700 1000 4750 1010
rect 5450 1000 5650 1010
rect 5800 1000 5950 1010
rect 6400 1000 6450 1010
rect 7400 1000 7450 1010
rect 7900 1000 7950 1010
rect 8150 1000 8250 1010
rect 8900 1000 9100 1010
rect 800 990 850 1000
rect 1500 990 1550 1000
rect 2750 990 2850 1000
rect 4800 990 4850 1000
rect 5300 990 5450 1000
rect 5500 990 6000 1000
rect 6400 990 6450 1000
rect 7400 990 7450 1000
rect 7900 990 7950 1000
rect 8150 990 8250 1000
rect 8900 990 9100 1000
rect 800 980 850 990
rect 1500 980 1550 990
rect 2750 980 2850 990
rect 4800 980 4850 990
rect 5300 980 5450 990
rect 5500 980 6000 990
rect 6400 980 6450 990
rect 7400 980 7450 990
rect 7900 980 7950 990
rect 8150 980 8250 990
rect 8900 980 9100 990
rect 800 970 850 980
rect 1500 970 1550 980
rect 2750 970 2850 980
rect 4800 970 4850 980
rect 5300 970 5450 980
rect 5500 970 6000 980
rect 6400 970 6450 980
rect 7400 970 7450 980
rect 7900 970 7950 980
rect 8150 970 8250 980
rect 8900 970 9100 980
rect 800 960 850 970
rect 1500 960 1550 970
rect 2750 960 2850 970
rect 4800 960 4850 970
rect 5300 960 5450 970
rect 5500 960 6000 970
rect 6400 960 6450 970
rect 7400 960 7450 970
rect 7900 960 7950 970
rect 8150 960 8250 970
rect 8900 960 9100 970
rect 800 950 850 960
rect 1500 950 1550 960
rect 2750 950 2850 960
rect 4800 950 4850 960
rect 5300 950 5450 960
rect 5500 950 6000 960
rect 6400 950 6450 960
rect 7400 950 7450 960
rect 7900 950 7950 960
rect 8150 950 8250 960
rect 8900 950 9100 960
rect 650 940 700 950
rect 800 940 850 950
rect 1300 940 1350 950
rect 1450 940 1500 950
rect 2750 940 2800 950
rect 5300 940 5350 950
rect 5800 940 6050 950
rect 6200 940 6300 950
rect 6400 940 6450 950
rect 7400 940 7450 950
rect 8150 940 8250 950
rect 8850 940 8950 950
rect 9050 940 9100 950
rect 650 930 700 940
rect 800 930 850 940
rect 1300 930 1350 940
rect 1450 930 1500 940
rect 2750 930 2800 940
rect 5300 930 5350 940
rect 5800 930 6050 940
rect 6200 930 6300 940
rect 6400 930 6450 940
rect 7400 930 7450 940
rect 8150 930 8250 940
rect 8850 930 8950 940
rect 9050 930 9100 940
rect 650 920 700 930
rect 800 920 850 930
rect 1300 920 1350 930
rect 1450 920 1500 930
rect 2750 920 2800 930
rect 5300 920 5350 930
rect 5800 920 6050 930
rect 6200 920 6300 930
rect 6400 920 6450 930
rect 7400 920 7450 930
rect 8150 920 8250 930
rect 8850 920 8950 930
rect 9050 920 9100 930
rect 650 910 700 920
rect 800 910 850 920
rect 1300 910 1350 920
rect 1450 910 1500 920
rect 2750 910 2800 920
rect 5300 910 5350 920
rect 5800 910 6050 920
rect 6200 910 6300 920
rect 6400 910 6450 920
rect 7400 910 7450 920
rect 8150 910 8250 920
rect 8850 910 8950 920
rect 9050 910 9100 920
rect 650 900 700 910
rect 800 900 850 910
rect 1300 900 1350 910
rect 1450 900 1500 910
rect 2750 900 2800 910
rect 5300 900 5350 910
rect 5800 900 6050 910
rect 6200 900 6300 910
rect 6400 900 6450 910
rect 7400 900 7450 910
rect 8150 900 8250 910
rect 8850 900 8950 910
rect 9050 900 9100 910
rect 800 890 900 900
rect 1250 890 1300 900
rect 1400 890 1450 900
rect 2700 890 2750 900
rect 3800 890 3850 900
rect 5300 890 5350 900
rect 5500 890 6050 900
rect 6200 890 6300 900
rect 6400 890 6450 900
rect 7400 890 7450 900
rect 8150 890 8250 900
rect 8800 890 8900 900
rect 9050 890 9150 900
rect 800 880 900 890
rect 1250 880 1300 890
rect 1400 880 1450 890
rect 2700 880 2750 890
rect 3800 880 3850 890
rect 5300 880 5350 890
rect 5500 880 6050 890
rect 6200 880 6300 890
rect 6400 880 6450 890
rect 7400 880 7450 890
rect 8150 880 8250 890
rect 8800 880 8900 890
rect 9050 880 9150 890
rect 800 870 900 880
rect 1250 870 1300 880
rect 1400 870 1450 880
rect 2700 870 2750 880
rect 3800 870 3850 880
rect 5300 870 5350 880
rect 5500 870 6050 880
rect 6200 870 6300 880
rect 6400 870 6450 880
rect 7400 870 7450 880
rect 8150 870 8250 880
rect 8800 870 8900 880
rect 9050 870 9150 880
rect 800 860 900 870
rect 1250 860 1300 870
rect 1400 860 1450 870
rect 2700 860 2750 870
rect 3800 860 3850 870
rect 5300 860 5350 870
rect 5500 860 6050 870
rect 6200 860 6300 870
rect 6400 860 6450 870
rect 7400 860 7450 870
rect 8150 860 8250 870
rect 8800 860 8900 870
rect 9050 860 9150 870
rect 800 850 900 860
rect 1250 850 1300 860
rect 1400 850 1450 860
rect 2700 850 2750 860
rect 3800 850 3850 860
rect 5300 850 5350 860
rect 5500 850 6050 860
rect 6200 850 6300 860
rect 6400 850 6450 860
rect 7400 850 7450 860
rect 8150 850 8250 860
rect 8800 850 8900 860
rect 9050 850 9150 860
rect 600 840 650 850
rect 800 840 900 850
rect 1350 840 1400 850
rect 2000 840 2050 850
rect 3850 840 3900 850
rect 5350 840 5600 850
rect 5750 840 6050 850
rect 6150 840 6300 850
rect 7400 840 7450 850
rect 7950 840 8000 850
rect 8150 840 8300 850
rect 8750 840 8900 850
rect 9050 840 9150 850
rect 600 830 650 840
rect 800 830 900 840
rect 1350 830 1400 840
rect 2000 830 2050 840
rect 3850 830 3900 840
rect 5350 830 5600 840
rect 5750 830 6050 840
rect 6150 830 6300 840
rect 7400 830 7450 840
rect 7950 830 8000 840
rect 8150 830 8300 840
rect 8750 830 8900 840
rect 9050 830 9150 840
rect 600 820 650 830
rect 800 820 900 830
rect 1350 820 1400 830
rect 2000 820 2050 830
rect 3850 820 3900 830
rect 5350 820 5600 830
rect 5750 820 6050 830
rect 6150 820 6300 830
rect 7400 820 7450 830
rect 7950 820 8000 830
rect 8150 820 8300 830
rect 8750 820 8900 830
rect 9050 820 9150 830
rect 600 810 650 820
rect 800 810 900 820
rect 1350 810 1400 820
rect 2000 810 2050 820
rect 3850 810 3900 820
rect 5350 810 5600 820
rect 5750 810 6050 820
rect 6150 810 6300 820
rect 7400 810 7450 820
rect 7950 810 8000 820
rect 8150 810 8300 820
rect 8750 810 8900 820
rect 9050 810 9150 820
rect 600 800 650 810
rect 800 800 900 810
rect 1350 800 1400 810
rect 2000 800 2050 810
rect 3850 800 3900 810
rect 5350 800 5600 810
rect 5750 800 6050 810
rect 6150 800 6300 810
rect 7400 800 7450 810
rect 7950 800 8000 810
rect 8150 800 8300 810
rect 8750 800 8900 810
rect 9050 800 9150 810
rect 600 790 650 800
rect 750 790 850 800
rect 1100 790 1150 800
rect 1300 790 1350 800
rect 2550 790 2600 800
rect 3550 790 3600 800
rect 3850 790 4000 800
rect 4900 790 4950 800
rect 5450 790 5550 800
rect 5750 790 6300 800
rect 6450 790 6500 800
rect 7950 790 8000 800
rect 8200 790 8300 800
rect 8750 790 8850 800
rect 600 780 650 790
rect 750 780 850 790
rect 1100 780 1150 790
rect 1300 780 1350 790
rect 2550 780 2600 790
rect 3550 780 3600 790
rect 3850 780 4000 790
rect 4900 780 4950 790
rect 5450 780 5550 790
rect 5750 780 6300 790
rect 6450 780 6500 790
rect 7950 780 8000 790
rect 8200 780 8300 790
rect 8750 780 8850 790
rect 600 770 650 780
rect 750 770 850 780
rect 1100 770 1150 780
rect 1300 770 1350 780
rect 2550 770 2600 780
rect 3550 770 3600 780
rect 3850 770 4000 780
rect 4900 770 4950 780
rect 5450 770 5550 780
rect 5750 770 6300 780
rect 6450 770 6500 780
rect 7950 770 8000 780
rect 8200 770 8300 780
rect 8750 770 8850 780
rect 600 760 650 770
rect 750 760 850 770
rect 1100 760 1150 770
rect 1300 760 1350 770
rect 2550 760 2600 770
rect 3550 760 3600 770
rect 3850 760 4000 770
rect 4900 760 4950 770
rect 5450 760 5550 770
rect 5750 760 6300 770
rect 6450 760 6500 770
rect 7950 760 8000 770
rect 8200 760 8300 770
rect 8750 760 8850 770
rect 600 750 650 760
rect 750 750 850 760
rect 1100 750 1150 760
rect 1300 750 1350 760
rect 2550 750 2600 760
rect 3550 750 3600 760
rect 3850 750 4000 760
rect 4900 750 4950 760
rect 5450 750 5550 760
rect 5750 750 6300 760
rect 6450 750 6500 760
rect 7950 750 8000 760
rect 8200 750 8300 760
rect 8750 750 8850 760
rect 750 740 800 750
rect 1050 740 1100 750
rect 1250 740 1300 750
rect 2050 740 2100 750
rect 2450 740 2500 750
rect 3350 740 3400 750
rect 3950 740 4000 750
rect 5500 740 5550 750
rect 5750 740 6200 750
rect 6250 740 6300 750
rect 6450 740 6500 750
rect 7950 740 8000 750
rect 8200 740 8350 750
rect 8700 740 8800 750
rect 9150 740 9200 750
rect 750 730 800 740
rect 1050 730 1100 740
rect 1250 730 1300 740
rect 2050 730 2100 740
rect 2450 730 2500 740
rect 3350 730 3400 740
rect 3950 730 4000 740
rect 5500 730 5550 740
rect 5750 730 6200 740
rect 6250 730 6300 740
rect 6450 730 6500 740
rect 7950 730 8000 740
rect 8200 730 8350 740
rect 8700 730 8800 740
rect 9150 730 9200 740
rect 750 720 800 730
rect 1050 720 1100 730
rect 1250 720 1300 730
rect 2050 720 2100 730
rect 2450 720 2500 730
rect 3350 720 3400 730
rect 3950 720 4000 730
rect 5500 720 5550 730
rect 5750 720 6200 730
rect 6250 720 6300 730
rect 6450 720 6500 730
rect 7950 720 8000 730
rect 8200 720 8350 730
rect 8700 720 8800 730
rect 9150 720 9200 730
rect 750 710 800 720
rect 1050 710 1100 720
rect 1250 710 1300 720
rect 2050 710 2100 720
rect 2450 710 2500 720
rect 3350 710 3400 720
rect 3950 710 4000 720
rect 5500 710 5550 720
rect 5750 710 6200 720
rect 6250 710 6300 720
rect 6450 710 6500 720
rect 7950 710 8000 720
rect 8200 710 8350 720
rect 8700 710 8800 720
rect 9150 710 9200 720
rect 750 700 800 710
rect 1050 700 1100 710
rect 1250 700 1300 710
rect 2050 700 2100 710
rect 2450 700 2500 710
rect 3350 700 3400 710
rect 3950 700 4000 710
rect 5500 700 5550 710
rect 5750 700 6200 710
rect 6250 700 6300 710
rect 6450 700 6500 710
rect 7950 700 8000 710
rect 8200 700 8350 710
rect 8700 700 8800 710
rect 9150 700 9200 710
rect 550 690 600 700
rect 700 690 900 700
rect 950 690 1050 700
rect 1250 690 1300 700
rect 3250 690 3300 700
rect 4750 690 4800 700
rect 5500 690 5700 700
rect 5750 690 6050 700
rect 6150 690 6300 700
rect 6500 690 6550 700
rect 7350 690 7400 700
rect 8250 690 8400 700
rect 8650 690 8750 700
rect 9100 690 9150 700
rect 550 680 600 690
rect 700 680 900 690
rect 950 680 1050 690
rect 1250 680 1300 690
rect 3250 680 3300 690
rect 4750 680 4800 690
rect 5500 680 5700 690
rect 5750 680 6050 690
rect 6150 680 6300 690
rect 6500 680 6550 690
rect 7350 680 7400 690
rect 8250 680 8400 690
rect 8650 680 8750 690
rect 9100 680 9150 690
rect 550 670 600 680
rect 700 670 900 680
rect 950 670 1050 680
rect 1250 670 1300 680
rect 3250 670 3300 680
rect 4750 670 4800 680
rect 5500 670 5700 680
rect 5750 670 6050 680
rect 6150 670 6300 680
rect 6500 670 6550 680
rect 7350 670 7400 680
rect 8250 670 8400 680
rect 8650 670 8750 680
rect 9100 670 9150 680
rect 550 660 600 670
rect 700 660 900 670
rect 950 660 1050 670
rect 1250 660 1300 670
rect 3250 660 3300 670
rect 4750 660 4800 670
rect 5500 660 5700 670
rect 5750 660 6050 670
rect 6150 660 6300 670
rect 6500 660 6550 670
rect 7350 660 7400 670
rect 8250 660 8400 670
rect 8650 660 8750 670
rect 9100 660 9150 670
rect 550 650 600 660
rect 700 650 900 660
rect 950 650 1050 660
rect 1250 650 1300 660
rect 3250 650 3300 660
rect 4750 650 4800 660
rect 5500 650 5700 660
rect 5750 650 6050 660
rect 6150 650 6300 660
rect 6500 650 6550 660
rect 7350 650 7400 660
rect 8250 650 8400 660
rect 8650 650 8750 660
rect 9100 650 9150 660
rect 350 640 450 650
rect 800 640 900 650
rect 1200 640 1350 650
rect 2300 640 2350 650
rect 3100 640 3150 650
rect 4700 640 4800 650
rect 5550 640 5700 650
rect 5750 640 5950 650
rect 6250 640 6300 650
rect 6500 640 6550 650
rect 7350 640 7400 650
rect 8000 640 8050 650
rect 8300 640 8450 650
rect 8550 640 8750 650
rect 9100 640 9150 650
rect 350 630 450 640
rect 800 630 900 640
rect 1200 630 1350 640
rect 2300 630 2350 640
rect 3100 630 3150 640
rect 4700 630 4800 640
rect 5550 630 5700 640
rect 5750 630 5950 640
rect 6250 630 6300 640
rect 6500 630 6550 640
rect 7350 630 7400 640
rect 8000 630 8050 640
rect 8300 630 8450 640
rect 8550 630 8750 640
rect 9100 630 9150 640
rect 350 620 450 630
rect 800 620 900 630
rect 1200 620 1350 630
rect 2300 620 2350 630
rect 3100 620 3150 630
rect 4700 620 4800 630
rect 5550 620 5700 630
rect 5750 620 5950 630
rect 6250 620 6300 630
rect 6500 620 6550 630
rect 7350 620 7400 630
rect 8000 620 8050 630
rect 8300 620 8450 630
rect 8550 620 8750 630
rect 9100 620 9150 630
rect 350 610 450 620
rect 800 610 900 620
rect 1200 610 1350 620
rect 2300 610 2350 620
rect 3100 610 3150 620
rect 4700 610 4800 620
rect 5550 610 5700 620
rect 5750 610 5950 620
rect 6250 610 6300 620
rect 6500 610 6550 620
rect 7350 610 7400 620
rect 8000 610 8050 620
rect 8300 610 8450 620
rect 8550 610 8750 620
rect 9100 610 9150 620
rect 350 600 450 610
rect 800 600 900 610
rect 1200 600 1350 610
rect 2300 600 2350 610
rect 3100 600 3150 610
rect 4700 600 4800 610
rect 5550 600 5700 610
rect 5750 600 5950 610
rect 6250 600 6300 610
rect 6500 600 6550 610
rect 7350 600 7400 610
rect 8000 600 8050 610
rect 8300 600 8450 610
rect 8550 600 8750 610
rect 9100 600 9150 610
rect 300 590 350 600
rect 800 590 850 600
rect 1100 590 1250 600
rect 2100 590 2250 600
rect 3000 590 3050 600
rect 4700 590 4750 600
rect 4950 590 5000 600
rect 5600 590 5700 600
rect 5850 590 6000 600
rect 6250 590 6350 600
rect 6550 590 6600 600
rect 7350 590 7400 600
rect 8050 590 8150 600
rect 8350 590 8700 600
rect 9050 590 9150 600
rect 300 580 350 590
rect 800 580 850 590
rect 1100 580 1250 590
rect 2100 580 2250 590
rect 3000 580 3050 590
rect 4700 580 4750 590
rect 4950 580 5000 590
rect 5600 580 5700 590
rect 5850 580 6000 590
rect 6250 580 6350 590
rect 6550 580 6600 590
rect 7350 580 7400 590
rect 8050 580 8150 590
rect 8350 580 8700 590
rect 9050 580 9150 590
rect 300 570 350 580
rect 800 570 850 580
rect 1100 570 1250 580
rect 2100 570 2250 580
rect 3000 570 3050 580
rect 4700 570 4750 580
rect 4950 570 5000 580
rect 5600 570 5700 580
rect 5850 570 6000 580
rect 6250 570 6350 580
rect 6550 570 6600 580
rect 7350 570 7400 580
rect 8050 570 8150 580
rect 8350 570 8700 580
rect 9050 570 9150 580
rect 300 560 350 570
rect 800 560 850 570
rect 1100 560 1250 570
rect 2100 560 2250 570
rect 3000 560 3050 570
rect 4700 560 4750 570
rect 4950 560 5000 570
rect 5600 560 5700 570
rect 5850 560 6000 570
rect 6250 560 6350 570
rect 6550 560 6600 570
rect 7350 560 7400 570
rect 8050 560 8150 570
rect 8350 560 8700 570
rect 9050 560 9150 570
rect 300 550 350 560
rect 800 550 850 560
rect 1100 550 1250 560
rect 2100 550 2250 560
rect 3000 550 3050 560
rect 4700 550 4750 560
rect 4950 550 5000 560
rect 5600 550 5700 560
rect 5850 550 6000 560
rect 6250 550 6350 560
rect 6550 550 6600 560
rect 7350 550 7400 560
rect 8050 550 8150 560
rect 8350 550 8700 560
rect 9050 550 9150 560
rect 150 540 300 550
rect 650 540 900 550
rect 1050 540 1200 550
rect 1500 540 1550 550
rect 2850 540 2950 550
rect 4450 540 4550 550
rect 4650 540 4750 550
rect 4950 540 5000 550
rect 5850 540 6050 550
rect 6250 540 6350 550
rect 6600 540 6650 550
rect 7350 540 7400 550
rect 8450 540 8550 550
rect 9050 540 9150 550
rect 150 530 300 540
rect 650 530 900 540
rect 1050 530 1200 540
rect 1500 530 1550 540
rect 2850 530 2950 540
rect 4450 530 4550 540
rect 4650 530 4750 540
rect 4950 530 5000 540
rect 5850 530 6050 540
rect 6250 530 6350 540
rect 6600 530 6650 540
rect 7350 530 7400 540
rect 8450 530 8550 540
rect 9050 530 9150 540
rect 150 520 300 530
rect 650 520 900 530
rect 1050 520 1200 530
rect 1500 520 1550 530
rect 2850 520 2950 530
rect 4450 520 4550 530
rect 4650 520 4750 530
rect 4950 520 5000 530
rect 5850 520 6050 530
rect 6250 520 6350 530
rect 6600 520 6650 530
rect 7350 520 7400 530
rect 8450 520 8550 530
rect 9050 520 9150 530
rect 150 510 300 520
rect 650 510 900 520
rect 1050 510 1200 520
rect 1500 510 1550 520
rect 2850 510 2950 520
rect 4450 510 4550 520
rect 4650 510 4750 520
rect 4950 510 5000 520
rect 5850 510 6050 520
rect 6250 510 6350 520
rect 6600 510 6650 520
rect 7350 510 7400 520
rect 8450 510 8550 520
rect 9050 510 9150 520
rect 150 500 300 510
rect 650 500 900 510
rect 1050 500 1200 510
rect 1500 500 1550 510
rect 2850 500 2950 510
rect 4450 500 4550 510
rect 4650 500 4750 510
rect 4950 500 5000 510
rect 5850 500 6050 510
rect 6250 500 6350 510
rect 6600 500 6650 510
rect 7350 500 7400 510
rect 8450 500 8550 510
rect 9050 500 9150 510
rect 100 490 150 500
rect 550 490 650 500
rect 900 490 1150 500
rect 2000 490 2100 500
rect 2200 490 2250 500
rect 2700 490 2750 500
rect 4250 490 4350 500
rect 4550 490 4750 500
rect 5800 490 6050 500
rect 6200 490 6300 500
rect 6600 490 6650 500
rect 7300 490 7400 500
rect 9000 490 9100 500
rect 100 480 150 490
rect 550 480 650 490
rect 900 480 1150 490
rect 2000 480 2100 490
rect 2200 480 2250 490
rect 2700 480 2750 490
rect 4250 480 4350 490
rect 4550 480 4750 490
rect 5800 480 6050 490
rect 6200 480 6300 490
rect 6600 480 6650 490
rect 7300 480 7400 490
rect 9000 480 9100 490
rect 100 470 150 480
rect 550 470 650 480
rect 900 470 1150 480
rect 2000 470 2100 480
rect 2200 470 2250 480
rect 2700 470 2750 480
rect 4250 470 4350 480
rect 4550 470 4750 480
rect 5800 470 6050 480
rect 6200 470 6300 480
rect 6600 470 6650 480
rect 7300 470 7400 480
rect 9000 470 9100 480
rect 100 460 150 470
rect 550 460 650 470
rect 900 460 1150 470
rect 2000 460 2100 470
rect 2200 460 2250 470
rect 2700 460 2750 470
rect 4250 460 4350 470
rect 4550 460 4750 470
rect 5800 460 6050 470
rect 6200 460 6300 470
rect 6600 460 6650 470
rect 7300 460 7400 470
rect 9000 460 9100 470
rect 100 450 150 460
rect 550 450 650 460
rect 900 450 1150 460
rect 2000 450 2100 460
rect 2200 450 2250 460
rect 2700 450 2750 460
rect 4250 450 4350 460
rect 4550 450 4750 460
rect 5800 450 6050 460
rect 6200 450 6300 460
rect 6600 450 6650 460
rect 7300 450 7400 460
rect 9000 450 9100 460
rect 50 440 100 450
rect 500 440 700 450
rect 1000 440 1100 450
rect 4250 440 4300 450
rect 4550 440 4650 450
rect 4700 440 4750 450
rect 5800 440 5900 450
rect 5950 440 6050 450
rect 6200 440 6300 450
rect 6650 440 6700 450
rect 7300 440 7350 450
rect 8950 440 9100 450
rect 50 430 100 440
rect 500 430 700 440
rect 1000 430 1100 440
rect 4250 430 4300 440
rect 4550 430 4650 440
rect 4700 430 4750 440
rect 5800 430 5900 440
rect 5950 430 6050 440
rect 6200 430 6300 440
rect 6650 430 6700 440
rect 7300 430 7350 440
rect 8950 430 9100 440
rect 50 420 100 430
rect 500 420 700 430
rect 1000 420 1100 430
rect 4250 420 4300 430
rect 4550 420 4650 430
rect 4700 420 4750 430
rect 5800 420 5900 430
rect 5950 420 6050 430
rect 6200 420 6300 430
rect 6650 420 6700 430
rect 7300 420 7350 430
rect 8950 420 9100 430
rect 50 410 100 420
rect 500 410 700 420
rect 1000 410 1100 420
rect 4250 410 4300 420
rect 4550 410 4650 420
rect 4700 410 4750 420
rect 5800 410 5900 420
rect 5950 410 6050 420
rect 6200 410 6300 420
rect 6650 410 6700 420
rect 7300 410 7350 420
rect 8950 410 9100 420
rect 50 400 100 410
rect 500 400 700 410
rect 1000 400 1100 410
rect 4250 400 4300 410
rect 4550 400 4650 410
rect 4700 400 4750 410
rect 5800 400 5900 410
rect 5950 400 6050 410
rect 6200 400 6300 410
rect 6650 400 6700 410
rect 7300 400 7350 410
rect 8950 400 9100 410
rect 0 390 50 400
rect 400 390 450 400
rect 500 390 700 400
rect 4250 390 4300 400
rect 4350 390 4400 400
rect 4550 390 4600 400
rect 5800 390 5850 400
rect 5950 390 6050 400
rect 6200 390 6300 400
rect 6700 390 6750 400
rect 7300 390 7350 400
rect 8800 390 8850 400
rect 8950 390 9100 400
rect 0 380 50 390
rect 400 380 450 390
rect 500 380 700 390
rect 4250 380 4300 390
rect 4350 380 4400 390
rect 4550 380 4600 390
rect 5800 380 5850 390
rect 5950 380 6050 390
rect 6200 380 6300 390
rect 6700 380 6750 390
rect 7300 380 7350 390
rect 8800 380 8850 390
rect 8950 380 9100 390
rect 0 370 50 380
rect 400 370 450 380
rect 500 370 700 380
rect 4250 370 4300 380
rect 4350 370 4400 380
rect 4550 370 4600 380
rect 5800 370 5850 380
rect 5950 370 6050 380
rect 6200 370 6300 380
rect 6700 370 6750 380
rect 7300 370 7350 380
rect 8800 370 8850 380
rect 8950 370 9100 380
rect 0 360 50 370
rect 400 360 450 370
rect 500 360 700 370
rect 4250 360 4300 370
rect 4350 360 4400 370
rect 4550 360 4600 370
rect 5800 360 5850 370
rect 5950 360 6050 370
rect 6200 360 6300 370
rect 6700 360 6750 370
rect 7300 360 7350 370
rect 8800 360 8850 370
rect 8950 360 9100 370
rect 0 350 50 360
rect 400 350 450 360
rect 500 350 700 360
rect 4250 350 4300 360
rect 4350 350 4400 360
rect 4550 350 4600 360
rect 5800 350 5850 360
rect 5950 350 6050 360
rect 6200 350 6300 360
rect 6700 350 6750 360
rect 7300 350 7350 360
rect 8800 350 8850 360
rect 8950 350 9100 360
rect 400 340 450 350
rect 700 340 800 350
rect 1000 340 1050 350
rect 4450 340 4600 350
rect 4650 340 4700 350
rect 6000 340 6150 350
rect 6200 340 6300 350
rect 6700 340 6750 350
rect 7250 340 7350 350
rect 8800 340 8850 350
rect 9000 340 9050 350
rect 9250 340 9400 350
rect 400 330 450 340
rect 700 330 800 340
rect 1000 330 1050 340
rect 4450 330 4600 340
rect 4650 330 4700 340
rect 6000 330 6150 340
rect 6200 330 6300 340
rect 6700 330 6750 340
rect 7250 330 7350 340
rect 8800 330 8850 340
rect 9000 330 9050 340
rect 9250 330 9400 340
rect 400 320 450 330
rect 700 320 800 330
rect 1000 320 1050 330
rect 4450 320 4600 330
rect 4650 320 4700 330
rect 6000 320 6150 330
rect 6200 320 6300 330
rect 6700 320 6750 330
rect 7250 320 7350 330
rect 8800 320 8850 330
rect 9000 320 9050 330
rect 9250 320 9400 330
rect 400 310 450 320
rect 700 310 800 320
rect 1000 310 1050 320
rect 4450 310 4600 320
rect 4650 310 4700 320
rect 6000 310 6150 320
rect 6200 310 6300 320
rect 6700 310 6750 320
rect 7250 310 7350 320
rect 8800 310 8850 320
rect 9000 310 9050 320
rect 9250 310 9400 320
rect 400 300 450 310
rect 700 300 800 310
rect 1000 300 1050 310
rect 4450 300 4600 310
rect 4650 300 4700 310
rect 6000 300 6150 310
rect 6200 300 6300 310
rect 6700 300 6750 310
rect 7250 300 7350 310
rect 8800 300 8850 310
rect 9000 300 9050 310
rect 9250 300 9400 310
rect 900 290 1000 300
rect 4550 290 4650 300
rect 6000 290 6300 300
rect 6750 290 6850 300
rect 7250 290 7350 300
rect 8850 290 8950 300
rect 9000 290 9050 300
rect 9250 290 9400 300
rect 900 280 1000 290
rect 4550 280 4650 290
rect 6000 280 6300 290
rect 6750 280 6850 290
rect 7250 280 7350 290
rect 8850 280 8950 290
rect 9000 280 9050 290
rect 9250 280 9400 290
rect 900 270 1000 280
rect 4550 270 4650 280
rect 6000 270 6300 280
rect 6750 270 6850 280
rect 7250 270 7350 280
rect 8850 270 8950 280
rect 9000 270 9050 280
rect 9250 270 9400 280
rect 900 260 1000 270
rect 4550 260 4650 270
rect 6000 260 6300 270
rect 6750 260 6850 270
rect 7250 260 7350 270
rect 8850 260 8950 270
rect 9000 260 9050 270
rect 9250 260 9400 270
rect 900 250 1000 260
rect 4550 250 4650 260
rect 6000 250 6300 260
rect 6750 250 6850 260
rect 7250 250 7350 260
rect 8850 250 8950 260
rect 9000 250 9050 260
rect 9250 250 9400 260
rect 150 240 200 250
rect 5000 240 5050 250
rect 6100 240 6300 250
rect 6800 240 6950 250
rect 7250 240 7350 250
rect 8950 240 9000 250
rect 9200 240 9250 250
rect 150 230 200 240
rect 5000 230 5050 240
rect 6100 230 6300 240
rect 6800 230 6950 240
rect 7250 230 7350 240
rect 8950 230 9000 240
rect 9200 230 9250 240
rect 150 220 200 230
rect 5000 220 5050 230
rect 6100 220 6300 230
rect 6800 220 6950 230
rect 7250 220 7350 230
rect 8950 220 9000 230
rect 9200 220 9250 230
rect 150 210 200 220
rect 5000 210 5050 220
rect 6100 210 6300 220
rect 6800 210 6950 220
rect 7250 210 7350 220
rect 8950 210 9000 220
rect 9200 210 9250 220
rect 150 200 200 210
rect 5000 200 5050 210
rect 6100 200 6300 210
rect 6800 200 6950 210
rect 7250 200 7350 210
rect 8950 200 9000 210
rect 9200 200 9250 210
rect 100 190 150 200
rect 350 190 450 200
rect 5000 190 5050 200
rect 6050 190 6150 200
rect 6250 190 6350 200
rect 6900 190 7050 200
rect 7250 190 7350 200
rect 8550 190 8750 200
rect 8800 190 8850 200
rect 8900 190 9000 200
rect 9200 190 9300 200
rect 9800 190 9850 200
rect 100 180 150 190
rect 350 180 450 190
rect 5000 180 5050 190
rect 6050 180 6150 190
rect 6250 180 6350 190
rect 6900 180 7050 190
rect 7250 180 7350 190
rect 8550 180 8750 190
rect 8800 180 8850 190
rect 8900 180 9000 190
rect 9200 180 9300 190
rect 9800 180 9850 190
rect 100 170 150 180
rect 350 170 450 180
rect 5000 170 5050 180
rect 6050 170 6150 180
rect 6250 170 6350 180
rect 6900 170 7050 180
rect 7250 170 7350 180
rect 8550 170 8750 180
rect 8800 170 8850 180
rect 8900 170 9000 180
rect 9200 170 9300 180
rect 9800 170 9850 180
rect 100 160 150 170
rect 350 160 450 170
rect 5000 160 5050 170
rect 6050 160 6150 170
rect 6250 160 6350 170
rect 6900 160 7050 170
rect 7250 160 7350 170
rect 8550 160 8750 170
rect 8800 160 8850 170
rect 8900 160 9000 170
rect 9200 160 9300 170
rect 9800 160 9850 170
rect 100 150 150 160
rect 350 150 450 160
rect 5000 150 5050 160
rect 6050 150 6150 160
rect 6250 150 6350 160
rect 6900 150 7050 160
rect 7250 150 7350 160
rect 8550 150 8750 160
rect 8800 150 8850 160
rect 8900 150 9000 160
rect 9200 150 9300 160
rect 9800 150 9850 160
rect 150 140 350 150
rect 500 140 700 150
rect 750 140 900 150
rect 4250 140 4500 150
rect 4850 140 4900 150
rect 5950 140 6150 150
rect 6250 140 6350 150
rect 7000 140 7100 150
rect 7250 140 7350 150
rect 8550 140 8800 150
rect 9050 140 9100 150
rect 9300 140 9350 150
rect 9750 140 9800 150
rect 9850 140 9900 150
rect 150 130 350 140
rect 500 130 700 140
rect 750 130 900 140
rect 4250 130 4500 140
rect 4850 130 4900 140
rect 5950 130 6150 140
rect 6250 130 6350 140
rect 7000 130 7100 140
rect 7250 130 7350 140
rect 8550 130 8800 140
rect 9050 130 9100 140
rect 9300 130 9350 140
rect 9750 130 9800 140
rect 9850 130 9900 140
rect 150 120 350 130
rect 500 120 700 130
rect 750 120 900 130
rect 4250 120 4500 130
rect 4850 120 4900 130
rect 5950 120 6150 130
rect 6250 120 6350 130
rect 7000 120 7100 130
rect 7250 120 7350 130
rect 8550 120 8800 130
rect 9050 120 9100 130
rect 9300 120 9350 130
rect 9750 120 9800 130
rect 9850 120 9900 130
rect 150 110 350 120
rect 500 110 700 120
rect 750 110 900 120
rect 4250 110 4500 120
rect 4850 110 4900 120
rect 5950 110 6150 120
rect 6250 110 6350 120
rect 7000 110 7100 120
rect 7250 110 7350 120
rect 8550 110 8800 120
rect 9050 110 9100 120
rect 9300 110 9350 120
rect 9750 110 9800 120
rect 9850 110 9900 120
rect 150 100 350 110
rect 500 100 700 110
rect 750 100 900 110
rect 4250 100 4500 110
rect 4850 100 4900 110
rect 5950 100 6150 110
rect 6250 100 6350 110
rect 7000 100 7100 110
rect 7250 100 7350 110
rect 8550 100 8800 110
rect 9050 100 9100 110
rect 9300 100 9350 110
rect 9750 100 9800 110
rect 9850 100 9900 110
rect 150 90 200 100
rect 250 90 350 100
rect 600 90 750 100
rect 800 90 950 100
rect 4300 90 4350 100
rect 4450 90 4600 100
rect 4800 90 4900 100
rect 5850 90 6000 100
rect 6050 90 6150 100
rect 6300 90 6400 100
rect 7050 90 7200 100
rect 7250 90 7350 100
rect 8600 90 8750 100
rect 8950 90 9000 100
rect 9350 90 9400 100
rect 9750 90 9800 100
rect 9850 90 9900 100
rect 150 80 200 90
rect 250 80 350 90
rect 600 80 750 90
rect 800 80 950 90
rect 4300 80 4350 90
rect 4450 80 4600 90
rect 4800 80 4900 90
rect 5850 80 6000 90
rect 6050 80 6150 90
rect 6300 80 6400 90
rect 7050 80 7200 90
rect 7250 80 7350 90
rect 8600 80 8750 90
rect 8950 80 9000 90
rect 9350 80 9400 90
rect 9750 80 9800 90
rect 9850 80 9900 90
rect 150 70 200 80
rect 250 70 350 80
rect 600 70 750 80
rect 800 70 950 80
rect 4300 70 4350 80
rect 4450 70 4600 80
rect 4800 70 4900 80
rect 5850 70 6000 80
rect 6050 70 6150 80
rect 6300 70 6400 80
rect 7050 70 7200 80
rect 7250 70 7350 80
rect 8600 70 8750 80
rect 8950 70 9000 80
rect 9350 70 9400 80
rect 9750 70 9800 80
rect 9850 70 9900 80
rect 150 60 200 70
rect 250 60 350 70
rect 600 60 750 70
rect 800 60 950 70
rect 4300 60 4350 70
rect 4450 60 4600 70
rect 4800 60 4900 70
rect 5850 60 6000 70
rect 6050 60 6150 70
rect 6300 60 6400 70
rect 7050 60 7200 70
rect 7250 60 7350 70
rect 8600 60 8750 70
rect 8950 60 9000 70
rect 9350 60 9400 70
rect 9750 60 9800 70
rect 9850 60 9900 70
rect 150 50 200 60
rect 250 50 350 60
rect 600 50 750 60
rect 800 50 950 60
rect 4300 50 4350 60
rect 4450 50 4600 60
rect 4800 50 4900 60
rect 5850 50 6000 60
rect 6050 50 6150 60
rect 6300 50 6400 60
rect 7050 50 7200 60
rect 7250 50 7350 60
rect 8600 50 8750 60
rect 8950 50 9000 60
rect 9350 50 9400 60
rect 9750 50 9800 60
rect 9850 50 9900 60
rect 150 40 200 50
rect 650 40 750 50
rect 850 40 950 50
rect 4550 40 4650 50
rect 4750 40 4900 50
rect 5050 40 5100 50
rect 6050 40 6150 50
rect 6350 40 6450 50
rect 7100 40 7200 50
rect 7250 40 7350 50
rect 8550 40 8600 50
rect 8650 40 8700 50
rect 150 30 200 40
rect 650 30 750 40
rect 850 30 950 40
rect 4550 30 4650 40
rect 4750 30 4900 40
rect 5050 30 5100 40
rect 6050 30 6150 40
rect 6350 30 6450 40
rect 7100 30 7200 40
rect 7250 30 7350 40
rect 8550 30 8600 40
rect 8650 30 8700 40
rect 150 20 200 30
rect 650 20 750 30
rect 850 20 950 30
rect 4550 20 4650 30
rect 4750 20 4900 30
rect 5050 20 5100 30
rect 6050 20 6150 30
rect 6350 20 6450 30
rect 7100 20 7200 30
rect 7250 20 7350 30
rect 8550 20 8600 30
rect 8650 20 8700 30
rect 150 10 200 20
rect 650 10 750 20
rect 850 10 950 20
rect 4550 10 4650 20
rect 4750 10 4900 20
rect 5050 10 5100 20
rect 6050 10 6150 20
rect 6350 10 6450 20
rect 7100 10 7200 20
rect 7250 10 7350 20
rect 8550 10 8600 20
rect 8650 10 8700 20
rect 150 0 200 10
rect 650 0 750 10
rect 850 0 950 10
rect 4550 0 4650 10
rect 4750 0 4900 10
rect 5050 0 5100 10
rect 6050 0 6150 10
rect 6350 0 6450 10
rect 7100 0 7200 10
rect 7250 0 7350 10
rect 8550 0 8600 10
rect 8650 0 8700 10
<< metal3 >>
rect 2150 7490 2200 7500
rect 3300 7490 3350 7500
rect 3550 7490 3600 7500
rect 3650 7490 3700 7500
rect 9650 7490 9800 7500
rect 2150 7480 2200 7490
rect 3300 7480 3350 7490
rect 3550 7480 3600 7490
rect 3650 7480 3700 7490
rect 9650 7480 9800 7490
rect 2150 7470 2200 7480
rect 3300 7470 3350 7480
rect 3550 7470 3600 7480
rect 3650 7470 3700 7480
rect 9650 7470 9800 7480
rect 2150 7460 2200 7470
rect 3300 7460 3350 7470
rect 3550 7460 3600 7470
rect 3650 7460 3700 7470
rect 9650 7460 9800 7470
rect 2150 7450 2200 7460
rect 3300 7450 3350 7460
rect 3550 7450 3600 7460
rect 3650 7450 3700 7460
rect 9650 7450 9800 7460
rect 2100 7440 2150 7450
rect 3300 7440 3350 7450
rect 9600 7440 9650 7450
rect 2100 7430 2150 7440
rect 3300 7430 3350 7440
rect 9600 7430 9650 7440
rect 2100 7420 2150 7430
rect 3300 7420 3350 7430
rect 9600 7420 9650 7430
rect 2100 7410 2150 7420
rect 3300 7410 3350 7420
rect 9600 7410 9650 7420
rect 2100 7400 2150 7410
rect 3300 7400 3350 7410
rect 9600 7400 9650 7410
rect 2050 7390 2100 7400
rect 9600 7390 9650 7400
rect 2050 7380 2100 7390
rect 9600 7380 9650 7390
rect 2050 7370 2100 7380
rect 9600 7370 9650 7380
rect 2050 7360 2100 7370
rect 9600 7360 9650 7370
rect 2050 7350 2100 7360
rect 9600 7350 9650 7360
rect 9600 7340 9650 7350
rect 9850 7340 9900 7350
rect 9600 7330 9650 7340
rect 9850 7330 9900 7340
rect 9600 7320 9650 7330
rect 9850 7320 9900 7330
rect 9600 7310 9650 7320
rect 9850 7310 9900 7320
rect 9600 7300 9650 7310
rect 9850 7300 9900 7310
rect 3350 7290 3400 7300
rect 9600 7290 9650 7300
rect 9800 7290 9900 7300
rect 3350 7280 3400 7290
rect 9600 7280 9650 7290
rect 9800 7280 9900 7290
rect 3350 7270 3400 7280
rect 9600 7270 9650 7280
rect 9800 7270 9900 7280
rect 3350 7260 3400 7270
rect 9600 7260 9650 7270
rect 9800 7260 9900 7270
rect 3350 7250 3400 7260
rect 9600 7250 9650 7260
rect 9800 7250 9900 7260
rect 1950 7240 2000 7250
rect 3400 7240 3450 7250
rect 3850 7240 3900 7250
rect 9600 7240 9800 7250
rect 1950 7230 2000 7240
rect 3400 7230 3450 7240
rect 3850 7230 3900 7240
rect 9600 7230 9800 7240
rect 1950 7220 2000 7230
rect 3400 7220 3450 7230
rect 3850 7220 3900 7230
rect 9600 7220 9800 7230
rect 1950 7210 2000 7220
rect 3400 7210 3450 7220
rect 3850 7210 3900 7220
rect 9600 7210 9800 7220
rect 1950 7200 2000 7210
rect 3400 7200 3450 7210
rect 3850 7200 3900 7210
rect 9600 7200 9800 7210
rect 3350 7190 3400 7200
rect 3800 7190 3850 7200
rect 9600 7190 9650 7200
rect 3350 7180 3400 7190
rect 3800 7180 3850 7190
rect 9600 7180 9650 7190
rect 3350 7170 3400 7180
rect 3800 7170 3850 7180
rect 9600 7170 9650 7180
rect 3350 7160 3400 7170
rect 3800 7160 3850 7170
rect 9600 7160 9650 7170
rect 3350 7150 3400 7160
rect 3800 7150 3850 7160
rect 9600 7150 9650 7160
rect 1900 7140 1950 7150
rect 3400 7140 3450 7150
rect 3650 7140 3700 7150
rect 3800 7140 3850 7150
rect 3900 7140 3950 7150
rect 9600 7140 9650 7150
rect 1900 7130 1950 7140
rect 3400 7130 3450 7140
rect 3650 7130 3700 7140
rect 3800 7130 3850 7140
rect 3900 7130 3950 7140
rect 9600 7130 9650 7140
rect 1900 7120 1950 7130
rect 3400 7120 3450 7130
rect 3650 7120 3700 7130
rect 3800 7120 3850 7130
rect 3900 7120 3950 7130
rect 9600 7120 9650 7130
rect 1900 7110 1950 7120
rect 3400 7110 3450 7120
rect 3650 7110 3700 7120
rect 3800 7110 3850 7120
rect 3900 7110 3950 7120
rect 9600 7110 9650 7120
rect 1900 7100 1950 7110
rect 3400 7100 3450 7110
rect 3650 7100 3700 7110
rect 3800 7100 3850 7110
rect 3900 7100 3950 7110
rect 9600 7100 9650 7110
rect 1900 7090 1950 7100
rect 3500 7090 3550 7100
rect 3700 7090 3850 7100
rect 3900 7090 3950 7100
rect 1900 7080 1950 7090
rect 3500 7080 3550 7090
rect 3700 7080 3850 7090
rect 3900 7080 3950 7090
rect 1900 7070 1950 7080
rect 3500 7070 3550 7080
rect 3700 7070 3850 7080
rect 3900 7070 3950 7080
rect 1900 7060 1950 7070
rect 3500 7060 3550 7070
rect 3700 7060 3850 7070
rect 3900 7060 3950 7070
rect 1900 7050 1950 7060
rect 3500 7050 3550 7060
rect 3700 7050 3850 7060
rect 3900 7050 3950 7060
rect 1900 7040 1950 7050
rect 3700 7040 3750 7050
rect 3800 7040 3950 7050
rect 9600 7040 9650 7050
rect 1900 7030 1950 7040
rect 3700 7030 3750 7040
rect 3800 7030 3950 7040
rect 9600 7030 9650 7040
rect 1900 7020 1950 7030
rect 3700 7020 3750 7030
rect 3800 7020 3950 7030
rect 9600 7020 9650 7030
rect 1900 7010 1950 7020
rect 3700 7010 3750 7020
rect 3800 7010 3950 7020
rect 9600 7010 9650 7020
rect 1900 7000 1950 7010
rect 3700 7000 3750 7010
rect 3800 7000 3950 7010
rect 9600 7000 9650 7010
rect 3150 6990 3300 7000
rect 3600 6990 3700 7000
rect 3850 6990 3950 7000
rect 9600 6990 9650 7000
rect 3150 6980 3300 6990
rect 3600 6980 3700 6990
rect 3850 6980 3950 6990
rect 9600 6980 9650 6990
rect 3150 6970 3300 6980
rect 3600 6970 3700 6980
rect 3850 6970 3950 6980
rect 9600 6970 9650 6980
rect 3150 6960 3300 6970
rect 3600 6960 3700 6970
rect 3850 6960 3950 6970
rect 9600 6960 9650 6970
rect 3150 6950 3300 6960
rect 3600 6950 3700 6960
rect 3850 6950 3950 6960
rect 9600 6950 9650 6960
rect 1900 6940 1950 6950
rect 2400 6940 2650 6950
rect 2750 6940 3250 6950
rect 3400 6940 3450 6950
rect 3750 6940 3900 6950
rect 9600 6940 9650 6950
rect 1900 6930 1950 6940
rect 2400 6930 2650 6940
rect 2750 6930 3250 6940
rect 3400 6930 3450 6940
rect 3750 6930 3900 6940
rect 9600 6930 9650 6940
rect 1900 6920 1950 6930
rect 2400 6920 2650 6930
rect 2750 6920 3250 6930
rect 3400 6920 3450 6930
rect 3750 6920 3900 6930
rect 9600 6920 9650 6930
rect 1900 6910 1950 6920
rect 2400 6910 2650 6920
rect 2750 6910 3250 6920
rect 3400 6910 3450 6920
rect 3750 6910 3900 6920
rect 9600 6910 9650 6920
rect 1900 6900 1950 6910
rect 2400 6900 2650 6910
rect 2750 6900 3250 6910
rect 3400 6900 3450 6910
rect 3750 6900 3900 6910
rect 9600 6900 9650 6910
rect 2500 6890 3250 6900
rect 3500 6890 3550 6900
rect 3800 6890 3900 6900
rect 9600 6890 9650 6900
rect 2500 6880 3250 6890
rect 3500 6880 3550 6890
rect 3800 6880 3900 6890
rect 9600 6880 9650 6890
rect 2500 6870 3250 6880
rect 3500 6870 3550 6880
rect 3800 6870 3900 6880
rect 9600 6870 9650 6880
rect 2500 6860 3250 6870
rect 3500 6860 3550 6870
rect 3800 6860 3900 6870
rect 9600 6860 9650 6870
rect 2500 6850 3250 6860
rect 3500 6850 3550 6860
rect 3800 6850 3900 6860
rect 9600 6850 9650 6860
rect 2550 6840 3100 6850
rect 3600 6840 3650 6850
rect 3850 6840 3900 6850
rect 9600 6840 9650 6850
rect 2550 6830 3100 6840
rect 3600 6830 3650 6840
rect 3850 6830 3900 6840
rect 9600 6830 9650 6840
rect 2550 6820 3100 6830
rect 3600 6820 3650 6830
rect 3850 6820 3900 6830
rect 9600 6820 9650 6830
rect 2550 6810 3100 6820
rect 3600 6810 3650 6820
rect 3850 6810 3900 6820
rect 9600 6810 9650 6820
rect 2550 6800 3100 6810
rect 3600 6800 3650 6810
rect 3850 6800 3900 6810
rect 9600 6800 9650 6810
rect 1850 6790 1900 6800
rect 2800 6790 3050 6800
rect 3900 6790 3950 6800
rect 1850 6780 1900 6790
rect 2800 6780 3050 6790
rect 3900 6780 3950 6790
rect 1850 6770 1900 6780
rect 2800 6770 3050 6780
rect 3900 6770 3950 6780
rect 1850 6760 1900 6770
rect 2800 6760 3050 6770
rect 3900 6760 3950 6770
rect 1850 6750 1900 6760
rect 2800 6750 3050 6760
rect 3900 6750 3950 6760
rect 1850 6740 1900 6750
rect 2250 6740 2350 6750
rect 2450 6740 2500 6750
rect 3200 6740 3300 6750
rect 3750 6740 3800 6750
rect 3900 6740 3950 6750
rect 9550 6740 9600 6750
rect 1850 6730 1900 6740
rect 2250 6730 2350 6740
rect 2450 6730 2500 6740
rect 3200 6730 3300 6740
rect 3750 6730 3800 6740
rect 3900 6730 3950 6740
rect 9550 6730 9600 6740
rect 1850 6720 1900 6730
rect 2250 6720 2350 6730
rect 2450 6720 2500 6730
rect 3200 6720 3300 6730
rect 3750 6720 3800 6730
rect 3900 6720 3950 6730
rect 9550 6720 9600 6730
rect 1850 6710 1900 6720
rect 2250 6710 2350 6720
rect 2450 6710 2500 6720
rect 3200 6710 3300 6720
rect 3750 6710 3800 6720
rect 3900 6710 3950 6720
rect 9550 6710 9600 6720
rect 1850 6700 1900 6710
rect 2250 6700 2350 6710
rect 2450 6700 2500 6710
rect 3200 6700 3300 6710
rect 3750 6700 3800 6710
rect 3900 6700 3950 6710
rect 9550 6700 9600 6710
rect 1850 6690 1900 6700
rect 2500 6690 2550 6700
rect 3450 6690 3500 6700
rect 3800 6690 3850 6700
rect 9500 6690 9550 6700
rect 9600 6690 9650 6700
rect 9900 6690 9950 6700
rect 1850 6680 1900 6690
rect 2500 6680 2550 6690
rect 3450 6680 3500 6690
rect 3800 6680 3850 6690
rect 9500 6680 9550 6690
rect 9600 6680 9650 6690
rect 9900 6680 9950 6690
rect 1850 6670 1900 6680
rect 2500 6670 2550 6680
rect 3450 6670 3500 6680
rect 3800 6670 3850 6680
rect 9500 6670 9550 6680
rect 9600 6670 9650 6680
rect 9900 6670 9950 6680
rect 1850 6660 1900 6670
rect 2500 6660 2550 6670
rect 3450 6660 3500 6670
rect 3800 6660 3850 6670
rect 9500 6660 9550 6670
rect 9600 6660 9650 6670
rect 9900 6660 9950 6670
rect 1850 6650 1900 6660
rect 2500 6650 2550 6660
rect 3450 6650 3500 6660
rect 3800 6650 3850 6660
rect 9500 6650 9550 6660
rect 9600 6650 9650 6660
rect 9900 6650 9950 6660
rect 1750 6640 1800 6650
rect 2200 6640 2250 6650
rect 2550 6640 2600 6650
rect 3600 6640 3650 6650
rect 3850 6640 3900 6650
rect 9500 6640 9550 6650
rect 9600 6640 9650 6650
rect 9750 6640 9800 6650
rect 1750 6630 1800 6640
rect 2200 6630 2250 6640
rect 2550 6630 2600 6640
rect 3600 6630 3650 6640
rect 3850 6630 3900 6640
rect 9500 6630 9550 6640
rect 9600 6630 9650 6640
rect 9750 6630 9800 6640
rect 1750 6620 1800 6630
rect 2200 6620 2250 6630
rect 2550 6620 2600 6630
rect 3600 6620 3650 6630
rect 3850 6620 3900 6630
rect 9500 6620 9550 6630
rect 9600 6620 9650 6630
rect 9750 6620 9800 6630
rect 1750 6610 1800 6620
rect 2200 6610 2250 6620
rect 2550 6610 2600 6620
rect 3600 6610 3650 6620
rect 3850 6610 3900 6620
rect 9500 6610 9550 6620
rect 9600 6610 9650 6620
rect 9750 6610 9800 6620
rect 1750 6600 1800 6610
rect 2200 6600 2250 6610
rect 2550 6600 2600 6610
rect 3600 6600 3650 6610
rect 3850 6600 3900 6610
rect 9500 6600 9550 6610
rect 9600 6600 9650 6610
rect 9750 6600 9800 6610
rect 1550 6590 1650 6600
rect 1750 6590 1800 6600
rect 2050 6590 2150 6600
rect 3700 6590 3750 6600
rect 3900 6590 4000 6600
rect 1550 6580 1650 6590
rect 1750 6580 1800 6590
rect 2050 6580 2150 6590
rect 3700 6580 3750 6590
rect 3900 6580 4000 6590
rect 1550 6570 1650 6580
rect 1750 6570 1800 6580
rect 2050 6570 2150 6580
rect 3700 6570 3750 6580
rect 3900 6570 4000 6580
rect 1550 6560 1650 6570
rect 1750 6560 1800 6570
rect 2050 6560 2150 6570
rect 3700 6560 3750 6570
rect 3900 6560 4000 6570
rect 1550 6550 1650 6560
rect 1750 6550 1800 6560
rect 2050 6550 2150 6560
rect 3700 6550 3750 6560
rect 3900 6550 4000 6560
rect 1350 6540 1450 6550
rect 1750 6540 1800 6550
rect 2050 6540 2100 6550
rect 2550 6540 2600 6550
rect 3800 6540 3850 6550
rect 3950 6540 4000 6550
rect 6150 6540 6600 6550
rect 1350 6530 1450 6540
rect 1750 6530 1800 6540
rect 2050 6530 2100 6540
rect 2550 6530 2600 6540
rect 3800 6530 3850 6540
rect 3950 6530 4000 6540
rect 6150 6530 6600 6540
rect 1350 6520 1450 6530
rect 1750 6520 1800 6530
rect 2050 6520 2100 6530
rect 2550 6520 2600 6530
rect 3800 6520 3850 6530
rect 3950 6520 4000 6530
rect 6150 6520 6600 6530
rect 1350 6510 1450 6520
rect 1750 6510 1800 6520
rect 2050 6510 2100 6520
rect 2550 6510 2600 6520
rect 3800 6510 3850 6520
rect 3950 6510 4000 6520
rect 6150 6510 6600 6520
rect 1350 6500 1450 6510
rect 1750 6500 1800 6510
rect 2050 6500 2100 6510
rect 2550 6500 2600 6510
rect 3800 6500 3850 6510
rect 3950 6500 4000 6510
rect 6150 6500 6600 6510
rect 1250 6490 1300 6500
rect 2100 6490 2150 6500
rect 6050 6490 6150 6500
rect 6200 6490 6350 6500
rect 6550 6490 6650 6500
rect 9800 6490 9900 6500
rect 1250 6480 1300 6490
rect 2100 6480 2150 6490
rect 6050 6480 6150 6490
rect 6200 6480 6350 6490
rect 6550 6480 6650 6490
rect 9800 6480 9900 6490
rect 1250 6470 1300 6480
rect 2100 6470 2150 6480
rect 6050 6470 6150 6480
rect 6200 6470 6350 6480
rect 6550 6470 6650 6480
rect 9800 6470 9900 6480
rect 1250 6460 1300 6470
rect 2100 6460 2150 6470
rect 6050 6460 6150 6470
rect 6200 6460 6350 6470
rect 6550 6460 6650 6470
rect 9800 6460 9900 6470
rect 1250 6450 1300 6460
rect 2100 6450 2150 6460
rect 6050 6450 6150 6460
rect 6200 6450 6350 6460
rect 6550 6450 6650 6460
rect 9800 6450 9900 6460
rect 1250 6440 1350 6450
rect 1750 6440 1950 6450
rect 2050 6440 2100 6450
rect 3950 6440 4000 6450
rect 6050 6440 6100 6450
rect 6600 6440 6700 6450
rect 9650 6440 9700 6450
rect 1250 6430 1350 6440
rect 1750 6430 1950 6440
rect 2050 6430 2100 6440
rect 3950 6430 4000 6440
rect 6050 6430 6100 6440
rect 6600 6430 6700 6440
rect 9650 6430 9700 6440
rect 1250 6420 1350 6430
rect 1750 6420 1950 6430
rect 2050 6420 2100 6430
rect 3950 6420 4000 6430
rect 6050 6420 6100 6430
rect 6600 6420 6700 6430
rect 9650 6420 9700 6430
rect 1250 6410 1350 6420
rect 1750 6410 1950 6420
rect 2050 6410 2100 6420
rect 3950 6410 4000 6420
rect 6050 6410 6100 6420
rect 6600 6410 6700 6420
rect 9650 6410 9700 6420
rect 1250 6400 1350 6410
rect 1750 6400 1950 6410
rect 2050 6400 2100 6410
rect 3950 6400 4000 6410
rect 6050 6400 6100 6410
rect 6600 6400 6700 6410
rect 9650 6400 9700 6410
rect 1400 6390 1450 6400
rect 1600 6390 1650 6400
rect 1700 6390 1850 6400
rect 5800 6390 5850 6400
rect 6150 6390 6250 6400
rect 6350 6390 6400 6400
rect 6650 6390 6800 6400
rect 1400 6380 1450 6390
rect 1600 6380 1650 6390
rect 1700 6380 1850 6390
rect 5800 6380 5850 6390
rect 6150 6380 6250 6390
rect 6350 6380 6400 6390
rect 6650 6380 6800 6390
rect 1400 6370 1450 6380
rect 1600 6370 1650 6380
rect 1700 6370 1850 6380
rect 5800 6370 5850 6380
rect 6150 6370 6250 6380
rect 6350 6370 6400 6380
rect 6650 6370 6800 6380
rect 1400 6360 1450 6370
rect 1600 6360 1650 6370
rect 1700 6360 1850 6370
rect 5800 6360 5850 6370
rect 6150 6360 6250 6370
rect 6350 6360 6400 6370
rect 6650 6360 6800 6370
rect 1400 6350 1450 6360
rect 1600 6350 1650 6360
rect 1700 6350 1850 6360
rect 5800 6350 5850 6360
rect 6150 6350 6250 6360
rect 6350 6350 6400 6360
rect 6650 6350 6800 6360
rect 1400 6340 1450 6350
rect 1600 6340 1700 6350
rect 2400 6340 2450 6350
rect 4100 6340 4150 6350
rect 5500 6340 5800 6350
rect 6400 6340 6500 6350
rect 6750 6340 6800 6350
rect 1400 6330 1450 6340
rect 1600 6330 1700 6340
rect 2400 6330 2450 6340
rect 4100 6330 4150 6340
rect 5500 6330 5800 6340
rect 6400 6330 6500 6340
rect 6750 6330 6800 6340
rect 1400 6320 1450 6330
rect 1600 6320 1700 6330
rect 2400 6320 2450 6330
rect 4100 6320 4150 6330
rect 5500 6320 5800 6330
rect 6400 6320 6500 6330
rect 6750 6320 6800 6330
rect 1400 6310 1450 6320
rect 1600 6310 1700 6320
rect 2400 6310 2450 6320
rect 4100 6310 4150 6320
rect 5500 6310 5800 6320
rect 6400 6310 6500 6320
rect 6750 6310 6800 6320
rect 1400 6300 1450 6310
rect 1600 6300 1700 6310
rect 2400 6300 2450 6310
rect 4100 6300 4150 6310
rect 5500 6300 5800 6310
rect 6400 6300 6500 6310
rect 6750 6300 6800 6310
rect 1250 6290 1300 6300
rect 1800 6290 1850 6300
rect 2400 6290 2450 6300
rect 4150 6290 4200 6300
rect 5350 6290 5400 6300
rect 5550 6290 5650 6300
rect 6500 6290 6550 6300
rect 6800 6290 6850 6300
rect 9850 6290 9990 6300
rect 1250 6280 1300 6290
rect 1800 6280 1850 6290
rect 2400 6280 2450 6290
rect 4150 6280 4200 6290
rect 5350 6280 5400 6290
rect 5550 6280 5650 6290
rect 6500 6280 6550 6290
rect 6800 6280 6850 6290
rect 9850 6280 9990 6290
rect 1250 6270 1300 6280
rect 1800 6270 1850 6280
rect 2400 6270 2450 6280
rect 4150 6270 4200 6280
rect 5350 6270 5400 6280
rect 5550 6270 5650 6280
rect 6500 6270 6550 6280
rect 6800 6270 6850 6280
rect 9850 6270 9990 6280
rect 1250 6260 1300 6270
rect 1800 6260 1850 6270
rect 2400 6260 2450 6270
rect 4150 6260 4200 6270
rect 5350 6260 5400 6270
rect 5550 6260 5650 6270
rect 6500 6260 6550 6270
rect 6800 6260 6850 6270
rect 9850 6260 9990 6270
rect 1250 6250 1300 6260
rect 1800 6250 1850 6260
rect 2400 6250 2450 6260
rect 4150 6250 4200 6260
rect 5350 6250 5400 6260
rect 5550 6250 5650 6260
rect 6500 6250 6550 6260
rect 6800 6250 6850 6260
rect 9850 6250 9990 6260
rect 1250 6240 1400 6250
rect 1750 6240 1800 6250
rect 2400 6240 2450 6250
rect 4200 6240 4250 6250
rect 5300 6240 5350 6250
rect 5500 6240 5550 6250
rect 6550 6240 6600 6250
rect 6800 6240 6850 6250
rect 9400 6240 9500 6250
rect 9600 6240 9650 6250
rect 1250 6230 1400 6240
rect 1750 6230 1800 6240
rect 2400 6230 2450 6240
rect 4200 6230 4250 6240
rect 5300 6230 5350 6240
rect 5500 6230 5550 6240
rect 6550 6230 6600 6240
rect 6800 6230 6850 6240
rect 9400 6230 9500 6240
rect 9600 6230 9650 6240
rect 1250 6220 1400 6230
rect 1750 6220 1800 6230
rect 2400 6220 2450 6230
rect 4200 6220 4250 6230
rect 5300 6220 5350 6230
rect 5500 6220 5550 6230
rect 6550 6220 6600 6230
rect 6800 6220 6850 6230
rect 9400 6220 9500 6230
rect 9600 6220 9650 6230
rect 1250 6210 1400 6220
rect 1750 6210 1800 6220
rect 2400 6210 2450 6220
rect 4200 6210 4250 6220
rect 5300 6210 5350 6220
rect 5500 6210 5550 6220
rect 6550 6210 6600 6220
rect 6800 6210 6850 6220
rect 9400 6210 9500 6220
rect 9600 6210 9650 6220
rect 1250 6200 1400 6210
rect 1750 6200 1800 6210
rect 2400 6200 2450 6210
rect 4200 6200 4250 6210
rect 5300 6200 5350 6210
rect 5500 6200 5550 6210
rect 6550 6200 6600 6210
rect 6800 6200 6850 6210
rect 9400 6200 9500 6210
rect 9600 6200 9650 6210
rect 1250 6190 1400 6200
rect 2400 6190 2450 6200
rect 5450 6190 5500 6200
rect 6650 6190 6700 6200
rect 6800 6190 6900 6200
rect 9250 6190 9300 6200
rect 9600 6190 9700 6200
rect 1250 6180 1400 6190
rect 2400 6180 2450 6190
rect 5450 6180 5500 6190
rect 6650 6180 6700 6190
rect 6800 6180 6900 6190
rect 9250 6180 9300 6190
rect 9600 6180 9700 6190
rect 1250 6170 1400 6180
rect 2400 6170 2450 6180
rect 5450 6170 5500 6180
rect 6650 6170 6700 6180
rect 6800 6170 6900 6180
rect 9250 6170 9300 6180
rect 9600 6170 9700 6180
rect 1250 6160 1400 6170
rect 2400 6160 2450 6170
rect 5450 6160 5500 6170
rect 6650 6160 6700 6170
rect 6800 6160 6900 6170
rect 9250 6160 9300 6170
rect 9600 6160 9700 6170
rect 1250 6150 1400 6160
rect 2400 6150 2450 6160
rect 5450 6150 5500 6160
rect 6650 6150 6700 6160
rect 6800 6150 6900 6160
rect 9250 6150 9300 6160
rect 9600 6150 9700 6160
rect 1250 6140 1300 6150
rect 1650 6140 1700 6150
rect 5250 6140 5300 6150
rect 5400 6140 5450 6150
rect 6850 6140 6950 6150
rect 9150 6140 9200 6150
rect 1250 6130 1300 6140
rect 1650 6130 1700 6140
rect 5250 6130 5300 6140
rect 5400 6130 5450 6140
rect 6850 6130 6950 6140
rect 9150 6130 9200 6140
rect 1250 6120 1300 6130
rect 1650 6120 1700 6130
rect 5250 6120 5300 6130
rect 5400 6120 5450 6130
rect 6850 6120 6950 6130
rect 9150 6120 9200 6130
rect 1250 6110 1300 6120
rect 1650 6110 1700 6120
rect 5250 6110 5300 6120
rect 5400 6110 5450 6120
rect 6850 6110 6950 6120
rect 9150 6110 9200 6120
rect 1250 6100 1300 6110
rect 1650 6100 1700 6110
rect 5250 6100 5300 6110
rect 5400 6100 5450 6110
rect 6850 6100 6950 6110
rect 9150 6100 9200 6110
rect 1250 6090 1300 6100
rect 1650 6090 1700 6100
rect 3950 6090 4000 6100
rect 5350 6090 5400 6100
rect 6700 6090 6750 6100
rect 6900 6090 6950 6100
rect 9050 6090 9100 6100
rect 1250 6080 1300 6090
rect 1650 6080 1700 6090
rect 3950 6080 4000 6090
rect 5350 6080 5400 6090
rect 6700 6080 6750 6090
rect 6900 6080 6950 6090
rect 9050 6080 9100 6090
rect 1250 6070 1300 6080
rect 1650 6070 1700 6080
rect 3950 6070 4000 6080
rect 5350 6070 5400 6080
rect 6700 6070 6750 6080
rect 6900 6070 6950 6080
rect 9050 6070 9100 6080
rect 1250 6060 1300 6070
rect 1650 6060 1700 6070
rect 3950 6060 4000 6070
rect 5350 6060 5400 6070
rect 6700 6060 6750 6070
rect 6900 6060 6950 6070
rect 9050 6060 9100 6070
rect 1250 6050 1300 6060
rect 1650 6050 1700 6060
rect 3950 6050 4000 6060
rect 5350 6050 5400 6060
rect 6700 6050 6750 6060
rect 6900 6050 6950 6060
rect 9050 6050 9100 6060
rect 850 6040 900 6050
rect 1150 6040 1200 6050
rect 1700 6040 1750 6050
rect 4000 6040 4050 6050
rect 5350 6040 5400 6050
rect 6950 6040 7000 6050
rect 8850 6040 8950 6050
rect 9100 6040 9200 6050
rect 9250 6040 9300 6050
rect 9850 6040 9900 6050
rect 850 6030 900 6040
rect 1150 6030 1200 6040
rect 1700 6030 1750 6040
rect 4000 6030 4050 6040
rect 5350 6030 5400 6040
rect 6950 6030 7000 6040
rect 8850 6030 8950 6040
rect 9100 6030 9200 6040
rect 9250 6030 9300 6040
rect 9850 6030 9900 6040
rect 850 6020 900 6030
rect 1150 6020 1200 6030
rect 1700 6020 1750 6030
rect 4000 6020 4050 6030
rect 5350 6020 5400 6030
rect 6950 6020 7000 6030
rect 8850 6020 8950 6030
rect 9100 6020 9200 6030
rect 9250 6020 9300 6030
rect 9850 6020 9900 6030
rect 850 6010 900 6020
rect 1150 6010 1200 6020
rect 1700 6010 1750 6020
rect 4000 6010 4050 6020
rect 5350 6010 5400 6020
rect 6950 6010 7000 6020
rect 8850 6010 8950 6020
rect 9100 6010 9200 6020
rect 9250 6010 9300 6020
rect 9850 6010 9900 6020
rect 850 6000 900 6010
rect 1150 6000 1200 6010
rect 1700 6000 1750 6010
rect 4000 6000 4050 6010
rect 5350 6000 5400 6010
rect 6950 6000 7000 6010
rect 8850 6000 8950 6010
rect 9100 6000 9200 6010
rect 9250 6000 9300 6010
rect 9850 6000 9900 6010
rect 800 5990 1000 6000
rect 1100 5990 1150 6000
rect 1700 5990 1750 6000
rect 2500 5990 2550 6000
rect 3750 5990 3800 6000
rect 5150 5990 5200 6000
rect 6750 5990 6800 6000
rect 6950 5990 7000 6000
rect 8700 5990 8750 6000
rect 8950 5990 9050 6000
rect 9150 5990 9200 6000
rect 9250 5990 9300 6000
rect 800 5980 1000 5990
rect 1100 5980 1150 5990
rect 1700 5980 1750 5990
rect 2500 5980 2550 5990
rect 3750 5980 3800 5990
rect 5150 5980 5200 5990
rect 6750 5980 6800 5990
rect 6950 5980 7000 5990
rect 8700 5980 8750 5990
rect 8950 5980 9050 5990
rect 9150 5980 9200 5990
rect 9250 5980 9300 5990
rect 800 5970 1000 5980
rect 1100 5970 1150 5980
rect 1700 5970 1750 5980
rect 2500 5970 2550 5980
rect 3750 5970 3800 5980
rect 5150 5970 5200 5980
rect 6750 5970 6800 5980
rect 6950 5970 7000 5980
rect 8700 5970 8750 5980
rect 8950 5970 9050 5980
rect 9150 5970 9200 5980
rect 9250 5970 9300 5980
rect 800 5960 1000 5970
rect 1100 5960 1150 5970
rect 1700 5960 1750 5970
rect 2500 5960 2550 5970
rect 3750 5960 3800 5970
rect 5150 5960 5200 5970
rect 6750 5960 6800 5970
rect 6950 5960 7000 5970
rect 8700 5960 8750 5970
rect 8950 5960 9050 5970
rect 9150 5960 9200 5970
rect 9250 5960 9300 5970
rect 800 5950 1000 5960
rect 1100 5950 1150 5960
rect 1700 5950 1750 5960
rect 2500 5950 2550 5960
rect 3750 5950 3800 5960
rect 5150 5950 5200 5960
rect 6750 5950 6800 5960
rect 6950 5950 7000 5960
rect 8700 5950 8750 5960
rect 8950 5950 9050 5960
rect 9150 5950 9200 5960
rect 9250 5950 9300 5960
rect 700 5940 800 5950
rect 1700 5940 1750 5950
rect 2500 5940 2550 5950
rect 3150 5940 3250 5950
rect 4300 5940 4350 5950
rect 6950 5940 7000 5950
rect 8550 5940 8600 5950
rect 8800 5940 8850 5950
rect 8900 5940 8950 5950
rect 9150 5940 9200 5950
rect 9250 5940 9300 5950
rect 9350 5940 9500 5950
rect 700 5930 800 5940
rect 1700 5930 1750 5940
rect 2500 5930 2550 5940
rect 3150 5930 3250 5940
rect 4300 5930 4350 5940
rect 6950 5930 7000 5940
rect 8550 5930 8600 5940
rect 8800 5930 8850 5940
rect 8900 5930 8950 5940
rect 9150 5930 9200 5940
rect 9250 5930 9300 5940
rect 9350 5930 9500 5940
rect 700 5920 800 5930
rect 1700 5920 1750 5930
rect 2500 5920 2550 5930
rect 3150 5920 3250 5930
rect 4300 5920 4350 5930
rect 6950 5920 7000 5930
rect 8550 5920 8600 5930
rect 8800 5920 8850 5930
rect 8900 5920 8950 5930
rect 9150 5920 9200 5930
rect 9250 5920 9300 5930
rect 9350 5920 9500 5930
rect 700 5910 800 5920
rect 1700 5910 1750 5920
rect 2500 5910 2550 5920
rect 3150 5910 3250 5920
rect 4300 5910 4350 5920
rect 6950 5910 7000 5920
rect 8550 5910 8600 5920
rect 8800 5910 8850 5920
rect 8900 5910 8950 5920
rect 9150 5910 9200 5920
rect 9250 5910 9300 5920
rect 9350 5910 9500 5920
rect 700 5900 800 5910
rect 1700 5900 1750 5910
rect 2500 5900 2550 5910
rect 3150 5900 3250 5910
rect 4300 5900 4350 5910
rect 6950 5900 7000 5910
rect 8550 5900 8600 5910
rect 8800 5900 8850 5910
rect 8900 5900 8950 5910
rect 9150 5900 9200 5910
rect 9250 5900 9300 5910
rect 9350 5900 9500 5910
rect 650 5890 700 5900
rect 750 5890 800 5900
rect 950 5890 1000 5900
rect 1800 5890 1850 5900
rect 2550 5890 2600 5900
rect 3050 5890 3150 5900
rect 3200 5890 3250 5900
rect 5100 5890 5150 5900
rect 5300 5890 5350 5900
rect 6950 5890 7000 5900
rect 8350 5890 8400 5900
rect 8750 5890 8800 5900
rect 8850 5890 8900 5900
rect 9150 5890 9200 5900
rect 9300 5890 9350 5900
rect 650 5880 700 5890
rect 750 5880 800 5890
rect 950 5880 1000 5890
rect 1800 5880 1850 5890
rect 2550 5880 2600 5890
rect 3050 5880 3150 5890
rect 3200 5880 3250 5890
rect 5100 5880 5150 5890
rect 5300 5880 5350 5890
rect 6950 5880 7000 5890
rect 8350 5880 8400 5890
rect 8750 5880 8800 5890
rect 8850 5880 8900 5890
rect 9150 5880 9200 5890
rect 9300 5880 9350 5890
rect 650 5870 700 5880
rect 750 5870 800 5880
rect 950 5870 1000 5880
rect 1800 5870 1850 5880
rect 2550 5870 2600 5880
rect 3050 5870 3150 5880
rect 3200 5870 3250 5880
rect 5100 5870 5150 5880
rect 5300 5870 5350 5880
rect 6950 5870 7000 5880
rect 8350 5870 8400 5880
rect 8750 5870 8800 5880
rect 8850 5870 8900 5880
rect 9150 5870 9200 5880
rect 9300 5870 9350 5880
rect 650 5860 700 5870
rect 750 5860 800 5870
rect 950 5860 1000 5870
rect 1800 5860 1850 5870
rect 2550 5860 2600 5870
rect 3050 5860 3150 5870
rect 3200 5860 3250 5870
rect 5100 5860 5150 5870
rect 5300 5860 5350 5870
rect 6950 5860 7000 5870
rect 8350 5860 8400 5870
rect 8750 5860 8800 5870
rect 8850 5860 8900 5870
rect 9150 5860 9200 5870
rect 9300 5860 9350 5870
rect 650 5850 700 5860
rect 750 5850 800 5860
rect 950 5850 1000 5860
rect 1800 5850 1850 5860
rect 2550 5850 2600 5860
rect 3050 5850 3150 5860
rect 3200 5850 3250 5860
rect 5100 5850 5150 5860
rect 5300 5850 5350 5860
rect 6950 5850 7000 5860
rect 8350 5850 8400 5860
rect 8750 5850 8800 5860
rect 8850 5850 8900 5860
rect 9150 5850 9200 5860
rect 9300 5850 9350 5860
rect 600 5840 650 5850
rect 700 5840 750 5850
rect 2300 5840 2350 5850
rect 2600 5840 2650 5850
rect 3000 5840 3050 5850
rect 3200 5840 3250 5850
rect 3750 5840 3850 5850
rect 5300 5840 5350 5850
rect 8200 5840 8250 5850
rect 8700 5840 8750 5850
rect 8850 5840 8900 5850
rect 8950 5840 9000 5850
rect 9050 5840 9200 5850
rect 9900 5840 9950 5850
rect 600 5830 650 5840
rect 700 5830 750 5840
rect 2300 5830 2350 5840
rect 2600 5830 2650 5840
rect 3000 5830 3050 5840
rect 3200 5830 3250 5840
rect 3750 5830 3850 5840
rect 5300 5830 5350 5840
rect 8200 5830 8250 5840
rect 8700 5830 8750 5840
rect 8850 5830 8900 5840
rect 8950 5830 9000 5840
rect 9050 5830 9200 5840
rect 9900 5830 9950 5840
rect 600 5820 650 5830
rect 700 5820 750 5830
rect 2300 5820 2350 5830
rect 2600 5820 2650 5830
rect 3000 5820 3050 5830
rect 3200 5820 3250 5830
rect 3750 5820 3850 5830
rect 5300 5820 5350 5830
rect 8200 5820 8250 5830
rect 8700 5820 8750 5830
rect 8850 5820 8900 5830
rect 8950 5820 9000 5830
rect 9050 5820 9200 5830
rect 9900 5820 9950 5830
rect 600 5810 650 5820
rect 700 5810 750 5820
rect 2300 5810 2350 5820
rect 2600 5810 2650 5820
rect 3000 5810 3050 5820
rect 3200 5810 3250 5820
rect 3750 5810 3850 5820
rect 5300 5810 5350 5820
rect 8200 5810 8250 5820
rect 8700 5810 8750 5820
rect 8850 5810 8900 5820
rect 8950 5810 9000 5820
rect 9050 5810 9200 5820
rect 9900 5810 9950 5820
rect 600 5800 650 5810
rect 700 5800 750 5810
rect 2300 5800 2350 5810
rect 2600 5800 2650 5810
rect 3000 5800 3050 5810
rect 3200 5800 3250 5810
rect 3750 5800 3850 5810
rect 5300 5800 5350 5810
rect 8200 5800 8250 5810
rect 8700 5800 8750 5810
rect 8850 5800 8900 5810
rect 8950 5800 9000 5810
rect 9050 5800 9200 5810
rect 9900 5800 9950 5810
rect 650 5790 700 5800
rect 800 5790 900 5800
rect 1850 5790 1900 5800
rect 2250 5790 2350 5800
rect 2550 5790 2650 5800
rect 2900 5790 3000 5800
rect 3200 5790 3250 5800
rect 3850 5790 3900 5800
rect 6800 5790 6850 5800
rect 6950 5790 7000 5800
rect 8050 5790 8100 5800
rect 8350 5790 8450 5800
rect 8650 5790 8700 5800
rect 8800 5790 8850 5800
rect 650 5780 700 5790
rect 800 5780 900 5790
rect 1850 5780 1900 5790
rect 2250 5780 2350 5790
rect 2550 5780 2650 5790
rect 2900 5780 3000 5790
rect 3200 5780 3250 5790
rect 3850 5780 3900 5790
rect 6800 5780 6850 5790
rect 6950 5780 7000 5790
rect 8050 5780 8100 5790
rect 8350 5780 8450 5790
rect 8650 5780 8700 5790
rect 8800 5780 8850 5790
rect 650 5770 700 5780
rect 800 5770 900 5780
rect 1850 5770 1900 5780
rect 2250 5770 2350 5780
rect 2550 5770 2650 5780
rect 2900 5770 3000 5780
rect 3200 5770 3250 5780
rect 3850 5770 3900 5780
rect 6800 5770 6850 5780
rect 6950 5770 7000 5780
rect 8050 5770 8100 5780
rect 8350 5770 8450 5780
rect 8650 5770 8700 5780
rect 8800 5770 8850 5780
rect 650 5760 700 5770
rect 800 5760 900 5770
rect 1850 5760 1900 5770
rect 2250 5760 2350 5770
rect 2550 5760 2650 5770
rect 2900 5760 3000 5770
rect 3200 5760 3250 5770
rect 3850 5760 3900 5770
rect 6800 5760 6850 5770
rect 6950 5760 7000 5770
rect 8050 5760 8100 5770
rect 8350 5760 8450 5770
rect 8650 5760 8700 5770
rect 8800 5760 8850 5770
rect 650 5750 700 5760
rect 800 5750 900 5760
rect 1850 5750 1900 5760
rect 2250 5750 2350 5760
rect 2550 5750 2650 5760
rect 2900 5750 3000 5760
rect 3200 5750 3250 5760
rect 3850 5750 3900 5760
rect 6800 5750 6850 5760
rect 6950 5750 7000 5760
rect 8050 5750 8100 5760
rect 8350 5750 8450 5760
rect 8650 5750 8700 5760
rect 8800 5750 8850 5760
rect 2200 5740 2300 5750
rect 2500 5740 2550 5750
rect 2800 5740 2950 5750
rect 3200 5740 3250 5750
rect 3950 5740 4000 5750
rect 6800 5740 6850 5750
rect 6950 5740 7000 5750
rect 7900 5740 7950 5750
rect 8150 5740 8300 5750
rect 8350 5740 8400 5750
rect 2200 5730 2300 5740
rect 2500 5730 2550 5740
rect 2800 5730 2950 5740
rect 3200 5730 3250 5740
rect 3950 5730 4000 5740
rect 6800 5730 6850 5740
rect 6950 5730 7000 5740
rect 7900 5730 7950 5740
rect 8150 5730 8300 5740
rect 8350 5730 8400 5740
rect 2200 5720 2300 5730
rect 2500 5720 2550 5730
rect 2800 5720 2950 5730
rect 3200 5720 3250 5730
rect 3950 5720 4000 5730
rect 6800 5720 6850 5730
rect 6950 5720 7000 5730
rect 7900 5720 7950 5730
rect 8150 5720 8300 5730
rect 8350 5720 8400 5730
rect 2200 5710 2300 5720
rect 2500 5710 2550 5720
rect 2800 5710 2950 5720
rect 3200 5710 3250 5720
rect 3950 5710 4000 5720
rect 6800 5710 6850 5720
rect 6950 5710 7000 5720
rect 7900 5710 7950 5720
rect 8150 5710 8300 5720
rect 8350 5710 8400 5720
rect 2200 5700 2300 5710
rect 2500 5700 2550 5710
rect 2800 5700 2950 5710
rect 3200 5700 3250 5710
rect 3950 5700 4000 5710
rect 6800 5700 6850 5710
rect 6950 5700 7000 5710
rect 7900 5700 7950 5710
rect 8150 5700 8300 5710
rect 8350 5700 8400 5710
rect 1900 5690 1950 5700
rect 2250 5690 2300 5700
rect 2450 5690 2500 5700
rect 2750 5690 2800 5700
rect 3200 5690 3250 5700
rect 3950 5690 4000 5700
rect 7700 5690 7750 5700
rect 7850 5690 7900 5700
rect 8000 5690 8100 5700
rect 8450 5690 8500 5700
rect 1900 5680 1950 5690
rect 2250 5680 2300 5690
rect 2450 5680 2500 5690
rect 2750 5680 2800 5690
rect 3200 5680 3250 5690
rect 3950 5680 4000 5690
rect 7700 5680 7750 5690
rect 7850 5680 7900 5690
rect 8000 5680 8100 5690
rect 8450 5680 8500 5690
rect 1900 5670 1950 5680
rect 2250 5670 2300 5680
rect 2450 5670 2500 5680
rect 2750 5670 2800 5680
rect 3200 5670 3250 5680
rect 3950 5670 4000 5680
rect 7700 5670 7750 5680
rect 7850 5670 7900 5680
rect 8000 5670 8100 5680
rect 8450 5670 8500 5680
rect 1900 5660 1950 5670
rect 2250 5660 2300 5670
rect 2450 5660 2500 5670
rect 2750 5660 2800 5670
rect 3200 5660 3250 5670
rect 3950 5660 4000 5670
rect 7700 5660 7750 5670
rect 7850 5660 7900 5670
rect 8000 5660 8100 5670
rect 8450 5660 8500 5670
rect 1900 5650 1950 5660
rect 2250 5650 2300 5660
rect 2450 5650 2500 5660
rect 2750 5650 2800 5660
rect 3200 5650 3250 5660
rect 3950 5650 4000 5660
rect 7700 5650 7750 5660
rect 7850 5650 7900 5660
rect 8000 5650 8100 5660
rect 8450 5650 8500 5660
rect 2150 5640 2200 5650
rect 2450 5640 2500 5650
rect 2700 5640 2800 5650
rect 3200 5640 3250 5650
rect 5100 5640 5150 5650
rect 5250 5640 5300 5650
rect 5600 5640 5800 5650
rect 6850 5640 6900 5650
rect 7550 5640 7700 5650
rect 7800 5640 7850 5650
rect 7900 5640 7950 5650
rect 8000 5640 8050 5650
rect 8300 5640 8400 5650
rect 2150 5630 2200 5640
rect 2450 5630 2500 5640
rect 2700 5630 2800 5640
rect 3200 5630 3250 5640
rect 5100 5630 5150 5640
rect 5250 5630 5300 5640
rect 5600 5630 5800 5640
rect 6850 5630 6900 5640
rect 7550 5630 7700 5640
rect 7800 5630 7850 5640
rect 7900 5630 7950 5640
rect 8000 5630 8050 5640
rect 8300 5630 8400 5640
rect 2150 5620 2200 5630
rect 2450 5620 2500 5630
rect 2700 5620 2800 5630
rect 3200 5620 3250 5630
rect 5100 5620 5150 5630
rect 5250 5620 5300 5630
rect 5600 5620 5800 5630
rect 6850 5620 6900 5630
rect 7550 5620 7700 5630
rect 7800 5620 7850 5630
rect 7900 5620 7950 5630
rect 8000 5620 8050 5630
rect 8300 5620 8400 5630
rect 2150 5610 2200 5620
rect 2450 5610 2500 5620
rect 2700 5610 2800 5620
rect 3200 5610 3250 5620
rect 5100 5610 5150 5620
rect 5250 5610 5300 5620
rect 5600 5610 5800 5620
rect 6850 5610 6900 5620
rect 7550 5610 7700 5620
rect 7800 5610 7850 5620
rect 7900 5610 7950 5620
rect 8000 5610 8050 5620
rect 8300 5610 8400 5620
rect 2150 5600 2200 5610
rect 2450 5600 2500 5610
rect 2700 5600 2800 5610
rect 3200 5600 3250 5610
rect 5100 5600 5150 5610
rect 5250 5600 5300 5610
rect 5600 5600 5800 5610
rect 6850 5600 6900 5610
rect 7550 5600 7700 5610
rect 7800 5600 7850 5610
rect 7900 5600 7950 5610
rect 8000 5600 8050 5610
rect 8300 5600 8400 5610
rect 650 5590 700 5600
rect 1950 5590 2000 5600
rect 2150 5590 2200 5600
rect 2400 5590 2450 5600
rect 2650 5590 2700 5600
rect 2850 5590 2950 5600
rect 3200 5590 3250 5600
rect 3750 5590 3800 5600
rect 5500 5590 5600 5600
rect 5850 5590 5950 5600
rect 6200 5590 6300 5600
rect 6450 5590 6550 5600
rect 7400 5590 7450 5600
rect 7600 5590 7700 5600
rect 7750 5590 7800 5600
rect 8000 5590 8050 5600
rect 8250 5590 8400 5600
rect 9050 5590 9100 5600
rect 650 5580 700 5590
rect 1950 5580 2000 5590
rect 2150 5580 2200 5590
rect 2400 5580 2450 5590
rect 2650 5580 2700 5590
rect 2850 5580 2950 5590
rect 3200 5580 3250 5590
rect 3750 5580 3800 5590
rect 5500 5580 5600 5590
rect 5850 5580 5950 5590
rect 6200 5580 6300 5590
rect 6450 5580 6550 5590
rect 7400 5580 7450 5590
rect 7600 5580 7700 5590
rect 7750 5580 7800 5590
rect 8000 5580 8050 5590
rect 8250 5580 8400 5590
rect 9050 5580 9100 5590
rect 650 5570 700 5580
rect 1950 5570 2000 5580
rect 2150 5570 2200 5580
rect 2400 5570 2450 5580
rect 2650 5570 2700 5580
rect 2850 5570 2950 5580
rect 3200 5570 3250 5580
rect 3750 5570 3800 5580
rect 5500 5570 5600 5580
rect 5850 5570 5950 5580
rect 6200 5570 6300 5580
rect 6450 5570 6550 5580
rect 7400 5570 7450 5580
rect 7600 5570 7700 5580
rect 7750 5570 7800 5580
rect 8000 5570 8050 5580
rect 8250 5570 8400 5580
rect 9050 5570 9100 5580
rect 650 5560 700 5570
rect 1950 5560 2000 5570
rect 2150 5560 2200 5570
rect 2400 5560 2450 5570
rect 2650 5560 2700 5570
rect 2850 5560 2950 5570
rect 3200 5560 3250 5570
rect 3750 5560 3800 5570
rect 5500 5560 5600 5570
rect 5850 5560 5950 5570
rect 6200 5560 6300 5570
rect 6450 5560 6550 5570
rect 7400 5560 7450 5570
rect 7600 5560 7700 5570
rect 7750 5560 7800 5570
rect 8000 5560 8050 5570
rect 8250 5560 8400 5570
rect 9050 5560 9100 5570
rect 650 5550 700 5560
rect 1950 5550 2000 5560
rect 2150 5550 2200 5560
rect 2400 5550 2450 5560
rect 2650 5550 2700 5560
rect 2850 5550 2950 5560
rect 3200 5550 3250 5560
rect 3750 5550 3800 5560
rect 5500 5550 5600 5560
rect 5850 5550 5950 5560
rect 6200 5550 6300 5560
rect 6450 5550 6550 5560
rect 7400 5550 7450 5560
rect 7600 5550 7700 5560
rect 7750 5550 7800 5560
rect 8000 5550 8050 5560
rect 8250 5550 8400 5560
rect 9050 5550 9100 5560
rect 500 5540 650 5550
rect 1950 5540 2000 5550
rect 2150 5540 2200 5550
rect 2350 5540 2400 5550
rect 2600 5540 2700 5550
rect 2800 5540 3000 5550
rect 3200 5540 3250 5550
rect 3700 5540 3750 5550
rect 5100 5540 5150 5550
rect 5500 5540 5650 5550
rect 5950 5540 6000 5550
rect 6150 5540 6200 5550
rect 6550 5540 6600 5550
rect 7350 5540 7400 5550
rect 7500 5540 7550 5550
rect 7700 5540 7750 5550
rect 8750 5540 8850 5550
rect 8900 5540 8950 5550
rect 9050 5540 9100 5550
rect 500 5530 650 5540
rect 1950 5530 2000 5540
rect 2150 5530 2200 5540
rect 2350 5530 2400 5540
rect 2600 5530 2700 5540
rect 2800 5530 3000 5540
rect 3200 5530 3250 5540
rect 3700 5530 3750 5540
rect 5100 5530 5150 5540
rect 5500 5530 5650 5540
rect 5950 5530 6000 5540
rect 6150 5530 6200 5540
rect 6550 5530 6600 5540
rect 7350 5530 7400 5540
rect 7500 5530 7550 5540
rect 7700 5530 7750 5540
rect 8750 5530 8850 5540
rect 8900 5530 8950 5540
rect 9050 5530 9100 5540
rect 500 5520 650 5530
rect 1950 5520 2000 5530
rect 2150 5520 2200 5530
rect 2350 5520 2400 5530
rect 2600 5520 2700 5530
rect 2800 5520 3000 5530
rect 3200 5520 3250 5530
rect 3700 5520 3750 5530
rect 5100 5520 5150 5530
rect 5500 5520 5650 5530
rect 5950 5520 6000 5530
rect 6150 5520 6200 5530
rect 6550 5520 6600 5530
rect 7350 5520 7400 5530
rect 7500 5520 7550 5530
rect 7700 5520 7750 5530
rect 8750 5520 8850 5530
rect 8900 5520 8950 5530
rect 9050 5520 9100 5530
rect 500 5510 650 5520
rect 1950 5510 2000 5520
rect 2150 5510 2200 5520
rect 2350 5510 2400 5520
rect 2600 5510 2700 5520
rect 2800 5510 3000 5520
rect 3200 5510 3250 5520
rect 3700 5510 3750 5520
rect 5100 5510 5150 5520
rect 5500 5510 5650 5520
rect 5950 5510 6000 5520
rect 6150 5510 6200 5520
rect 6550 5510 6600 5520
rect 7350 5510 7400 5520
rect 7500 5510 7550 5520
rect 7700 5510 7750 5520
rect 8750 5510 8850 5520
rect 8900 5510 8950 5520
rect 9050 5510 9100 5520
rect 500 5500 650 5510
rect 1950 5500 2000 5510
rect 2150 5500 2200 5510
rect 2350 5500 2400 5510
rect 2600 5500 2700 5510
rect 2800 5500 3000 5510
rect 3200 5500 3250 5510
rect 3700 5500 3750 5510
rect 5100 5500 5150 5510
rect 5500 5500 5650 5510
rect 5950 5500 6000 5510
rect 6150 5500 6200 5510
rect 6550 5500 6600 5510
rect 7350 5500 7400 5510
rect 7500 5500 7550 5510
rect 7700 5500 7750 5510
rect 8750 5500 8850 5510
rect 8900 5500 8950 5510
rect 9050 5500 9100 5510
rect 1950 5490 2000 5500
rect 2150 5490 2200 5500
rect 2350 5490 2400 5500
rect 2600 5490 2850 5500
rect 2950 5490 3050 5500
rect 3150 5490 3200 5500
rect 3600 5490 3650 5500
rect 5450 5490 5550 5500
rect 5600 5490 5650 5500
rect 6150 5490 6200 5500
rect 6500 5490 6600 5500
rect 6900 5490 6950 5500
rect 7350 5490 7400 5500
rect 8600 5490 8700 5500
rect 9000 5490 9050 5500
rect 9100 5490 9150 5500
rect 1950 5480 2000 5490
rect 2150 5480 2200 5490
rect 2350 5480 2400 5490
rect 2600 5480 2850 5490
rect 2950 5480 3050 5490
rect 3150 5480 3200 5490
rect 3600 5480 3650 5490
rect 5450 5480 5550 5490
rect 5600 5480 5650 5490
rect 6150 5480 6200 5490
rect 6500 5480 6600 5490
rect 6900 5480 6950 5490
rect 7350 5480 7400 5490
rect 8600 5480 8700 5490
rect 9000 5480 9050 5490
rect 9100 5480 9150 5490
rect 1950 5470 2000 5480
rect 2150 5470 2200 5480
rect 2350 5470 2400 5480
rect 2600 5470 2850 5480
rect 2950 5470 3050 5480
rect 3150 5470 3200 5480
rect 3600 5470 3650 5480
rect 5450 5470 5550 5480
rect 5600 5470 5650 5480
rect 6150 5470 6200 5480
rect 6500 5470 6600 5480
rect 6900 5470 6950 5480
rect 7350 5470 7400 5480
rect 8600 5470 8700 5480
rect 9000 5470 9050 5480
rect 9100 5470 9150 5480
rect 1950 5460 2000 5470
rect 2150 5460 2200 5470
rect 2350 5460 2400 5470
rect 2600 5460 2850 5470
rect 2950 5460 3050 5470
rect 3150 5460 3200 5470
rect 3600 5460 3650 5470
rect 5450 5460 5550 5470
rect 5600 5460 5650 5470
rect 6150 5460 6200 5470
rect 6500 5460 6600 5470
rect 6900 5460 6950 5470
rect 7350 5460 7400 5470
rect 8600 5460 8700 5470
rect 9000 5460 9050 5470
rect 9100 5460 9150 5470
rect 1950 5450 2000 5460
rect 2150 5450 2200 5460
rect 2350 5450 2400 5460
rect 2600 5450 2850 5460
rect 2950 5450 3050 5460
rect 3150 5450 3200 5460
rect 3600 5450 3650 5460
rect 5450 5450 5550 5460
rect 5600 5450 5650 5460
rect 6150 5450 6200 5460
rect 6500 5450 6600 5460
rect 6900 5450 6950 5460
rect 7350 5450 7400 5460
rect 8600 5450 8700 5460
rect 9000 5450 9050 5460
rect 9100 5450 9150 5460
rect 550 5440 600 5450
rect 2000 5440 2050 5450
rect 2150 5440 2250 5450
rect 2350 5440 2400 5450
rect 2650 5440 2850 5450
rect 3050 5440 3150 5450
rect 3550 5440 3600 5450
rect 5200 5440 5250 5450
rect 6150 5440 6200 5450
rect 6600 5440 6650 5450
rect 7250 5440 7350 5450
rect 7750 5440 7950 5450
rect 8350 5440 8400 5450
rect 8450 5440 8500 5450
rect 8950 5440 9000 5450
rect 9550 5440 9600 5450
rect 550 5430 600 5440
rect 2000 5430 2050 5440
rect 2150 5430 2250 5440
rect 2350 5430 2400 5440
rect 2650 5430 2850 5440
rect 3050 5430 3150 5440
rect 3550 5430 3600 5440
rect 5200 5430 5250 5440
rect 6150 5430 6200 5440
rect 6600 5430 6650 5440
rect 7250 5430 7350 5440
rect 7750 5430 7950 5440
rect 8350 5430 8400 5440
rect 8450 5430 8500 5440
rect 8950 5430 9000 5440
rect 9550 5430 9600 5440
rect 550 5420 600 5430
rect 2000 5420 2050 5430
rect 2150 5420 2250 5430
rect 2350 5420 2400 5430
rect 2650 5420 2850 5430
rect 3050 5420 3150 5430
rect 3550 5420 3600 5430
rect 5200 5420 5250 5430
rect 6150 5420 6200 5430
rect 6600 5420 6650 5430
rect 7250 5420 7350 5430
rect 7750 5420 7950 5430
rect 8350 5420 8400 5430
rect 8450 5420 8500 5430
rect 8950 5420 9000 5430
rect 9550 5420 9600 5430
rect 550 5410 600 5420
rect 2000 5410 2050 5420
rect 2150 5410 2250 5420
rect 2350 5410 2400 5420
rect 2650 5410 2850 5420
rect 3050 5410 3150 5420
rect 3550 5410 3600 5420
rect 5200 5410 5250 5420
rect 6150 5410 6200 5420
rect 6600 5410 6650 5420
rect 7250 5410 7350 5420
rect 7750 5410 7950 5420
rect 8350 5410 8400 5420
rect 8450 5410 8500 5420
rect 8950 5410 9000 5420
rect 9550 5410 9600 5420
rect 550 5400 600 5410
rect 2000 5400 2050 5410
rect 2150 5400 2250 5410
rect 2350 5400 2400 5410
rect 2650 5400 2850 5410
rect 3050 5400 3150 5410
rect 3550 5400 3600 5410
rect 5200 5400 5250 5410
rect 6150 5400 6200 5410
rect 6600 5400 6650 5410
rect 7250 5400 7350 5410
rect 7750 5400 7950 5410
rect 8350 5400 8400 5410
rect 8450 5400 8500 5410
rect 8950 5400 9000 5410
rect 9550 5400 9600 5410
rect 350 5390 400 5400
rect 450 5390 500 5400
rect 2000 5390 2250 5400
rect 2350 5390 2400 5400
rect 5200 5390 5250 5400
rect 5400 5390 5450 5400
rect 5900 5390 5950 5400
rect 6150 5390 6200 5400
rect 7300 5390 7350 5400
rect 7500 5390 7550 5400
rect 7600 5390 7750 5400
rect 8250 5390 8300 5400
rect 8500 5390 8550 5400
rect 8850 5390 8950 5400
rect 9400 5390 9450 5400
rect 9550 5390 9600 5400
rect 350 5380 400 5390
rect 450 5380 500 5390
rect 2000 5380 2250 5390
rect 2350 5380 2400 5390
rect 5200 5380 5250 5390
rect 5400 5380 5450 5390
rect 5900 5380 5950 5390
rect 6150 5380 6200 5390
rect 7300 5380 7350 5390
rect 7500 5380 7550 5390
rect 7600 5380 7750 5390
rect 8250 5380 8300 5390
rect 8500 5380 8550 5390
rect 8850 5380 8950 5390
rect 9400 5380 9450 5390
rect 9550 5380 9600 5390
rect 350 5370 400 5380
rect 450 5370 500 5380
rect 2000 5370 2250 5380
rect 2350 5370 2400 5380
rect 5200 5370 5250 5380
rect 5400 5370 5450 5380
rect 5900 5370 5950 5380
rect 6150 5370 6200 5380
rect 7300 5370 7350 5380
rect 7500 5370 7550 5380
rect 7600 5370 7750 5380
rect 8250 5370 8300 5380
rect 8500 5370 8550 5380
rect 8850 5370 8950 5380
rect 9400 5370 9450 5380
rect 9550 5370 9600 5380
rect 350 5360 400 5370
rect 450 5360 500 5370
rect 2000 5360 2250 5370
rect 2350 5360 2400 5370
rect 5200 5360 5250 5370
rect 5400 5360 5450 5370
rect 5900 5360 5950 5370
rect 6150 5360 6200 5370
rect 7300 5360 7350 5370
rect 7500 5360 7550 5370
rect 7600 5360 7750 5370
rect 8250 5360 8300 5370
rect 8500 5360 8550 5370
rect 8850 5360 8950 5370
rect 9400 5360 9450 5370
rect 9550 5360 9600 5370
rect 350 5350 400 5360
rect 450 5350 500 5360
rect 2000 5350 2250 5360
rect 2350 5350 2400 5360
rect 5200 5350 5250 5360
rect 5400 5350 5450 5360
rect 5900 5350 5950 5360
rect 6150 5350 6200 5360
rect 7300 5350 7350 5360
rect 7500 5350 7550 5360
rect 7600 5350 7750 5360
rect 8250 5350 8300 5360
rect 8500 5350 8550 5360
rect 8850 5350 8950 5360
rect 9400 5350 9450 5360
rect 9550 5350 9600 5360
rect 250 5340 450 5350
rect 2050 5340 2250 5350
rect 2350 5340 2400 5350
rect 5100 5340 5150 5350
rect 5200 5340 5250 5350
rect 5650 5340 5700 5350
rect 5850 5340 5900 5350
rect 6150 5340 6200 5350
rect 7300 5340 7350 5350
rect 8050 5340 8100 5350
rect 8150 5340 8250 5350
rect 8300 5340 8350 5350
rect 8500 5340 8550 5350
rect 8700 5340 8800 5350
rect 9300 5340 9350 5350
rect 9400 5340 9450 5350
rect 9500 5340 9550 5350
rect 250 5330 450 5340
rect 2050 5330 2250 5340
rect 2350 5330 2400 5340
rect 5100 5330 5150 5340
rect 5200 5330 5250 5340
rect 5650 5330 5700 5340
rect 5850 5330 5900 5340
rect 6150 5330 6200 5340
rect 7300 5330 7350 5340
rect 8050 5330 8100 5340
rect 8150 5330 8250 5340
rect 8300 5330 8350 5340
rect 8500 5330 8550 5340
rect 8700 5330 8800 5340
rect 9300 5330 9350 5340
rect 9400 5330 9450 5340
rect 9500 5330 9550 5340
rect 250 5320 450 5330
rect 2050 5320 2250 5330
rect 2350 5320 2400 5330
rect 5100 5320 5150 5330
rect 5200 5320 5250 5330
rect 5650 5320 5700 5330
rect 5850 5320 5900 5330
rect 6150 5320 6200 5330
rect 7300 5320 7350 5330
rect 8050 5320 8100 5330
rect 8150 5320 8250 5330
rect 8300 5320 8350 5330
rect 8500 5320 8550 5330
rect 8700 5320 8800 5330
rect 9300 5320 9350 5330
rect 9400 5320 9450 5330
rect 9500 5320 9550 5330
rect 250 5310 450 5320
rect 2050 5310 2250 5320
rect 2350 5310 2400 5320
rect 5100 5310 5150 5320
rect 5200 5310 5250 5320
rect 5650 5310 5700 5320
rect 5850 5310 5900 5320
rect 6150 5310 6200 5320
rect 7300 5310 7350 5320
rect 8050 5310 8100 5320
rect 8150 5310 8250 5320
rect 8300 5310 8350 5320
rect 8500 5310 8550 5320
rect 8700 5310 8800 5320
rect 9300 5310 9350 5320
rect 9400 5310 9450 5320
rect 9500 5310 9550 5320
rect 250 5300 450 5310
rect 2050 5300 2250 5310
rect 2350 5300 2400 5310
rect 5100 5300 5150 5310
rect 5200 5300 5250 5310
rect 5650 5300 5700 5310
rect 5850 5300 5900 5310
rect 6150 5300 6200 5310
rect 7300 5300 7350 5310
rect 8050 5300 8100 5310
rect 8150 5300 8250 5310
rect 8300 5300 8350 5310
rect 8500 5300 8550 5310
rect 8700 5300 8800 5310
rect 9300 5300 9350 5310
rect 9400 5300 9450 5310
rect 9500 5300 9550 5310
rect 300 5290 350 5300
rect 550 5290 600 5300
rect 2050 5290 2250 5300
rect 2350 5290 2400 5300
rect 2450 5290 2600 5300
rect 2650 5290 2750 5300
rect 3500 5290 3550 5300
rect 5100 5290 5150 5300
rect 5650 5290 5850 5300
rect 6200 5290 6250 5300
rect 6450 5290 6500 5300
rect 7250 5290 7300 5300
rect 7950 5290 8000 5300
rect 8350 5290 8400 5300
rect 8550 5290 8600 5300
rect 9050 5290 9200 5300
rect 9250 5290 9600 5300
rect 9850 5290 9900 5300
rect 9950 5290 9990 5300
rect 300 5280 350 5290
rect 550 5280 600 5290
rect 2050 5280 2250 5290
rect 2350 5280 2400 5290
rect 2450 5280 2600 5290
rect 2650 5280 2750 5290
rect 3500 5280 3550 5290
rect 5100 5280 5150 5290
rect 5650 5280 5850 5290
rect 6200 5280 6250 5290
rect 6450 5280 6500 5290
rect 7250 5280 7300 5290
rect 7950 5280 8000 5290
rect 8350 5280 8400 5290
rect 8550 5280 8600 5290
rect 9050 5280 9200 5290
rect 9250 5280 9600 5290
rect 9850 5280 9900 5290
rect 9950 5280 9990 5290
rect 300 5270 350 5280
rect 550 5270 600 5280
rect 2050 5270 2250 5280
rect 2350 5270 2400 5280
rect 2450 5270 2600 5280
rect 2650 5270 2750 5280
rect 3500 5270 3550 5280
rect 5100 5270 5150 5280
rect 5650 5270 5850 5280
rect 6200 5270 6250 5280
rect 6450 5270 6500 5280
rect 7250 5270 7300 5280
rect 7950 5270 8000 5280
rect 8350 5270 8400 5280
rect 8550 5270 8600 5280
rect 9050 5270 9200 5280
rect 9250 5270 9600 5280
rect 9850 5270 9900 5280
rect 9950 5270 9990 5280
rect 300 5260 350 5270
rect 550 5260 600 5270
rect 2050 5260 2250 5270
rect 2350 5260 2400 5270
rect 2450 5260 2600 5270
rect 2650 5260 2750 5270
rect 3500 5260 3550 5270
rect 5100 5260 5150 5270
rect 5650 5260 5850 5270
rect 6200 5260 6250 5270
rect 6450 5260 6500 5270
rect 7250 5260 7300 5270
rect 7950 5260 8000 5270
rect 8350 5260 8400 5270
rect 8550 5260 8600 5270
rect 9050 5260 9200 5270
rect 9250 5260 9600 5270
rect 9850 5260 9900 5270
rect 9950 5260 9990 5270
rect 300 5250 350 5260
rect 550 5250 600 5260
rect 2050 5250 2250 5260
rect 2350 5250 2400 5260
rect 2450 5250 2600 5260
rect 2650 5250 2750 5260
rect 3500 5250 3550 5260
rect 5100 5250 5150 5260
rect 5650 5250 5850 5260
rect 6200 5250 6250 5260
rect 6450 5250 6500 5260
rect 7250 5250 7300 5260
rect 7950 5250 8000 5260
rect 8350 5250 8400 5260
rect 8550 5250 8600 5260
rect 9050 5250 9200 5260
rect 9250 5250 9600 5260
rect 9850 5250 9900 5260
rect 9950 5250 9990 5260
rect 2050 5240 2250 5250
rect 2350 5240 2500 5250
rect 2650 5240 2900 5250
rect 5050 5240 5100 5250
rect 5150 5240 5200 5250
rect 6350 5240 6550 5250
rect 7950 5240 8000 5250
rect 8350 5240 8400 5250
rect 8850 5240 8950 5250
rect 9300 5240 9400 5250
rect 9700 5240 9750 5250
rect 9800 5240 9850 5250
rect 9900 5240 9950 5250
rect 2050 5230 2250 5240
rect 2350 5230 2500 5240
rect 2650 5230 2900 5240
rect 5050 5230 5100 5240
rect 5150 5230 5200 5240
rect 6350 5230 6550 5240
rect 7950 5230 8000 5240
rect 8350 5230 8400 5240
rect 8850 5230 8950 5240
rect 9300 5230 9400 5240
rect 9700 5230 9750 5240
rect 9800 5230 9850 5240
rect 9900 5230 9950 5240
rect 2050 5220 2250 5230
rect 2350 5220 2500 5230
rect 2650 5220 2900 5230
rect 5050 5220 5100 5230
rect 5150 5220 5200 5230
rect 6350 5220 6550 5230
rect 7950 5220 8000 5230
rect 8350 5220 8400 5230
rect 8850 5220 8950 5230
rect 9300 5220 9400 5230
rect 9700 5220 9750 5230
rect 9800 5220 9850 5230
rect 9900 5220 9950 5230
rect 2050 5210 2250 5220
rect 2350 5210 2500 5220
rect 2650 5210 2900 5220
rect 5050 5210 5100 5220
rect 5150 5210 5200 5220
rect 6350 5210 6550 5220
rect 7950 5210 8000 5220
rect 8350 5210 8400 5220
rect 8850 5210 8950 5220
rect 9300 5210 9400 5220
rect 9700 5210 9750 5220
rect 9800 5210 9850 5220
rect 9900 5210 9950 5220
rect 2050 5200 2250 5210
rect 2350 5200 2500 5210
rect 2650 5200 2900 5210
rect 5050 5200 5100 5210
rect 5150 5200 5200 5210
rect 6350 5200 6550 5210
rect 7950 5200 8000 5210
rect 8350 5200 8400 5210
rect 8850 5200 8950 5210
rect 9300 5200 9400 5210
rect 9700 5200 9750 5210
rect 9800 5200 9850 5210
rect 9900 5200 9950 5210
rect 2050 5190 2250 5200
rect 2350 5190 2500 5200
rect 2800 5190 2900 5200
rect 3450 5190 3500 5200
rect 7300 5190 7350 5200
rect 8000 5190 8050 5200
rect 8200 5190 8250 5200
rect 8600 5190 8650 5200
rect 8700 5190 8750 5200
rect 8800 5190 8950 5200
rect 9000 5190 9200 5200
rect 9500 5190 9600 5200
rect 9800 5190 9950 5200
rect 2050 5180 2250 5190
rect 2350 5180 2500 5190
rect 2800 5180 2900 5190
rect 3450 5180 3500 5190
rect 7300 5180 7350 5190
rect 8000 5180 8050 5190
rect 8200 5180 8250 5190
rect 8600 5180 8650 5190
rect 8700 5180 8750 5190
rect 8800 5180 8950 5190
rect 9000 5180 9200 5190
rect 9500 5180 9600 5190
rect 9800 5180 9950 5190
rect 2050 5170 2250 5180
rect 2350 5170 2500 5180
rect 2800 5170 2900 5180
rect 3450 5170 3500 5180
rect 7300 5170 7350 5180
rect 8000 5170 8050 5180
rect 8200 5170 8250 5180
rect 8600 5170 8650 5180
rect 8700 5170 8750 5180
rect 8800 5170 8950 5180
rect 9000 5170 9200 5180
rect 9500 5170 9600 5180
rect 9800 5170 9950 5180
rect 2050 5160 2250 5170
rect 2350 5160 2500 5170
rect 2800 5160 2900 5170
rect 3450 5160 3500 5170
rect 7300 5160 7350 5170
rect 8000 5160 8050 5170
rect 8200 5160 8250 5170
rect 8600 5160 8650 5170
rect 8700 5160 8750 5170
rect 8800 5160 8950 5170
rect 9000 5160 9200 5170
rect 9500 5160 9600 5170
rect 9800 5160 9950 5170
rect 2050 5150 2250 5160
rect 2350 5150 2500 5160
rect 2800 5150 2900 5160
rect 3450 5150 3500 5160
rect 7300 5150 7350 5160
rect 8000 5150 8050 5160
rect 8200 5150 8250 5160
rect 8600 5150 8650 5160
rect 8700 5150 8750 5160
rect 8800 5150 8950 5160
rect 9000 5150 9200 5160
rect 9500 5150 9600 5160
rect 9800 5150 9950 5160
rect 500 5140 600 5150
rect 2100 5140 2300 5150
rect 2400 5140 2500 5150
rect 2700 5140 2750 5150
rect 7300 5140 7350 5150
rect 8050 5140 8100 5150
rect 8450 5140 8500 5150
rect 8750 5140 8850 5150
rect 8900 5140 9050 5150
rect 9250 5140 9400 5150
rect 9500 5140 9650 5150
rect 9700 5140 9800 5150
rect 500 5130 600 5140
rect 2100 5130 2300 5140
rect 2400 5130 2500 5140
rect 2700 5130 2750 5140
rect 7300 5130 7350 5140
rect 8050 5130 8100 5140
rect 8450 5130 8500 5140
rect 8750 5130 8850 5140
rect 8900 5130 9050 5140
rect 9250 5130 9400 5140
rect 9500 5130 9650 5140
rect 9700 5130 9800 5140
rect 500 5120 600 5130
rect 2100 5120 2300 5130
rect 2400 5120 2500 5130
rect 2700 5120 2750 5130
rect 7300 5120 7350 5130
rect 8050 5120 8100 5130
rect 8450 5120 8500 5130
rect 8750 5120 8850 5130
rect 8900 5120 9050 5130
rect 9250 5120 9400 5130
rect 9500 5120 9650 5130
rect 9700 5120 9800 5130
rect 500 5110 600 5120
rect 2100 5110 2300 5120
rect 2400 5110 2500 5120
rect 2700 5110 2750 5120
rect 7300 5110 7350 5120
rect 8050 5110 8100 5120
rect 8450 5110 8500 5120
rect 8750 5110 8850 5120
rect 8900 5110 9050 5120
rect 9250 5110 9400 5120
rect 9500 5110 9650 5120
rect 9700 5110 9800 5120
rect 500 5100 600 5110
rect 2100 5100 2300 5110
rect 2400 5100 2500 5110
rect 2700 5100 2750 5110
rect 7300 5100 7350 5110
rect 8050 5100 8100 5110
rect 8450 5100 8500 5110
rect 8750 5100 8850 5110
rect 8900 5100 9050 5110
rect 9250 5100 9400 5110
rect 9500 5100 9650 5110
rect 9700 5100 9800 5110
rect 350 5090 500 5100
rect 2150 5090 2300 5100
rect 2400 5090 2500 5100
rect 2650 5090 2800 5100
rect 5150 5090 5200 5100
rect 8400 5090 8450 5100
rect 8650 5090 8700 5100
rect 9100 5090 9150 5100
rect 9300 5090 9400 5100
rect 9450 5090 9600 5100
rect 350 5080 500 5090
rect 2150 5080 2300 5090
rect 2400 5080 2500 5090
rect 2650 5080 2800 5090
rect 5150 5080 5200 5090
rect 8400 5080 8450 5090
rect 8650 5080 8700 5090
rect 9100 5080 9150 5090
rect 9300 5080 9400 5090
rect 9450 5080 9600 5090
rect 350 5070 500 5080
rect 2150 5070 2300 5080
rect 2400 5070 2500 5080
rect 2650 5070 2800 5080
rect 5150 5070 5200 5080
rect 8400 5070 8450 5080
rect 8650 5070 8700 5080
rect 9100 5070 9150 5080
rect 9300 5070 9400 5080
rect 9450 5070 9600 5080
rect 350 5060 500 5070
rect 2150 5060 2300 5070
rect 2400 5060 2500 5070
rect 2650 5060 2800 5070
rect 5150 5060 5200 5070
rect 8400 5060 8450 5070
rect 8650 5060 8700 5070
rect 9100 5060 9150 5070
rect 9300 5060 9400 5070
rect 9450 5060 9600 5070
rect 350 5050 500 5060
rect 2150 5050 2300 5060
rect 2400 5050 2500 5060
rect 2650 5050 2800 5060
rect 5150 5050 5200 5060
rect 8400 5050 8450 5060
rect 8650 5050 8700 5060
rect 9100 5050 9150 5060
rect 9300 5050 9400 5060
rect 9450 5050 9600 5060
rect 150 5040 200 5050
rect 350 5040 400 5050
rect 2200 5040 2300 5050
rect 2400 5040 2750 5050
rect 5150 5040 5200 5050
rect 7300 5040 7350 5050
rect 8000 5040 8050 5050
rect 8100 5040 8150 5050
rect 8400 5040 8450 5050
rect 8500 5040 8550 5050
rect 8950 5040 9150 5050
rect 9250 5040 9350 5050
rect 9450 5040 9500 5050
rect 9550 5040 9600 5050
rect 150 5030 200 5040
rect 350 5030 400 5040
rect 2200 5030 2300 5040
rect 2400 5030 2750 5040
rect 5150 5030 5200 5040
rect 7300 5030 7350 5040
rect 8000 5030 8050 5040
rect 8100 5030 8150 5040
rect 8400 5030 8450 5040
rect 8500 5030 8550 5040
rect 8950 5030 9150 5040
rect 9250 5030 9350 5040
rect 9450 5030 9500 5040
rect 9550 5030 9600 5040
rect 150 5020 200 5030
rect 350 5020 400 5030
rect 2200 5020 2300 5030
rect 2400 5020 2750 5030
rect 5150 5020 5200 5030
rect 7300 5020 7350 5030
rect 8000 5020 8050 5030
rect 8100 5020 8150 5030
rect 8400 5020 8450 5030
rect 8500 5020 8550 5030
rect 8950 5020 9150 5030
rect 9250 5020 9350 5030
rect 9450 5020 9500 5030
rect 9550 5020 9600 5030
rect 150 5010 200 5020
rect 350 5010 400 5020
rect 2200 5010 2300 5020
rect 2400 5010 2750 5020
rect 5150 5010 5200 5020
rect 7300 5010 7350 5020
rect 8000 5010 8050 5020
rect 8100 5010 8150 5020
rect 8400 5010 8450 5020
rect 8500 5010 8550 5020
rect 8950 5010 9150 5020
rect 9250 5010 9350 5020
rect 9450 5010 9500 5020
rect 9550 5010 9600 5020
rect 150 5000 200 5010
rect 350 5000 400 5010
rect 2200 5000 2300 5010
rect 2400 5000 2750 5010
rect 5150 5000 5200 5010
rect 7300 5000 7350 5010
rect 8000 5000 8050 5010
rect 8100 5000 8150 5010
rect 8400 5000 8450 5010
rect 8500 5000 8550 5010
rect 8950 5000 9150 5010
rect 9250 5000 9350 5010
rect 9450 5000 9500 5010
rect 9550 5000 9600 5010
rect 150 4990 400 5000
rect 2300 4990 2350 5000
rect 2450 4990 2600 5000
rect 3350 4990 3400 5000
rect 4200 4990 4350 5000
rect 5650 4990 5700 5000
rect 6350 4990 6400 5000
rect 7300 4990 7350 5000
rect 7850 4990 7950 5000
rect 8200 4990 8250 5000
rect 8450 4990 8500 5000
rect 8800 4990 8900 5000
rect 9000 4990 9100 5000
rect 9650 4990 9700 5000
rect 150 4980 400 4990
rect 2300 4980 2350 4990
rect 2450 4980 2600 4990
rect 3350 4980 3400 4990
rect 4200 4980 4350 4990
rect 5650 4980 5700 4990
rect 6350 4980 6400 4990
rect 7300 4980 7350 4990
rect 7850 4980 7950 4990
rect 8200 4980 8250 4990
rect 8450 4980 8500 4990
rect 8800 4980 8900 4990
rect 9000 4980 9100 4990
rect 9650 4980 9700 4990
rect 150 4970 400 4980
rect 2300 4970 2350 4980
rect 2450 4970 2600 4980
rect 3350 4970 3400 4980
rect 4200 4970 4350 4980
rect 5650 4970 5700 4980
rect 6350 4970 6400 4980
rect 7300 4970 7350 4980
rect 7850 4970 7950 4980
rect 8200 4970 8250 4980
rect 8450 4970 8500 4980
rect 8800 4970 8900 4980
rect 9000 4970 9100 4980
rect 9650 4970 9700 4980
rect 150 4960 400 4970
rect 2300 4960 2350 4970
rect 2450 4960 2600 4970
rect 3350 4960 3400 4970
rect 4200 4960 4350 4970
rect 5650 4960 5700 4970
rect 6350 4960 6400 4970
rect 7300 4960 7350 4970
rect 7850 4960 7950 4970
rect 8200 4960 8250 4970
rect 8450 4960 8500 4970
rect 8800 4960 8900 4970
rect 9000 4960 9100 4970
rect 9650 4960 9700 4970
rect 150 4950 400 4960
rect 2300 4950 2350 4960
rect 2450 4950 2600 4960
rect 3350 4950 3400 4960
rect 4200 4950 4350 4960
rect 5650 4950 5700 4960
rect 6350 4950 6400 4960
rect 7300 4950 7350 4960
rect 7850 4950 7950 4960
rect 8200 4950 8250 4960
rect 8450 4950 8500 4960
rect 8800 4950 8900 4960
rect 9000 4950 9100 4960
rect 9650 4950 9700 4960
rect 50 4940 200 4950
rect 2350 4940 2400 4950
rect 2450 4940 2600 4950
rect 4050 4940 4100 4950
rect 4150 4940 4200 4950
rect 4450 4940 4500 4950
rect 5550 4940 5600 4950
rect 5700 4940 5850 4950
rect 5900 4940 6000 4950
rect 6050 4940 6300 4950
rect 6450 4940 6500 4950
rect 7750 4940 7850 4950
rect 8150 4940 8200 4950
rect 8250 4940 8300 4950
rect 8500 4940 8550 4950
rect 8650 4940 8700 4950
rect 8850 4940 8900 4950
rect 9000 4940 9150 4950
rect 9500 4940 9550 4950
rect 9650 4940 9700 4950
rect 50 4930 200 4940
rect 2350 4930 2400 4940
rect 2450 4930 2600 4940
rect 4050 4930 4100 4940
rect 4150 4930 4200 4940
rect 4450 4930 4500 4940
rect 5550 4930 5600 4940
rect 5700 4930 5850 4940
rect 5900 4930 6000 4940
rect 6050 4930 6300 4940
rect 6450 4930 6500 4940
rect 7750 4930 7850 4940
rect 8150 4930 8200 4940
rect 8250 4930 8300 4940
rect 8500 4930 8550 4940
rect 8650 4930 8700 4940
rect 8850 4930 8900 4940
rect 9000 4930 9150 4940
rect 9500 4930 9550 4940
rect 9650 4930 9700 4940
rect 50 4920 200 4930
rect 2350 4920 2400 4930
rect 2450 4920 2600 4930
rect 4050 4920 4100 4930
rect 4150 4920 4200 4930
rect 4450 4920 4500 4930
rect 5550 4920 5600 4930
rect 5700 4920 5850 4930
rect 5900 4920 6000 4930
rect 6050 4920 6300 4930
rect 6450 4920 6500 4930
rect 7750 4920 7850 4930
rect 8150 4920 8200 4930
rect 8250 4920 8300 4930
rect 8500 4920 8550 4930
rect 8650 4920 8700 4930
rect 8850 4920 8900 4930
rect 9000 4920 9150 4930
rect 9500 4920 9550 4930
rect 9650 4920 9700 4930
rect 50 4910 200 4920
rect 2350 4910 2400 4920
rect 2450 4910 2600 4920
rect 4050 4910 4100 4920
rect 4150 4910 4200 4920
rect 4450 4910 4500 4920
rect 5550 4910 5600 4920
rect 5700 4910 5850 4920
rect 5900 4910 6000 4920
rect 6050 4910 6300 4920
rect 6450 4910 6500 4920
rect 7750 4910 7850 4920
rect 8150 4910 8200 4920
rect 8250 4910 8300 4920
rect 8500 4910 8550 4920
rect 8650 4910 8700 4920
rect 8850 4910 8900 4920
rect 9000 4910 9150 4920
rect 9500 4910 9550 4920
rect 9650 4910 9700 4920
rect 50 4900 200 4910
rect 2350 4900 2400 4910
rect 2450 4900 2600 4910
rect 4050 4900 4100 4910
rect 4150 4900 4200 4910
rect 4450 4900 4500 4910
rect 5550 4900 5600 4910
rect 5700 4900 5850 4910
rect 5900 4900 6000 4910
rect 6050 4900 6300 4910
rect 6450 4900 6500 4910
rect 7750 4900 7850 4910
rect 8150 4900 8200 4910
rect 8250 4900 8300 4910
rect 8500 4900 8550 4910
rect 8650 4900 8700 4910
rect 8850 4900 8900 4910
rect 9000 4900 9150 4910
rect 9500 4900 9550 4910
rect 9650 4900 9700 4910
rect 0 4890 50 4900
rect 2350 4890 2400 4900
rect 2500 4890 2650 4900
rect 3850 4890 3900 4900
rect 4000 4890 4050 4900
rect 4800 4890 4850 4900
rect 5500 4890 5550 4900
rect 5700 4890 5850 4900
rect 6450 4890 6550 4900
rect 8000 4890 8100 4900
rect 8450 4890 8500 4900
rect 8550 4890 8600 4900
rect 8900 4890 8950 4900
rect 9050 4890 9100 4900
rect 9350 4890 9450 4900
rect 9600 4890 9650 4900
rect 0 4880 50 4890
rect 2350 4880 2400 4890
rect 2500 4880 2650 4890
rect 3850 4880 3900 4890
rect 4000 4880 4050 4890
rect 4800 4880 4850 4890
rect 5500 4880 5550 4890
rect 5700 4880 5850 4890
rect 6450 4880 6550 4890
rect 8000 4880 8100 4890
rect 8450 4880 8500 4890
rect 8550 4880 8600 4890
rect 8900 4880 8950 4890
rect 9050 4880 9100 4890
rect 9350 4880 9450 4890
rect 9600 4880 9650 4890
rect 0 4870 50 4880
rect 2350 4870 2400 4880
rect 2500 4870 2650 4880
rect 3850 4870 3900 4880
rect 4000 4870 4050 4880
rect 4800 4870 4850 4880
rect 5500 4870 5550 4880
rect 5700 4870 5850 4880
rect 6450 4870 6550 4880
rect 8000 4870 8100 4880
rect 8450 4870 8500 4880
rect 8550 4870 8600 4880
rect 8900 4870 8950 4880
rect 9050 4870 9100 4880
rect 9350 4870 9450 4880
rect 9600 4870 9650 4880
rect 0 4860 50 4870
rect 2350 4860 2400 4870
rect 2500 4860 2650 4870
rect 3850 4860 3900 4870
rect 4000 4860 4050 4870
rect 4800 4860 4850 4870
rect 5500 4860 5550 4870
rect 5700 4860 5850 4870
rect 6450 4860 6550 4870
rect 8000 4860 8100 4870
rect 8450 4860 8500 4870
rect 8550 4860 8600 4870
rect 8900 4860 8950 4870
rect 9050 4860 9100 4870
rect 9350 4860 9450 4870
rect 9600 4860 9650 4870
rect 0 4850 50 4860
rect 2350 4850 2400 4860
rect 2500 4850 2650 4860
rect 3850 4850 3900 4860
rect 4000 4850 4050 4860
rect 4800 4850 4850 4860
rect 5500 4850 5550 4860
rect 5700 4850 5850 4860
rect 6450 4850 6550 4860
rect 8000 4850 8100 4860
rect 8450 4850 8500 4860
rect 8550 4850 8600 4860
rect 8900 4850 8950 4860
rect 9050 4850 9100 4860
rect 9350 4850 9450 4860
rect 9600 4850 9650 4860
rect 2350 4840 2450 4850
rect 2600 4840 2700 4850
rect 3350 4840 3400 4850
rect 4950 4840 5000 4850
rect 5450 4840 5500 4850
rect 5700 4840 5750 4850
rect 5850 4840 5950 4850
rect 6500 4840 6600 4850
rect 7800 4840 7850 4850
rect 7900 4840 7950 4850
rect 8200 4840 8300 4850
rect 8450 4840 8500 4850
rect 8550 4840 8650 4850
rect 8700 4840 8750 4850
rect 9450 4840 9500 4850
rect 9550 4840 9650 4850
rect 9700 4840 9750 4850
rect 2350 4830 2450 4840
rect 2600 4830 2700 4840
rect 3350 4830 3400 4840
rect 4950 4830 5000 4840
rect 5450 4830 5500 4840
rect 5700 4830 5750 4840
rect 5850 4830 5950 4840
rect 6500 4830 6600 4840
rect 7800 4830 7850 4840
rect 7900 4830 7950 4840
rect 8200 4830 8300 4840
rect 8450 4830 8500 4840
rect 8550 4830 8650 4840
rect 8700 4830 8750 4840
rect 9450 4830 9500 4840
rect 9550 4830 9650 4840
rect 9700 4830 9750 4840
rect 2350 4820 2450 4830
rect 2600 4820 2700 4830
rect 3350 4820 3400 4830
rect 4950 4820 5000 4830
rect 5450 4820 5500 4830
rect 5700 4820 5750 4830
rect 5850 4820 5950 4830
rect 6500 4820 6600 4830
rect 7800 4820 7850 4830
rect 7900 4820 7950 4830
rect 8200 4820 8300 4830
rect 8450 4820 8500 4830
rect 8550 4820 8650 4830
rect 8700 4820 8750 4830
rect 9450 4820 9500 4830
rect 9550 4820 9650 4830
rect 9700 4820 9750 4830
rect 2350 4810 2450 4820
rect 2600 4810 2700 4820
rect 3350 4810 3400 4820
rect 4950 4810 5000 4820
rect 5450 4810 5500 4820
rect 5700 4810 5750 4820
rect 5850 4810 5950 4820
rect 6500 4810 6600 4820
rect 7800 4810 7850 4820
rect 7900 4810 7950 4820
rect 8200 4810 8300 4820
rect 8450 4810 8500 4820
rect 8550 4810 8650 4820
rect 8700 4810 8750 4820
rect 9450 4810 9500 4820
rect 9550 4810 9650 4820
rect 9700 4810 9750 4820
rect 2350 4800 2450 4810
rect 2600 4800 2700 4810
rect 3350 4800 3400 4810
rect 4950 4800 5000 4810
rect 5450 4800 5500 4810
rect 5700 4800 5750 4810
rect 5850 4800 5950 4810
rect 6500 4800 6600 4810
rect 7800 4800 7850 4810
rect 7900 4800 7950 4810
rect 8200 4800 8300 4810
rect 8450 4800 8500 4810
rect 8550 4800 8650 4810
rect 8700 4800 8750 4810
rect 9450 4800 9500 4810
rect 9550 4800 9650 4810
rect 9700 4800 9750 4810
rect 2450 4790 2500 4800
rect 2650 4790 2750 4800
rect 5400 4790 5450 4800
rect 5650 4790 5700 4800
rect 5950 4790 6000 4800
rect 6550 4790 6650 4800
rect 8250 4790 8300 4800
rect 8500 4790 8550 4800
rect 8900 4790 9000 4800
rect 9400 4790 9500 4800
rect 2450 4780 2500 4790
rect 2650 4780 2750 4790
rect 5400 4780 5450 4790
rect 5650 4780 5700 4790
rect 5950 4780 6000 4790
rect 6550 4780 6650 4790
rect 8250 4780 8300 4790
rect 8500 4780 8550 4790
rect 8900 4780 9000 4790
rect 9400 4780 9500 4790
rect 2450 4770 2500 4780
rect 2650 4770 2750 4780
rect 5400 4770 5450 4780
rect 5650 4770 5700 4780
rect 5950 4770 6000 4780
rect 6550 4770 6650 4780
rect 8250 4770 8300 4780
rect 8500 4770 8550 4780
rect 8900 4770 9000 4780
rect 9400 4770 9500 4780
rect 2450 4760 2500 4770
rect 2650 4760 2750 4770
rect 5400 4760 5450 4770
rect 5650 4760 5700 4770
rect 5950 4760 6000 4770
rect 6550 4760 6650 4770
rect 8250 4760 8300 4770
rect 8500 4760 8550 4770
rect 8900 4760 9000 4770
rect 9400 4760 9500 4770
rect 2450 4750 2500 4760
rect 2650 4750 2750 4760
rect 5400 4750 5450 4760
rect 5650 4750 5700 4760
rect 5950 4750 6000 4760
rect 6550 4750 6650 4760
rect 8250 4750 8300 4760
rect 8500 4750 8550 4760
rect 8900 4750 9000 4760
rect 9400 4750 9500 4760
rect 0 4740 50 4750
rect 2500 4740 2750 4750
rect 3250 4740 3300 4750
rect 3500 4740 3550 4750
rect 5400 4740 5450 4750
rect 5650 4740 5700 4750
rect 6000 4740 6350 4750
rect 6600 4740 6650 4750
rect 7350 4740 7400 4750
rect 7750 4740 7800 4750
rect 7950 4740 8000 4750
rect 8250 4740 8300 4750
rect 8350 4740 8400 4750
rect 9300 4740 9350 4750
rect 0 4730 50 4740
rect 2500 4730 2750 4740
rect 3250 4730 3300 4740
rect 3500 4730 3550 4740
rect 5400 4730 5450 4740
rect 5650 4730 5700 4740
rect 6000 4730 6350 4740
rect 6600 4730 6650 4740
rect 7350 4730 7400 4740
rect 7750 4730 7800 4740
rect 7950 4730 8000 4740
rect 8250 4730 8300 4740
rect 8350 4730 8400 4740
rect 9300 4730 9350 4740
rect 0 4720 50 4730
rect 2500 4720 2750 4730
rect 3250 4720 3300 4730
rect 3500 4720 3550 4730
rect 5400 4720 5450 4730
rect 5650 4720 5700 4730
rect 6000 4720 6350 4730
rect 6600 4720 6650 4730
rect 7350 4720 7400 4730
rect 7750 4720 7800 4730
rect 7950 4720 8000 4730
rect 8250 4720 8300 4730
rect 8350 4720 8400 4730
rect 9300 4720 9350 4730
rect 0 4710 50 4720
rect 2500 4710 2750 4720
rect 3250 4710 3300 4720
rect 3500 4710 3550 4720
rect 5400 4710 5450 4720
rect 5650 4710 5700 4720
rect 6000 4710 6350 4720
rect 6600 4710 6650 4720
rect 7350 4710 7400 4720
rect 7750 4710 7800 4720
rect 7950 4710 8000 4720
rect 8250 4710 8300 4720
rect 8350 4710 8400 4720
rect 9300 4710 9350 4720
rect 0 4700 50 4710
rect 2500 4700 2750 4710
rect 3250 4700 3300 4710
rect 3500 4700 3550 4710
rect 5400 4700 5450 4710
rect 5650 4700 5700 4710
rect 6000 4700 6350 4710
rect 6600 4700 6650 4710
rect 7350 4700 7400 4710
rect 7750 4700 7800 4710
rect 7950 4700 8000 4710
rect 8250 4700 8300 4710
rect 8350 4700 8400 4710
rect 9300 4700 9350 4710
rect 5150 4690 5200 4700
rect 5350 4690 5450 4700
rect 5700 4690 5800 4700
rect 5950 4690 6350 4700
rect 6600 4690 6650 4700
rect 7600 4690 7750 4700
rect 7850 4690 7900 4700
rect 7950 4690 8000 4700
rect 8100 4690 8200 4700
rect 8500 4690 8600 4700
rect 8800 4690 8950 4700
rect 9250 4690 9300 4700
rect 5150 4680 5200 4690
rect 5350 4680 5450 4690
rect 5700 4680 5800 4690
rect 5950 4680 6350 4690
rect 6600 4680 6650 4690
rect 7600 4680 7750 4690
rect 7850 4680 7900 4690
rect 7950 4680 8000 4690
rect 8100 4680 8200 4690
rect 8500 4680 8600 4690
rect 8800 4680 8950 4690
rect 9250 4680 9300 4690
rect 5150 4670 5200 4680
rect 5350 4670 5450 4680
rect 5700 4670 5800 4680
rect 5950 4670 6350 4680
rect 6600 4670 6650 4680
rect 7600 4670 7750 4680
rect 7850 4670 7900 4680
rect 7950 4670 8000 4680
rect 8100 4670 8200 4680
rect 8500 4670 8600 4680
rect 8800 4670 8950 4680
rect 9250 4670 9300 4680
rect 5150 4660 5200 4670
rect 5350 4660 5450 4670
rect 5700 4660 5800 4670
rect 5950 4660 6350 4670
rect 6600 4660 6650 4670
rect 7600 4660 7750 4670
rect 7850 4660 7900 4670
rect 7950 4660 8000 4670
rect 8100 4660 8200 4670
rect 8500 4660 8600 4670
rect 8800 4660 8950 4670
rect 9250 4660 9300 4670
rect 5150 4650 5200 4660
rect 5350 4650 5450 4660
rect 5700 4650 5800 4660
rect 5950 4650 6350 4660
rect 6600 4650 6650 4660
rect 7600 4650 7750 4660
rect 7850 4650 7900 4660
rect 7950 4650 8000 4660
rect 8100 4650 8200 4660
rect 8500 4650 8600 4660
rect 8800 4650 8950 4660
rect 9250 4650 9300 4660
rect 3450 4640 3500 4650
rect 5350 4640 5450 4650
rect 5950 4640 6000 4650
rect 6600 4640 6650 4650
rect 7450 4640 7500 4650
rect 7650 4640 7750 4650
rect 7800 4640 7850 4650
rect 7950 4640 8000 4650
rect 8050 4640 8100 4650
rect 8250 4640 8300 4650
rect 8350 4640 8400 4650
rect 8550 4640 8650 4650
rect 8800 4640 8900 4650
rect 3450 4630 3500 4640
rect 5350 4630 5450 4640
rect 5950 4630 6000 4640
rect 6600 4630 6650 4640
rect 7450 4630 7500 4640
rect 7650 4630 7750 4640
rect 7800 4630 7850 4640
rect 7950 4630 8000 4640
rect 8050 4630 8100 4640
rect 8250 4630 8300 4640
rect 8350 4630 8400 4640
rect 8550 4630 8650 4640
rect 8800 4630 8900 4640
rect 3450 4620 3500 4630
rect 5350 4620 5450 4630
rect 5950 4620 6000 4630
rect 6600 4620 6650 4630
rect 7450 4620 7500 4630
rect 7650 4620 7750 4630
rect 7800 4620 7850 4630
rect 7950 4620 8000 4630
rect 8050 4620 8100 4630
rect 8250 4620 8300 4630
rect 8350 4620 8400 4630
rect 8550 4620 8650 4630
rect 8800 4620 8900 4630
rect 3450 4610 3500 4620
rect 5350 4610 5450 4620
rect 5950 4610 6000 4620
rect 6600 4610 6650 4620
rect 7450 4610 7500 4620
rect 7650 4610 7750 4620
rect 7800 4610 7850 4620
rect 7950 4610 8000 4620
rect 8050 4610 8100 4620
rect 8250 4610 8300 4620
rect 8350 4610 8400 4620
rect 8550 4610 8650 4620
rect 8800 4610 8900 4620
rect 3450 4600 3500 4610
rect 5350 4600 5450 4610
rect 5950 4600 6000 4610
rect 6600 4600 6650 4610
rect 7450 4600 7500 4610
rect 7650 4600 7750 4610
rect 7800 4600 7850 4610
rect 7950 4600 8000 4610
rect 8050 4600 8100 4610
rect 8250 4600 8300 4610
rect 8350 4600 8400 4610
rect 8550 4600 8650 4610
rect 8800 4600 8900 4610
rect 5200 4590 5250 4600
rect 5400 4590 5500 4600
rect 5600 4590 5650 4600
rect 6050 4590 6150 4600
rect 6550 4590 6600 4600
rect 7450 4590 7500 4600
rect 7550 4590 7600 4600
rect 7650 4590 7850 4600
rect 8100 4590 8150 4600
rect 8200 4590 8300 4600
rect 8600 4590 8650 4600
rect 5200 4580 5250 4590
rect 5400 4580 5500 4590
rect 5600 4580 5650 4590
rect 6050 4580 6150 4590
rect 6550 4580 6600 4590
rect 7450 4580 7500 4590
rect 7550 4580 7600 4590
rect 7650 4580 7850 4590
rect 8100 4580 8150 4590
rect 8200 4580 8300 4590
rect 8600 4580 8650 4590
rect 5200 4570 5250 4580
rect 5400 4570 5500 4580
rect 5600 4570 5650 4580
rect 6050 4570 6150 4580
rect 6550 4570 6600 4580
rect 7450 4570 7500 4580
rect 7550 4570 7600 4580
rect 7650 4570 7850 4580
rect 8100 4570 8150 4580
rect 8200 4570 8300 4580
rect 8600 4570 8650 4580
rect 5200 4560 5250 4570
rect 5400 4560 5500 4570
rect 5600 4560 5650 4570
rect 6050 4560 6150 4570
rect 6550 4560 6600 4570
rect 7450 4560 7500 4570
rect 7550 4560 7600 4570
rect 7650 4560 7850 4570
rect 8100 4560 8150 4570
rect 8200 4560 8300 4570
rect 8600 4560 8650 4570
rect 5200 4550 5250 4560
rect 5400 4550 5500 4560
rect 5600 4550 5650 4560
rect 6050 4550 6150 4560
rect 6550 4550 6600 4560
rect 7450 4550 7500 4560
rect 7550 4550 7600 4560
rect 7650 4550 7850 4560
rect 8100 4550 8150 4560
rect 8200 4550 8300 4560
rect 8600 4550 8650 4560
rect 3400 4540 3450 4550
rect 5250 4540 5350 4550
rect 5450 4540 5500 4550
rect 5600 4540 5700 4550
rect 5800 4540 5850 4550
rect 6200 4540 6250 4550
rect 6500 4540 6550 4550
rect 7500 4540 7550 4550
rect 7650 4540 7700 4550
rect 7950 4540 8000 4550
rect 8250 4540 8300 4550
rect 8500 4540 8550 4550
rect 9950 4540 9990 4550
rect 3400 4530 3450 4540
rect 5250 4530 5350 4540
rect 5450 4530 5500 4540
rect 5600 4530 5700 4540
rect 5800 4530 5850 4540
rect 6200 4530 6250 4540
rect 6500 4530 6550 4540
rect 7500 4530 7550 4540
rect 7650 4530 7700 4540
rect 7950 4530 8000 4540
rect 8250 4530 8300 4540
rect 8500 4530 8550 4540
rect 9950 4530 9990 4540
rect 3400 4520 3450 4530
rect 5250 4520 5350 4530
rect 5450 4520 5500 4530
rect 5600 4520 5700 4530
rect 5800 4520 5850 4530
rect 6200 4520 6250 4530
rect 6500 4520 6550 4530
rect 7500 4520 7550 4530
rect 7650 4520 7700 4530
rect 7950 4520 8000 4530
rect 8250 4520 8300 4530
rect 8500 4520 8550 4530
rect 9950 4520 9990 4530
rect 3400 4510 3450 4520
rect 5250 4510 5350 4520
rect 5450 4510 5500 4520
rect 5600 4510 5700 4520
rect 5800 4510 5850 4520
rect 6200 4510 6250 4520
rect 6500 4510 6550 4520
rect 7500 4510 7550 4520
rect 7650 4510 7700 4520
rect 7950 4510 8000 4520
rect 8250 4510 8300 4520
rect 8500 4510 8550 4520
rect 9950 4510 9990 4520
rect 3400 4500 3450 4510
rect 5250 4500 5350 4510
rect 5450 4500 5500 4510
rect 5600 4500 5700 4510
rect 5800 4500 5850 4510
rect 6200 4500 6250 4510
rect 6500 4500 6550 4510
rect 7500 4500 7550 4510
rect 7650 4500 7700 4510
rect 7950 4500 8000 4510
rect 8250 4500 8300 4510
rect 8500 4500 8550 4510
rect 9950 4500 9990 4510
rect 3000 4490 3050 4500
rect 3250 4490 3300 4500
rect 5300 4490 5600 4500
rect 5700 4490 5750 4500
rect 5800 4490 5850 4500
rect 6150 4490 6200 4500
rect 6500 4490 6550 4500
rect 7400 4490 7450 4500
rect 7750 4490 7800 4500
rect 7850 4490 7900 4500
rect 8250 4490 8350 4500
rect 9200 4490 9250 4500
rect 9900 4490 9950 4500
rect 3000 4480 3050 4490
rect 3250 4480 3300 4490
rect 5300 4480 5600 4490
rect 5700 4480 5750 4490
rect 5800 4480 5850 4490
rect 6150 4480 6200 4490
rect 6500 4480 6550 4490
rect 7400 4480 7450 4490
rect 7750 4480 7800 4490
rect 7850 4480 7900 4490
rect 8250 4480 8350 4490
rect 9200 4480 9250 4490
rect 9900 4480 9950 4490
rect 3000 4470 3050 4480
rect 3250 4470 3300 4480
rect 5300 4470 5600 4480
rect 5700 4470 5750 4480
rect 5800 4470 5850 4480
rect 6150 4470 6200 4480
rect 6500 4470 6550 4480
rect 7400 4470 7450 4480
rect 7750 4470 7800 4480
rect 7850 4470 7900 4480
rect 8250 4470 8350 4480
rect 9200 4470 9250 4480
rect 9900 4470 9950 4480
rect 3000 4460 3050 4470
rect 3250 4460 3300 4470
rect 5300 4460 5600 4470
rect 5700 4460 5750 4470
rect 5800 4460 5850 4470
rect 6150 4460 6200 4470
rect 6500 4460 6550 4470
rect 7400 4460 7450 4470
rect 7750 4460 7800 4470
rect 7850 4460 7900 4470
rect 8250 4460 8350 4470
rect 9200 4460 9250 4470
rect 9900 4460 9950 4470
rect 3000 4450 3050 4460
rect 3250 4450 3300 4460
rect 5300 4450 5600 4460
rect 5700 4450 5750 4460
rect 5800 4450 5850 4460
rect 6150 4450 6200 4460
rect 6500 4450 6550 4460
rect 7400 4450 7450 4460
rect 7750 4450 7800 4460
rect 7850 4450 7900 4460
rect 8250 4450 8350 4460
rect 9200 4450 9250 4460
rect 9900 4450 9950 4460
rect 3250 4440 3300 4450
rect 5300 4440 5600 4450
rect 5750 4440 6150 4450
rect 6500 4440 6550 4450
rect 7400 4440 7450 4450
rect 7850 4440 7900 4450
rect 8000 4440 8150 4450
rect 9850 4440 9900 4450
rect 3250 4430 3300 4440
rect 5300 4430 5600 4440
rect 5750 4430 6150 4440
rect 6500 4430 6550 4440
rect 7400 4430 7450 4440
rect 7850 4430 7900 4440
rect 8000 4430 8150 4440
rect 9850 4430 9900 4440
rect 3250 4420 3300 4430
rect 5300 4420 5600 4430
rect 5750 4420 6150 4430
rect 6500 4420 6550 4430
rect 7400 4420 7450 4430
rect 7850 4420 7900 4430
rect 8000 4420 8150 4430
rect 9850 4420 9900 4430
rect 3250 4410 3300 4420
rect 5300 4410 5600 4420
rect 5750 4410 6150 4420
rect 6500 4410 6550 4420
rect 7400 4410 7450 4420
rect 7850 4410 7900 4420
rect 8000 4410 8150 4420
rect 9850 4410 9900 4420
rect 3250 4400 3300 4410
rect 5300 4400 5600 4410
rect 5750 4400 6150 4410
rect 6500 4400 6550 4410
rect 7400 4400 7450 4410
rect 7850 4400 7900 4410
rect 8000 4400 8150 4410
rect 9850 4400 9900 4410
rect 2950 4390 3000 4400
rect 3250 4390 3350 4400
rect 4600 4390 4750 4400
rect 5300 4390 5350 4400
rect 5400 4390 5600 4400
rect 5950 4390 6050 4400
rect 6450 4390 6500 4400
rect 7400 4390 7450 4400
rect 7800 4390 7850 4400
rect 7900 4390 8000 4400
rect 8650 4390 8700 4400
rect 2950 4380 3000 4390
rect 3250 4380 3350 4390
rect 4600 4380 4750 4390
rect 5300 4380 5350 4390
rect 5400 4380 5600 4390
rect 5950 4380 6050 4390
rect 6450 4380 6500 4390
rect 7400 4380 7450 4390
rect 7800 4380 7850 4390
rect 7900 4380 8000 4390
rect 8650 4380 8700 4390
rect 2950 4370 3000 4380
rect 3250 4370 3350 4380
rect 4600 4370 4750 4380
rect 5300 4370 5350 4380
rect 5400 4370 5600 4380
rect 5950 4370 6050 4380
rect 6450 4370 6500 4380
rect 7400 4370 7450 4380
rect 7800 4370 7850 4380
rect 7900 4370 8000 4380
rect 8650 4370 8700 4380
rect 2950 4360 3000 4370
rect 3250 4360 3350 4370
rect 4600 4360 4750 4370
rect 5300 4360 5350 4370
rect 5400 4360 5600 4370
rect 5950 4360 6050 4370
rect 6450 4360 6500 4370
rect 7400 4360 7450 4370
rect 7800 4360 7850 4370
rect 7900 4360 8000 4370
rect 8650 4360 8700 4370
rect 2950 4350 3000 4360
rect 3250 4350 3350 4360
rect 4600 4350 4750 4360
rect 5300 4350 5350 4360
rect 5400 4350 5600 4360
rect 5950 4350 6050 4360
rect 6450 4350 6500 4360
rect 7400 4350 7450 4360
rect 7800 4350 7850 4360
rect 7900 4350 8000 4360
rect 8650 4350 8700 4360
rect 2950 4340 3050 4350
rect 4550 4340 4600 4350
rect 4850 4340 4900 4350
rect 5400 4340 5500 4350
rect 5950 4340 6200 4350
rect 6300 4340 6500 4350
rect 8450 4340 8750 4350
rect 2950 4330 3050 4340
rect 4550 4330 4600 4340
rect 4850 4330 4900 4340
rect 5400 4330 5500 4340
rect 5950 4330 6200 4340
rect 6300 4330 6500 4340
rect 8450 4330 8750 4340
rect 2950 4320 3050 4330
rect 4550 4320 4600 4330
rect 4850 4320 4900 4330
rect 5400 4320 5500 4330
rect 5950 4320 6200 4330
rect 6300 4320 6500 4330
rect 8450 4320 8750 4330
rect 2950 4310 3050 4320
rect 4550 4310 4600 4320
rect 4850 4310 4900 4320
rect 5400 4310 5500 4320
rect 5950 4310 6200 4320
rect 6300 4310 6500 4320
rect 8450 4310 8750 4320
rect 2950 4300 3050 4310
rect 4550 4300 4600 4310
rect 4850 4300 4900 4310
rect 5400 4300 5500 4310
rect 5950 4300 6200 4310
rect 6300 4300 6500 4310
rect 8450 4300 8750 4310
rect 3200 4290 3250 4300
rect 4200 4290 4300 4300
rect 4550 4290 4600 4300
rect 4900 4290 4950 4300
rect 5450 4290 5550 4300
rect 5950 4290 6100 4300
rect 6200 4290 6450 4300
rect 6500 4290 6600 4300
rect 7150 4290 7200 4300
rect 8500 4290 8550 4300
rect 9750 4290 9800 4300
rect 3200 4280 3250 4290
rect 4200 4280 4300 4290
rect 4550 4280 4600 4290
rect 4900 4280 4950 4290
rect 5450 4280 5550 4290
rect 5950 4280 6100 4290
rect 6200 4280 6450 4290
rect 6500 4280 6600 4290
rect 7150 4280 7200 4290
rect 8500 4280 8550 4290
rect 9750 4280 9800 4290
rect 3200 4270 3250 4280
rect 4200 4270 4300 4280
rect 4550 4270 4600 4280
rect 4900 4270 4950 4280
rect 5450 4270 5550 4280
rect 5950 4270 6100 4280
rect 6200 4270 6450 4280
rect 6500 4270 6600 4280
rect 7150 4270 7200 4280
rect 8500 4270 8550 4280
rect 9750 4270 9800 4280
rect 3200 4260 3250 4270
rect 4200 4260 4300 4270
rect 4550 4260 4600 4270
rect 4900 4260 4950 4270
rect 5450 4260 5550 4270
rect 5950 4260 6100 4270
rect 6200 4260 6450 4270
rect 6500 4260 6600 4270
rect 7150 4260 7200 4270
rect 8500 4260 8550 4270
rect 9750 4260 9800 4270
rect 3200 4250 3250 4260
rect 4200 4250 4300 4260
rect 4550 4250 4600 4260
rect 4900 4250 4950 4260
rect 5450 4250 5550 4260
rect 5950 4250 6100 4260
rect 6200 4250 6450 4260
rect 6500 4250 6600 4260
rect 7150 4250 7200 4260
rect 8500 4250 8550 4260
rect 9750 4250 9800 4260
rect 3200 4240 3250 4250
rect 4150 4240 4200 4250
rect 4300 4240 4350 4250
rect 4500 4240 4550 4250
rect 4900 4240 4950 4250
rect 5350 4240 5400 4250
rect 5500 4240 5600 4250
rect 6000 4240 6350 4250
rect 6500 4240 6600 4250
rect 7150 4240 7400 4250
rect 8800 4240 8850 4250
rect 9800 4240 9850 4250
rect 3200 4230 3250 4240
rect 4150 4230 4200 4240
rect 4300 4230 4350 4240
rect 4500 4230 4550 4240
rect 4900 4230 4950 4240
rect 5350 4230 5400 4240
rect 5500 4230 5600 4240
rect 6000 4230 6350 4240
rect 6500 4230 6600 4240
rect 7150 4230 7400 4240
rect 8800 4230 8850 4240
rect 9800 4230 9850 4240
rect 3200 4220 3250 4230
rect 4150 4220 4200 4230
rect 4300 4220 4350 4230
rect 4500 4220 4550 4230
rect 4900 4220 4950 4230
rect 5350 4220 5400 4230
rect 5500 4220 5600 4230
rect 6000 4220 6350 4230
rect 6500 4220 6600 4230
rect 7150 4220 7400 4230
rect 8800 4220 8850 4230
rect 9800 4220 9850 4230
rect 3200 4210 3250 4220
rect 4150 4210 4200 4220
rect 4300 4210 4350 4220
rect 4500 4210 4550 4220
rect 4900 4210 4950 4220
rect 5350 4210 5400 4220
rect 5500 4210 5600 4220
rect 6000 4210 6350 4220
rect 6500 4210 6600 4220
rect 7150 4210 7400 4220
rect 8800 4210 8850 4220
rect 9800 4210 9850 4220
rect 3200 4200 3250 4210
rect 4150 4200 4200 4210
rect 4300 4200 4350 4210
rect 4500 4200 4550 4210
rect 4900 4200 4950 4210
rect 5350 4200 5400 4210
rect 5500 4200 5600 4210
rect 6000 4200 6350 4210
rect 6500 4200 6600 4210
rect 7150 4200 7400 4210
rect 8800 4200 8850 4210
rect 9800 4200 9850 4210
rect 4100 4190 4150 4200
rect 4350 4190 4500 4200
rect 4650 4190 4700 4200
rect 4950 4190 5000 4200
rect 6450 4190 6600 4200
rect 7300 4190 7350 4200
rect 7450 4190 7500 4200
rect 9800 4190 9900 4200
rect 4100 4180 4150 4190
rect 4350 4180 4500 4190
rect 4650 4180 4700 4190
rect 4950 4180 5000 4190
rect 6450 4180 6600 4190
rect 7300 4180 7350 4190
rect 7450 4180 7500 4190
rect 9800 4180 9900 4190
rect 4100 4170 4150 4180
rect 4350 4170 4500 4180
rect 4650 4170 4700 4180
rect 4950 4170 5000 4180
rect 6450 4170 6600 4180
rect 7300 4170 7350 4180
rect 7450 4170 7500 4180
rect 9800 4170 9900 4180
rect 4100 4160 4150 4170
rect 4350 4160 4500 4170
rect 4650 4160 4700 4170
rect 4950 4160 5000 4170
rect 6450 4160 6600 4170
rect 7300 4160 7350 4170
rect 7450 4160 7500 4170
rect 9800 4160 9900 4170
rect 4100 4150 4150 4160
rect 4350 4150 4500 4160
rect 4650 4150 4700 4160
rect 4950 4150 5000 4160
rect 6450 4150 6600 4160
rect 7300 4150 7350 4160
rect 7450 4150 7500 4160
rect 9800 4150 9900 4160
rect 3200 4140 3300 4150
rect 4550 4140 4650 4150
rect 4900 4140 5050 4150
rect 6400 4140 6550 4150
rect 9850 4140 9990 4150
rect 3200 4130 3300 4140
rect 4550 4130 4650 4140
rect 4900 4130 5050 4140
rect 6400 4130 6550 4140
rect 9850 4130 9990 4140
rect 3200 4120 3300 4130
rect 4550 4120 4650 4130
rect 4900 4120 5050 4130
rect 6400 4120 6550 4130
rect 9850 4120 9990 4130
rect 3200 4110 3300 4120
rect 4550 4110 4650 4120
rect 4900 4110 5050 4120
rect 6400 4110 6550 4120
rect 9850 4110 9990 4120
rect 3200 4100 3300 4110
rect 4550 4100 4650 4110
rect 4900 4100 5050 4110
rect 6400 4100 6550 4110
rect 9850 4100 9990 4110
rect 3100 4090 3200 4100
rect 3250 4090 3300 4100
rect 4050 4090 4100 4100
rect 4550 4090 4600 4100
rect 4800 4090 4850 4100
rect 5050 4090 5100 4100
rect 5400 4090 5450 4100
rect 5700 4090 5750 4100
rect 6300 4090 6450 4100
rect 7200 4090 7250 4100
rect 9950 4090 9990 4100
rect 3100 4080 3200 4090
rect 3250 4080 3300 4090
rect 4050 4080 4100 4090
rect 4550 4080 4600 4090
rect 4800 4080 4850 4090
rect 5050 4080 5100 4090
rect 5400 4080 5450 4090
rect 5700 4080 5750 4090
rect 6300 4080 6450 4090
rect 7200 4080 7250 4090
rect 9950 4080 9990 4090
rect 3100 4070 3200 4080
rect 3250 4070 3300 4080
rect 4050 4070 4100 4080
rect 4550 4070 4600 4080
rect 4800 4070 4850 4080
rect 5050 4070 5100 4080
rect 5400 4070 5450 4080
rect 5700 4070 5750 4080
rect 6300 4070 6450 4080
rect 7200 4070 7250 4080
rect 9950 4070 9990 4080
rect 3100 4060 3200 4070
rect 3250 4060 3300 4070
rect 4050 4060 4100 4070
rect 4550 4060 4600 4070
rect 4800 4060 4850 4070
rect 5050 4060 5100 4070
rect 5400 4060 5450 4070
rect 5700 4060 5750 4070
rect 6300 4060 6450 4070
rect 7200 4060 7250 4070
rect 9950 4060 9990 4070
rect 3100 4050 3200 4060
rect 3250 4050 3300 4060
rect 4050 4050 4100 4060
rect 4550 4050 4600 4060
rect 4800 4050 4850 4060
rect 5050 4050 5100 4060
rect 5400 4050 5450 4060
rect 5700 4050 5750 4060
rect 6300 4050 6450 4060
rect 7200 4050 7250 4060
rect 9950 4050 9990 4060
rect 3100 4040 3200 4050
rect 3250 4040 3300 4050
rect 4550 4040 4600 4050
rect 5750 4040 6050 4050
rect 6200 4040 6400 4050
rect 8550 4040 8650 4050
rect 8750 4040 8800 4050
rect 3100 4030 3200 4040
rect 3250 4030 3300 4040
rect 4550 4030 4600 4040
rect 5750 4030 6050 4040
rect 6200 4030 6400 4040
rect 8550 4030 8650 4040
rect 8750 4030 8800 4040
rect 3100 4020 3200 4030
rect 3250 4020 3300 4030
rect 4550 4020 4600 4030
rect 5750 4020 6050 4030
rect 6200 4020 6400 4030
rect 8550 4020 8650 4030
rect 8750 4020 8800 4030
rect 3100 4010 3200 4020
rect 3250 4010 3300 4020
rect 4550 4010 4600 4020
rect 5750 4010 6050 4020
rect 6200 4010 6400 4020
rect 8550 4010 8650 4020
rect 8750 4010 8800 4020
rect 3100 4000 3200 4010
rect 3250 4000 3300 4010
rect 4550 4000 4600 4010
rect 5750 4000 6050 4010
rect 6200 4000 6400 4010
rect 8550 4000 8650 4010
rect 8750 4000 8800 4010
rect 3100 3990 3200 4000
rect 4150 3990 4300 4000
rect 4550 3990 4700 4000
rect 5100 3990 5150 4000
rect 5400 3990 5500 4000
rect 6100 3990 6150 4000
rect 6350 3990 6400 4000
rect 8250 3990 8350 4000
rect 8400 3990 8450 4000
rect 8500 3990 8550 4000
rect 8650 3990 8750 4000
rect 3100 3980 3200 3990
rect 4150 3980 4300 3990
rect 4550 3980 4700 3990
rect 5100 3980 5150 3990
rect 5400 3980 5500 3990
rect 6100 3980 6150 3990
rect 6350 3980 6400 3990
rect 8250 3980 8350 3990
rect 8400 3980 8450 3990
rect 8500 3980 8550 3990
rect 8650 3980 8750 3990
rect 3100 3970 3200 3980
rect 4150 3970 4300 3980
rect 4550 3970 4700 3980
rect 5100 3970 5150 3980
rect 5400 3970 5500 3980
rect 6100 3970 6150 3980
rect 6350 3970 6400 3980
rect 8250 3970 8350 3980
rect 8400 3970 8450 3980
rect 8500 3970 8550 3980
rect 8650 3970 8750 3980
rect 3100 3960 3200 3970
rect 4150 3960 4300 3970
rect 4550 3960 4700 3970
rect 5100 3960 5150 3970
rect 5400 3960 5500 3970
rect 6100 3960 6150 3970
rect 6350 3960 6400 3970
rect 8250 3960 8350 3970
rect 8400 3960 8450 3970
rect 8500 3960 8550 3970
rect 8650 3960 8750 3970
rect 3100 3950 3200 3960
rect 4150 3950 4300 3960
rect 4550 3950 4700 3960
rect 5100 3950 5150 3960
rect 5400 3950 5500 3960
rect 6100 3950 6150 3960
rect 6350 3950 6400 3960
rect 8250 3950 8350 3960
rect 8400 3950 8450 3960
rect 8500 3950 8550 3960
rect 8650 3950 8750 3960
rect 3150 3940 3250 3950
rect 4100 3940 4150 3950
rect 4300 3940 4350 3950
rect 5150 3940 5200 3950
rect 6350 3940 6450 3950
rect 8000 3940 8050 3950
rect 8150 3940 8200 3950
rect 8500 3940 8700 3950
rect 9650 3940 9750 3950
rect 3150 3930 3250 3940
rect 4100 3930 4150 3940
rect 4300 3930 4350 3940
rect 5150 3930 5200 3940
rect 6350 3930 6450 3940
rect 8000 3930 8050 3940
rect 8150 3930 8200 3940
rect 8500 3930 8700 3940
rect 9650 3930 9750 3940
rect 3150 3920 3250 3930
rect 4100 3920 4150 3930
rect 4300 3920 4350 3930
rect 5150 3920 5200 3930
rect 6350 3920 6450 3930
rect 8000 3920 8050 3930
rect 8150 3920 8200 3930
rect 8500 3920 8700 3930
rect 9650 3920 9750 3930
rect 3150 3910 3250 3920
rect 4100 3910 4150 3920
rect 4300 3910 4350 3920
rect 5150 3910 5200 3920
rect 6350 3910 6450 3920
rect 8000 3910 8050 3920
rect 8150 3910 8200 3920
rect 8500 3910 8700 3920
rect 9650 3910 9750 3920
rect 3150 3900 3250 3910
rect 4100 3900 4150 3910
rect 4300 3900 4350 3910
rect 5150 3900 5200 3910
rect 6350 3900 6450 3910
rect 8000 3900 8050 3910
rect 8150 3900 8200 3910
rect 8500 3900 8700 3910
rect 9650 3900 9750 3910
rect 3100 3890 3200 3900
rect 3250 3890 3300 3900
rect 4050 3890 4100 3900
rect 4300 3890 4350 3900
rect 6400 3890 6500 3900
rect 8000 3890 8050 3900
rect 8300 3890 8350 3900
rect 8550 3890 8700 3900
rect 9550 3890 9600 3900
rect 9700 3890 9750 3900
rect 3100 3880 3200 3890
rect 3250 3880 3300 3890
rect 4050 3880 4100 3890
rect 4300 3880 4350 3890
rect 6400 3880 6500 3890
rect 8000 3880 8050 3890
rect 8300 3880 8350 3890
rect 8550 3880 8700 3890
rect 9550 3880 9600 3890
rect 9700 3880 9750 3890
rect 3100 3870 3200 3880
rect 3250 3870 3300 3880
rect 4050 3870 4100 3880
rect 4300 3870 4350 3880
rect 6400 3870 6500 3880
rect 8000 3870 8050 3880
rect 8300 3870 8350 3880
rect 8550 3870 8700 3880
rect 9550 3870 9600 3880
rect 9700 3870 9750 3880
rect 3100 3860 3200 3870
rect 3250 3860 3300 3870
rect 4050 3860 4100 3870
rect 4300 3860 4350 3870
rect 6400 3860 6500 3870
rect 8000 3860 8050 3870
rect 8300 3860 8350 3870
rect 8550 3860 8700 3870
rect 9550 3860 9600 3870
rect 9700 3860 9750 3870
rect 3100 3850 3200 3860
rect 3250 3850 3300 3860
rect 4050 3850 4100 3860
rect 4300 3850 4350 3860
rect 6400 3850 6500 3860
rect 8000 3850 8050 3860
rect 8300 3850 8350 3860
rect 8550 3850 8700 3860
rect 9550 3850 9600 3860
rect 9700 3850 9750 3860
rect 3000 3840 3200 3850
rect 3250 3840 3300 3850
rect 4000 3840 4050 3850
rect 4300 3840 4350 3850
rect 5200 3840 5250 3850
rect 6400 3840 6550 3850
rect 9750 3840 9800 3850
rect 3000 3830 3200 3840
rect 3250 3830 3300 3840
rect 4000 3830 4050 3840
rect 4300 3830 4350 3840
rect 5200 3830 5250 3840
rect 6400 3830 6550 3840
rect 9750 3830 9800 3840
rect 3000 3820 3200 3830
rect 3250 3820 3300 3830
rect 4000 3820 4050 3830
rect 4300 3820 4350 3830
rect 5200 3820 5250 3830
rect 6400 3820 6550 3830
rect 9750 3820 9800 3830
rect 3000 3810 3200 3820
rect 3250 3810 3300 3820
rect 4000 3810 4050 3820
rect 4300 3810 4350 3820
rect 5200 3810 5250 3820
rect 6400 3810 6550 3820
rect 9750 3810 9800 3820
rect 3000 3800 3200 3810
rect 3250 3800 3300 3810
rect 4000 3800 4050 3810
rect 4300 3800 4350 3810
rect 5200 3800 5250 3810
rect 6400 3800 6550 3810
rect 9750 3800 9800 3810
rect 2950 3790 3100 3800
rect 3250 3790 3300 3800
rect 3900 3790 4000 3800
rect 4200 3790 4300 3800
rect 5200 3790 5250 3800
rect 6450 3790 6550 3800
rect 7050 3790 7100 3800
rect 8250 3790 8350 3800
rect 9750 3790 9850 3800
rect 2950 3780 3100 3790
rect 3250 3780 3300 3790
rect 3900 3780 4000 3790
rect 4200 3780 4300 3790
rect 5200 3780 5250 3790
rect 6450 3780 6550 3790
rect 7050 3780 7100 3790
rect 8250 3780 8350 3790
rect 9750 3780 9850 3790
rect 2950 3770 3100 3780
rect 3250 3770 3300 3780
rect 3900 3770 4000 3780
rect 4200 3770 4300 3780
rect 5200 3770 5250 3780
rect 6450 3770 6550 3780
rect 7050 3770 7100 3780
rect 8250 3770 8350 3780
rect 9750 3770 9850 3780
rect 2950 3760 3100 3770
rect 3250 3760 3300 3770
rect 3900 3760 4000 3770
rect 4200 3760 4300 3770
rect 5200 3760 5250 3770
rect 6450 3760 6550 3770
rect 7050 3760 7100 3770
rect 8250 3760 8350 3770
rect 9750 3760 9850 3770
rect 2950 3750 3100 3760
rect 3250 3750 3300 3760
rect 3900 3750 4000 3760
rect 4200 3750 4300 3760
rect 5200 3750 5250 3760
rect 6450 3750 6550 3760
rect 7050 3750 7100 3760
rect 8250 3750 8350 3760
rect 9750 3750 9850 3760
rect 2950 3740 3200 3750
rect 3250 3740 3300 3750
rect 3900 3740 3950 3750
rect 4150 3740 4250 3750
rect 4850 3740 4950 3750
rect 5250 3740 5300 3750
rect 6500 3740 6550 3750
rect 8200 3740 8450 3750
rect 8550 3740 8600 3750
rect 2950 3730 3200 3740
rect 3250 3730 3300 3740
rect 3900 3730 3950 3740
rect 4150 3730 4250 3740
rect 4850 3730 4950 3740
rect 5250 3730 5300 3740
rect 6500 3730 6550 3740
rect 8200 3730 8450 3740
rect 8550 3730 8600 3740
rect 2950 3720 3200 3730
rect 3250 3720 3300 3730
rect 3900 3720 3950 3730
rect 4150 3720 4250 3730
rect 4850 3720 4950 3730
rect 5250 3720 5300 3730
rect 6500 3720 6550 3730
rect 8200 3720 8450 3730
rect 8550 3720 8600 3730
rect 2950 3710 3200 3720
rect 3250 3710 3300 3720
rect 3900 3710 3950 3720
rect 4150 3710 4250 3720
rect 4850 3710 4950 3720
rect 5250 3710 5300 3720
rect 6500 3710 6550 3720
rect 8200 3710 8450 3720
rect 8550 3710 8600 3720
rect 2950 3700 3200 3710
rect 3250 3700 3300 3710
rect 3900 3700 3950 3710
rect 4150 3700 4250 3710
rect 4850 3700 4950 3710
rect 5250 3700 5300 3710
rect 6500 3700 6550 3710
rect 8200 3700 8450 3710
rect 8550 3700 8600 3710
rect 3100 3690 3150 3700
rect 3200 3690 3300 3700
rect 4850 3690 5100 3700
rect 5250 3690 5300 3700
rect 6500 3690 6550 3700
rect 8550 3690 8600 3700
rect 3100 3680 3150 3690
rect 3200 3680 3300 3690
rect 4850 3680 5100 3690
rect 5250 3680 5300 3690
rect 6500 3680 6550 3690
rect 8550 3680 8600 3690
rect 3100 3670 3150 3680
rect 3200 3670 3300 3680
rect 4850 3670 5100 3680
rect 5250 3670 5300 3680
rect 6500 3670 6550 3680
rect 8550 3670 8600 3680
rect 3100 3660 3150 3670
rect 3200 3660 3300 3670
rect 4850 3660 5100 3670
rect 5250 3660 5300 3670
rect 6500 3660 6550 3670
rect 8550 3660 8600 3670
rect 3100 3650 3150 3660
rect 3200 3650 3300 3660
rect 4850 3650 5100 3660
rect 5250 3650 5300 3660
rect 6500 3650 6550 3660
rect 8550 3650 8600 3660
rect 3200 3640 3300 3650
rect 3950 3640 4000 3650
rect 4950 3640 5150 3650
rect 5250 3640 5300 3650
rect 6500 3640 6550 3650
rect 8350 3640 8400 3650
rect 8500 3640 8550 3650
rect 9550 3640 9650 3650
rect 3200 3630 3300 3640
rect 3950 3630 4000 3640
rect 4950 3630 5150 3640
rect 5250 3630 5300 3640
rect 6500 3630 6550 3640
rect 8350 3630 8400 3640
rect 8500 3630 8550 3640
rect 9550 3630 9650 3640
rect 3200 3620 3300 3630
rect 3950 3620 4000 3630
rect 4950 3620 5150 3630
rect 5250 3620 5300 3630
rect 6500 3620 6550 3630
rect 8350 3620 8400 3630
rect 8500 3620 8550 3630
rect 9550 3620 9650 3630
rect 3200 3610 3300 3620
rect 3950 3610 4000 3620
rect 4950 3610 5150 3620
rect 5250 3610 5300 3620
rect 6500 3610 6550 3620
rect 8350 3610 8400 3620
rect 8500 3610 8550 3620
rect 9550 3610 9650 3620
rect 3200 3600 3300 3610
rect 3950 3600 4000 3610
rect 4950 3600 5150 3610
rect 5250 3600 5300 3610
rect 6500 3600 6550 3610
rect 8350 3600 8400 3610
rect 8500 3600 8550 3610
rect 9550 3600 9650 3610
rect 3250 3590 3350 3600
rect 3950 3590 4000 3600
rect 4750 3590 4800 3600
rect 5050 3590 5150 3600
rect 6450 3590 6550 3600
rect 6900 3590 6950 3600
rect 9400 3590 9550 3600
rect 3250 3580 3350 3590
rect 3950 3580 4000 3590
rect 4750 3580 4800 3590
rect 5050 3580 5150 3590
rect 6450 3580 6550 3590
rect 6900 3580 6950 3590
rect 9400 3580 9550 3590
rect 3250 3570 3350 3580
rect 3950 3570 4000 3580
rect 4750 3570 4800 3580
rect 5050 3570 5150 3580
rect 6450 3570 6550 3580
rect 6900 3570 6950 3580
rect 9400 3570 9550 3580
rect 3250 3560 3350 3570
rect 3950 3560 4000 3570
rect 4750 3560 4800 3570
rect 5050 3560 5150 3570
rect 6450 3560 6550 3570
rect 6900 3560 6950 3570
rect 9400 3560 9550 3570
rect 3250 3550 3350 3560
rect 3950 3550 4000 3560
rect 4750 3550 4800 3560
rect 5050 3550 5150 3560
rect 6450 3550 6550 3560
rect 6900 3550 6950 3560
rect 9400 3550 9550 3560
rect 3300 3540 3350 3550
rect 3950 3540 4000 3550
rect 4300 3540 4400 3550
rect 4650 3540 4700 3550
rect 4750 3540 4800 3550
rect 5000 3540 5150 3550
rect 6400 3540 6500 3550
rect 6850 3540 6900 3550
rect 8400 3540 8450 3550
rect 9250 3540 9300 3550
rect 9400 3540 9450 3550
rect 3300 3530 3350 3540
rect 3950 3530 4000 3540
rect 4300 3530 4400 3540
rect 4650 3530 4700 3540
rect 4750 3530 4800 3540
rect 5000 3530 5150 3540
rect 6400 3530 6500 3540
rect 6850 3530 6900 3540
rect 8400 3530 8450 3540
rect 9250 3530 9300 3540
rect 9400 3530 9450 3540
rect 3300 3520 3350 3530
rect 3950 3520 4000 3530
rect 4300 3520 4400 3530
rect 4650 3520 4700 3530
rect 4750 3520 4800 3530
rect 5000 3520 5150 3530
rect 6400 3520 6500 3530
rect 6850 3520 6900 3530
rect 8400 3520 8450 3530
rect 9250 3520 9300 3530
rect 9400 3520 9450 3530
rect 3300 3510 3350 3520
rect 3950 3510 4000 3520
rect 4300 3510 4400 3520
rect 4650 3510 4700 3520
rect 4750 3510 4800 3520
rect 5000 3510 5150 3520
rect 6400 3510 6500 3520
rect 6850 3510 6900 3520
rect 8400 3510 8450 3520
rect 9250 3510 9300 3520
rect 9400 3510 9450 3520
rect 3300 3500 3350 3510
rect 3950 3500 4000 3510
rect 4300 3500 4400 3510
rect 4650 3500 4700 3510
rect 4750 3500 4800 3510
rect 5000 3500 5150 3510
rect 6400 3500 6500 3510
rect 6850 3500 6900 3510
rect 8400 3500 8450 3510
rect 9250 3500 9300 3510
rect 9400 3500 9450 3510
rect 2350 3490 2400 3500
rect 2700 3490 2800 3500
rect 3350 3490 3400 3500
rect 3950 3490 4000 3500
rect 4250 3490 4300 3500
rect 4350 3490 4500 3500
rect 4700 3490 4750 3500
rect 6400 3490 6500 3500
rect 8400 3490 8450 3500
rect 8500 3490 8550 3500
rect 9150 3490 9200 3500
rect 9300 3490 9350 3500
rect 9550 3490 9600 3500
rect 2350 3480 2400 3490
rect 2700 3480 2800 3490
rect 3350 3480 3400 3490
rect 3950 3480 4000 3490
rect 4250 3480 4300 3490
rect 4350 3480 4500 3490
rect 4700 3480 4750 3490
rect 6400 3480 6500 3490
rect 8400 3480 8450 3490
rect 8500 3480 8550 3490
rect 9150 3480 9200 3490
rect 9300 3480 9350 3490
rect 9550 3480 9600 3490
rect 2350 3470 2400 3480
rect 2700 3470 2800 3480
rect 3350 3470 3400 3480
rect 3950 3470 4000 3480
rect 4250 3470 4300 3480
rect 4350 3470 4500 3480
rect 4700 3470 4750 3480
rect 6400 3470 6500 3480
rect 8400 3470 8450 3480
rect 8500 3470 8550 3480
rect 9150 3470 9200 3480
rect 9300 3470 9350 3480
rect 9550 3470 9600 3480
rect 2350 3460 2400 3470
rect 2700 3460 2800 3470
rect 3350 3460 3400 3470
rect 3950 3460 4000 3470
rect 4250 3460 4300 3470
rect 4350 3460 4500 3470
rect 4700 3460 4750 3470
rect 6400 3460 6500 3470
rect 8400 3460 8450 3470
rect 8500 3460 8550 3470
rect 9150 3460 9200 3470
rect 9300 3460 9350 3470
rect 9550 3460 9600 3470
rect 2350 3450 2400 3460
rect 2700 3450 2800 3460
rect 3350 3450 3400 3460
rect 3950 3450 4000 3460
rect 4250 3450 4300 3460
rect 4350 3450 4500 3460
rect 4700 3450 4750 3460
rect 6400 3450 6500 3460
rect 8400 3450 8450 3460
rect 8500 3450 8550 3460
rect 9150 3450 9200 3460
rect 9300 3450 9350 3460
rect 9550 3450 9600 3460
rect 2250 3440 2300 3450
rect 2900 3440 2950 3450
rect 4000 3440 4050 3450
rect 4250 3440 4300 3450
rect 4350 3440 4450 3450
rect 4700 3440 4800 3450
rect 4850 3440 4900 3450
rect 5000 3440 5050 3450
rect 6350 3440 6450 3450
rect 8500 3440 8550 3450
rect 9100 3440 9150 3450
rect 9200 3440 9250 3450
rect 9450 3440 9600 3450
rect 2250 3430 2300 3440
rect 2900 3430 2950 3440
rect 4000 3430 4050 3440
rect 4250 3430 4300 3440
rect 4350 3430 4450 3440
rect 4700 3430 4800 3440
rect 4850 3430 4900 3440
rect 5000 3430 5050 3440
rect 6350 3430 6450 3440
rect 8500 3430 8550 3440
rect 9100 3430 9150 3440
rect 9200 3430 9250 3440
rect 9450 3430 9600 3440
rect 2250 3420 2300 3430
rect 2900 3420 2950 3430
rect 4000 3420 4050 3430
rect 4250 3420 4300 3430
rect 4350 3420 4450 3430
rect 4700 3420 4800 3430
rect 4850 3420 4900 3430
rect 5000 3420 5050 3430
rect 6350 3420 6450 3430
rect 8500 3420 8550 3430
rect 9100 3420 9150 3430
rect 9200 3420 9250 3430
rect 9450 3420 9600 3430
rect 2250 3410 2300 3420
rect 2900 3410 2950 3420
rect 4000 3410 4050 3420
rect 4250 3410 4300 3420
rect 4350 3410 4450 3420
rect 4700 3410 4800 3420
rect 4850 3410 4900 3420
rect 5000 3410 5050 3420
rect 6350 3410 6450 3420
rect 8500 3410 8550 3420
rect 9100 3410 9150 3420
rect 9200 3410 9250 3420
rect 9450 3410 9600 3420
rect 2250 3400 2300 3410
rect 2900 3400 2950 3410
rect 4000 3400 4050 3410
rect 4250 3400 4300 3410
rect 4350 3400 4450 3410
rect 4700 3400 4800 3410
rect 4850 3400 4900 3410
rect 5000 3400 5050 3410
rect 6350 3400 6450 3410
rect 8500 3400 8550 3410
rect 9100 3400 9150 3410
rect 9200 3400 9250 3410
rect 9450 3400 9600 3410
rect 3000 3390 3050 3400
rect 4000 3390 4100 3400
rect 4200 3390 4250 3400
rect 4350 3390 4400 3400
rect 4450 3390 4700 3400
rect 4900 3390 5000 3400
rect 5250 3390 5300 3400
rect 6250 3390 6400 3400
rect 6700 3390 6750 3400
rect 8500 3390 8550 3400
rect 9050 3390 9100 3400
rect 9450 3390 9550 3400
rect 3000 3380 3050 3390
rect 4000 3380 4100 3390
rect 4200 3380 4250 3390
rect 4350 3380 4400 3390
rect 4450 3380 4700 3390
rect 4900 3380 5000 3390
rect 5250 3380 5300 3390
rect 6250 3380 6400 3390
rect 6700 3380 6750 3390
rect 8500 3380 8550 3390
rect 9050 3380 9100 3390
rect 9450 3380 9550 3390
rect 3000 3370 3050 3380
rect 4000 3370 4100 3380
rect 4200 3370 4250 3380
rect 4350 3370 4400 3380
rect 4450 3370 4700 3380
rect 4900 3370 5000 3380
rect 5250 3370 5300 3380
rect 6250 3370 6400 3380
rect 6700 3370 6750 3380
rect 8500 3370 8550 3380
rect 9050 3370 9100 3380
rect 9450 3370 9550 3380
rect 3000 3360 3050 3370
rect 4000 3360 4100 3370
rect 4200 3360 4250 3370
rect 4350 3360 4400 3370
rect 4450 3360 4700 3370
rect 4900 3360 5000 3370
rect 5250 3360 5300 3370
rect 6250 3360 6400 3370
rect 6700 3360 6750 3370
rect 8500 3360 8550 3370
rect 9050 3360 9100 3370
rect 9450 3360 9550 3370
rect 3000 3350 3050 3360
rect 4000 3350 4100 3360
rect 4200 3350 4250 3360
rect 4350 3350 4400 3360
rect 4450 3350 4700 3360
rect 4900 3350 5000 3360
rect 5250 3350 5300 3360
rect 6250 3350 6400 3360
rect 6700 3350 6750 3360
rect 8500 3350 8550 3360
rect 9050 3350 9100 3360
rect 9450 3350 9550 3360
rect 3500 3340 3600 3350
rect 4050 3340 4250 3350
rect 4550 3340 4600 3350
rect 4850 3340 4900 3350
rect 4950 3340 5000 3350
rect 5250 3340 5300 3350
rect 6200 3340 6350 3350
rect 6650 3340 6700 3350
rect 9100 3340 9150 3350
rect 9400 3340 9500 3350
rect 9650 3340 9750 3350
rect 3500 3330 3600 3340
rect 4050 3330 4250 3340
rect 4550 3330 4600 3340
rect 4850 3330 4900 3340
rect 4950 3330 5000 3340
rect 5250 3330 5300 3340
rect 6200 3330 6350 3340
rect 6650 3330 6700 3340
rect 9100 3330 9150 3340
rect 9400 3330 9500 3340
rect 9650 3330 9750 3340
rect 3500 3320 3600 3330
rect 4050 3320 4250 3330
rect 4550 3320 4600 3330
rect 4850 3320 4900 3330
rect 4950 3320 5000 3330
rect 5250 3320 5300 3330
rect 6200 3320 6350 3330
rect 6650 3320 6700 3330
rect 9100 3320 9150 3330
rect 9400 3320 9500 3330
rect 9650 3320 9750 3330
rect 3500 3310 3600 3320
rect 4050 3310 4250 3320
rect 4550 3310 4600 3320
rect 4850 3310 4900 3320
rect 4950 3310 5000 3320
rect 5250 3310 5300 3320
rect 6200 3310 6350 3320
rect 6650 3310 6700 3320
rect 9100 3310 9150 3320
rect 9400 3310 9500 3320
rect 9650 3310 9750 3320
rect 3500 3300 3600 3310
rect 4050 3300 4250 3310
rect 4550 3300 4600 3310
rect 4850 3300 4900 3310
rect 4950 3300 5000 3310
rect 5250 3300 5300 3310
rect 6200 3300 6350 3310
rect 6650 3300 6700 3310
rect 9100 3300 9150 3310
rect 9400 3300 9500 3310
rect 9650 3300 9750 3310
rect 2100 3290 2150 3300
rect 3100 3290 3150 3300
rect 4150 3290 4200 3300
rect 4350 3290 4500 3300
rect 4750 3290 4800 3300
rect 4950 3290 5000 3300
rect 5250 3290 5300 3300
rect 6200 3290 6300 3300
rect 6550 3290 6650 3300
rect 9050 3290 9100 3300
rect 9400 3290 9450 3300
rect 9600 3290 9650 3300
rect 2100 3280 2150 3290
rect 3100 3280 3150 3290
rect 4150 3280 4200 3290
rect 4350 3280 4500 3290
rect 4750 3280 4800 3290
rect 4950 3280 5000 3290
rect 5250 3280 5300 3290
rect 6200 3280 6300 3290
rect 6550 3280 6650 3290
rect 9050 3280 9100 3290
rect 9400 3280 9450 3290
rect 9600 3280 9650 3290
rect 2100 3270 2150 3280
rect 3100 3270 3150 3280
rect 4150 3270 4200 3280
rect 4350 3270 4500 3280
rect 4750 3270 4800 3280
rect 4950 3270 5000 3280
rect 5250 3270 5300 3280
rect 6200 3270 6300 3280
rect 6550 3270 6650 3280
rect 9050 3270 9100 3280
rect 9400 3270 9450 3280
rect 9600 3270 9650 3280
rect 2100 3260 2150 3270
rect 3100 3260 3150 3270
rect 4150 3260 4200 3270
rect 4350 3260 4500 3270
rect 4750 3260 4800 3270
rect 4950 3260 5000 3270
rect 5250 3260 5300 3270
rect 6200 3260 6300 3270
rect 6550 3260 6650 3270
rect 9050 3260 9100 3270
rect 9400 3260 9450 3270
rect 9600 3260 9650 3270
rect 2100 3250 2150 3260
rect 3100 3250 3150 3260
rect 4150 3250 4200 3260
rect 4350 3250 4500 3260
rect 4750 3250 4800 3260
rect 4950 3250 5000 3260
rect 5250 3250 5300 3260
rect 6200 3250 6300 3260
rect 6550 3250 6650 3260
rect 9050 3250 9100 3260
rect 9400 3250 9450 3260
rect 9600 3250 9650 3260
rect 4650 3240 4750 3250
rect 4900 3240 5000 3250
rect 5250 3240 5300 3250
rect 6250 3240 6300 3250
rect 6400 3240 6500 3250
rect 9050 3240 9100 3250
rect 9300 3240 9350 3250
rect 9400 3240 9550 3250
rect 9600 3240 9650 3250
rect 4650 3230 4750 3240
rect 4900 3230 5000 3240
rect 5250 3230 5300 3240
rect 6250 3230 6300 3240
rect 6400 3230 6500 3240
rect 9050 3230 9100 3240
rect 9300 3230 9350 3240
rect 9400 3230 9550 3240
rect 9600 3230 9650 3240
rect 4650 3220 4750 3230
rect 4900 3220 5000 3230
rect 5250 3220 5300 3230
rect 6250 3220 6300 3230
rect 6400 3220 6500 3230
rect 9050 3220 9100 3230
rect 9300 3220 9350 3230
rect 9400 3220 9550 3230
rect 9600 3220 9650 3230
rect 4650 3210 4750 3220
rect 4900 3210 5000 3220
rect 5250 3210 5300 3220
rect 6250 3210 6300 3220
rect 6400 3210 6500 3220
rect 9050 3210 9100 3220
rect 9300 3210 9350 3220
rect 9400 3210 9550 3220
rect 9600 3210 9650 3220
rect 4650 3200 4750 3210
rect 4900 3200 5000 3210
rect 5250 3200 5300 3210
rect 6250 3200 6300 3210
rect 6400 3200 6500 3210
rect 9050 3200 9100 3210
rect 9300 3200 9350 3210
rect 9400 3200 9550 3210
rect 9600 3200 9650 3210
rect 2050 3190 2100 3200
rect 3150 3190 3200 3200
rect 4200 3190 4300 3200
rect 4550 3190 4650 3200
rect 4850 3190 4900 3200
rect 6300 3190 6350 3200
rect 9000 3190 9050 3200
rect 9400 3190 9450 3200
rect 9550 3190 9600 3200
rect 2050 3180 2100 3190
rect 3150 3180 3200 3190
rect 4200 3180 4300 3190
rect 4550 3180 4650 3190
rect 4850 3180 4900 3190
rect 6300 3180 6350 3190
rect 9000 3180 9050 3190
rect 9400 3180 9450 3190
rect 9550 3180 9600 3190
rect 2050 3170 2100 3180
rect 3150 3170 3200 3180
rect 4200 3170 4300 3180
rect 4550 3170 4650 3180
rect 4850 3170 4900 3180
rect 6300 3170 6350 3180
rect 9000 3170 9050 3180
rect 9400 3170 9450 3180
rect 9550 3170 9600 3180
rect 2050 3160 2100 3170
rect 3150 3160 3200 3170
rect 4200 3160 4300 3170
rect 4550 3160 4650 3170
rect 4850 3160 4900 3170
rect 6300 3160 6350 3170
rect 9000 3160 9050 3170
rect 9400 3160 9450 3170
rect 9550 3160 9600 3170
rect 2050 3150 2100 3160
rect 3150 3150 3200 3160
rect 4200 3150 4300 3160
rect 4550 3150 4650 3160
rect 4850 3150 4900 3160
rect 6300 3150 6350 3160
rect 9000 3150 9050 3160
rect 9400 3150 9450 3160
rect 9550 3150 9600 3160
rect 2050 3140 2100 3150
rect 3150 3140 3200 3150
rect 4200 3140 4250 3150
rect 4300 3140 4350 3150
rect 4450 3140 4500 3150
rect 4550 3140 4650 3150
rect 4750 3140 4850 3150
rect 4900 3140 4950 3150
rect 8900 3140 9050 3150
rect 9850 3140 9990 3150
rect 2050 3130 2100 3140
rect 3150 3130 3200 3140
rect 4200 3130 4250 3140
rect 4300 3130 4350 3140
rect 4450 3130 4500 3140
rect 4550 3130 4650 3140
rect 4750 3130 4850 3140
rect 4900 3130 4950 3140
rect 8900 3130 9050 3140
rect 9850 3130 9990 3140
rect 2050 3120 2100 3130
rect 3150 3120 3200 3130
rect 4200 3120 4250 3130
rect 4300 3120 4350 3130
rect 4450 3120 4500 3130
rect 4550 3120 4650 3130
rect 4750 3120 4850 3130
rect 4900 3120 4950 3130
rect 8900 3120 9050 3130
rect 9850 3120 9990 3130
rect 2050 3110 2100 3120
rect 3150 3110 3200 3120
rect 4200 3110 4250 3120
rect 4300 3110 4350 3120
rect 4450 3110 4500 3120
rect 4550 3110 4650 3120
rect 4750 3110 4850 3120
rect 4900 3110 4950 3120
rect 8900 3110 9050 3120
rect 9850 3110 9990 3120
rect 2050 3100 2100 3110
rect 3150 3100 3200 3110
rect 4200 3100 4250 3110
rect 4300 3100 4350 3110
rect 4450 3100 4500 3110
rect 4550 3100 4650 3110
rect 4750 3100 4850 3110
rect 4900 3100 4950 3110
rect 8900 3100 9050 3110
rect 9850 3100 9990 3110
rect 3150 3090 3200 3100
rect 4250 3090 4300 3100
rect 4900 3090 4950 3100
rect 5200 3090 5250 3100
rect 8350 3090 8400 3100
rect 9000 3090 9050 3100
rect 9800 3090 9900 3100
rect 3150 3080 3200 3090
rect 4250 3080 4300 3090
rect 4900 3080 4950 3090
rect 5200 3080 5250 3090
rect 8350 3080 8400 3090
rect 9000 3080 9050 3090
rect 9800 3080 9900 3090
rect 3150 3070 3200 3080
rect 4250 3070 4300 3080
rect 4900 3070 4950 3080
rect 5200 3070 5250 3080
rect 8350 3070 8400 3080
rect 9000 3070 9050 3080
rect 9800 3070 9900 3080
rect 3150 3060 3200 3070
rect 4250 3060 4300 3070
rect 4900 3060 4950 3070
rect 5200 3060 5250 3070
rect 8350 3060 8400 3070
rect 9000 3060 9050 3070
rect 9800 3060 9900 3070
rect 3150 3050 3200 3060
rect 4250 3050 4300 3060
rect 4900 3050 4950 3060
rect 5200 3050 5250 3060
rect 8350 3050 8400 3060
rect 9000 3050 9050 3060
rect 9800 3050 9900 3060
rect 3850 3040 3900 3050
rect 4300 3040 4350 3050
rect 4450 3040 4550 3050
rect 4850 3040 4900 3050
rect 8900 3040 9000 3050
rect 9450 3040 9500 3050
rect 9800 3040 9900 3050
rect 3850 3030 3900 3040
rect 4300 3030 4350 3040
rect 4450 3030 4550 3040
rect 4850 3030 4900 3040
rect 8900 3030 9000 3040
rect 9450 3030 9500 3040
rect 9800 3030 9900 3040
rect 3850 3020 3900 3030
rect 4300 3020 4350 3030
rect 4450 3020 4550 3030
rect 4850 3020 4900 3030
rect 8900 3020 9000 3030
rect 9450 3020 9500 3030
rect 9800 3020 9900 3030
rect 3850 3010 3900 3020
rect 4300 3010 4350 3020
rect 4450 3010 4550 3020
rect 4850 3010 4900 3020
rect 8900 3010 9000 3020
rect 9450 3010 9500 3020
rect 9800 3010 9900 3020
rect 3850 3000 3900 3010
rect 4300 3000 4350 3010
rect 4450 3000 4550 3010
rect 4850 3000 4900 3010
rect 8900 3000 9000 3010
rect 9450 3000 9500 3010
rect 9800 3000 9900 3010
rect 4000 2990 4150 3000
rect 4350 2990 4400 3000
rect 4450 2990 4550 3000
rect 4850 2990 4950 3000
rect 5150 2990 5200 3000
rect 8400 2990 8450 3000
rect 8700 2990 8950 3000
rect 9400 2990 9450 3000
rect 4000 2980 4150 2990
rect 4350 2980 4400 2990
rect 4450 2980 4550 2990
rect 4850 2980 4950 2990
rect 5150 2980 5200 2990
rect 8400 2980 8450 2990
rect 8700 2980 8950 2990
rect 9400 2980 9450 2990
rect 4000 2970 4150 2980
rect 4350 2970 4400 2980
rect 4450 2970 4550 2980
rect 4850 2970 4950 2980
rect 5150 2970 5200 2980
rect 8400 2970 8450 2980
rect 8700 2970 8950 2980
rect 9400 2970 9450 2980
rect 4000 2960 4150 2970
rect 4350 2960 4400 2970
rect 4450 2960 4550 2970
rect 4850 2960 4950 2970
rect 5150 2960 5200 2970
rect 8400 2960 8450 2970
rect 8700 2960 8950 2970
rect 9400 2960 9450 2970
rect 4000 2950 4150 2960
rect 4350 2950 4400 2960
rect 4450 2950 4550 2960
rect 4850 2950 4950 2960
rect 5150 2950 5200 2960
rect 8400 2950 8450 2960
rect 8700 2950 8950 2960
rect 9400 2950 9450 2960
rect 2000 2940 2050 2950
rect 3900 2940 4050 2950
rect 4200 2940 4250 2950
rect 4400 2940 4550 2950
rect 4600 2940 5000 2950
rect 5100 2940 5150 2950
rect 8250 2940 8300 2950
rect 8650 2940 8900 2950
rect 9150 2940 9200 2950
rect 2000 2930 2050 2940
rect 3900 2930 4050 2940
rect 4200 2930 4250 2940
rect 4400 2930 4550 2940
rect 4600 2930 5000 2940
rect 5100 2930 5150 2940
rect 8250 2930 8300 2940
rect 8650 2930 8900 2940
rect 9150 2930 9200 2940
rect 2000 2920 2050 2930
rect 3900 2920 4050 2930
rect 4200 2920 4250 2930
rect 4400 2920 4550 2930
rect 4600 2920 5000 2930
rect 5100 2920 5150 2930
rect 8250 2920 8300 2930
rect 8650 2920 8900 2930
rect 9150 2920 9200 2930
rect 2000 2910 2050 2920
rect 3900 2910 4050 2920
rect 4200 2910 4250 2920
rect 4400 2910 4550 2920
rect 4600 2910 5000 2920
rect 5100 2910 5150 2920
rect 8250 2910 8300 2920
rect 8650 2910 8900 2920
rect 9150 2910 9200 2920
rect 2000 2900 2050 2910
rect 3900 2900 4050 2910
rect 4200 2900 4250 2910
rect 4400 2900 4550 2910
rect 4600 2900 5000 2910
rect 5100 2900 5150 2910
rect 8250 2900 8300 2910
rect 8650 2900 8900 2910
rect 9150 2900 9200 2910
rect 2000 2890 2050 2900
rect 4500 2890 4600 2900
rect 4750 2890 5100 2900
rect 7300 2890 7350 2900
rect 7400 2890 7500 2900
rect 8600 2890 8900 2900
rect 9100 2890 9200 2900
rect 9300 2890 9400 2900
rect 2000 2880 2050 2890
rect 4500 2880 4600 2890
rect 4750 2880 5100 2890
rect 7300 2880 7350 2890
rect 7400 2880 7500 2890
rect 8600 2880 8900 2890
rect 9100 2880 9200 2890
rect 9300 2880 9400 2890
rect 2000 2870 2050 2880
rect 4500 2870 4600 2880
rect 4750 2870 5100 2880
rect 7300 2870 7350 2880
rect 7400 2870 7500 2880
rect 8600 2870 8900 2880
rect 9100 2870 9200 2880
rect 9300 2870 9400 2880
rect 2000 2860 2050 2870
rect 4500 2860 4600 2870
rect 4750 2860 5100 2870
rect 7300 2860 7350 2870
rect 7400 2860 7500 2870
rect 8600 2860 8900 2870
rect 9100 2860 9200 2870
rect 9300 2860 9400 2870
rect 2000 2850 2050 2860
rect 4500 2850 4600 2860
rect 4750 2850 5100 2860
rect 7300 2850 7350 2860
rect 7400 2850 7500 2860
rect 8600 2850 8900 2860
rect 9100 2850 9200 2860
rect 9300 2850 9400 2860
rect 2000 2840 2050 2850
rect 3100 2840 3150 2850
rect 3950 2840 4000 2850
rect 4850 2840 4900 2850
rect 8600 2840 8900 2850
rect 9050 2840 9100 2850
rect 9150 2840 9400 2850
rect 2000 2830 2050 2840
rect 3100 2830 3150 2840
rect 3950 2830 4000 2840
rect 4850 2830 4900 2840
rect 8600 2830 8900 2840
rect 9050 2830 9100 2840
rect 9150 2830 9400 2840
rect 2000 2820 2050 2830
rect 3100 2820 3150 2830
rect 3950 2820 4000 2830
rect 4850 2820 4900 2830
rect 8600 2820 8900 2830
rect 9050 2820 9100 2830
rect 9150 2820 9400 2830
rect 2000 2810 2050 2820
rect 3100 2810 3150 2820
rect 3950 2810 4000 2820
rect 4850 2810 4900 2820
rect 8600 2810 8900 2820
rect 9050 2810 9100 2820
rect 9150 2810 9400 2820
rect 2000 2800 2050 2810
rect 3100 2800 3150 2810
rect 3950 2800 4000 2810
rect 4850 2800 4900 2810
rect 8600 2800 8900 2810
rect 9050 2800 9100 2810
rect 9150 2800 9400 2810
rect 2000 2790 2050 2800
rect 3100 2790 3150 2800
rect 4250 2790 4300 2800
rect 7100 2790 7150 2800
rect 7600 2790 7650 2800
rect 8150 2790 8200 2800
rect 8600 2790 8750 2800
rect 9000 2790 9300 2800
rect 9400 2790 9450 2800
rect 9650 2790 9700 2800
rect 9950 2790 9990 2800
rect 2000 2780 2050 2790
rect 3100 2780 3150 2790
rect 4250 2780 4300 2790
rect 7100 2780 7150 2790
rect 7600 2780 7650 2790
rect 8150 2780 8200 2790
rect 8600 2780 8750 2790
rect 9000 2780 9300 2790
rect 9400 2780 9450 2790
rect 9650 2780 9700 2790
rect 9950 2780 9990 2790
rect 2000 2770 2050 2780
rect 3100 2770 3150 2780
rect 4250 2770 4300 2780
rect 7100 2770 7150 2780
rect 7600 2770 7650 2780
rect 8150 2770 8200 2780
rect 8600 2770 8750 2780
rect 9000 2770 9300 2780
rect 9400 2770 9450 2780
rect 9650 2770 9700 2780
rect 9950 2770 9990 2780
rect 2000 2760 2050 2770
rect 3100 2760 3150 2770
rect 4250 2760 4300 2770
rect 7100 2760 7150 2770
rect 7600 2760 7650 2770
rect 8150 2760 8200 2770
rect 8600 2760 8750 2770
rect 9000 2760 9300 2770
rect 9400 2760 9450 2770
rect 9650 2760 9700 2770
rect 9950 2760 9990 2770
rect 2000 2750 2050 2760
rect 3100 2750 3150 2760
rect 4250 2750 4300 2760
rect 7100 2750 7150 2760
rect 7600 2750 7650 2760
rect 8150 2750 8200 2760
rect 8600 2750 8750 2760
rect 9000 2750 9300 2760
rect 9400 2750 9450 2760
rect 9650 2750 9700 2760
rect 9950 2750 9990 2760
rect 2000 2740 2050 2750
rect 3900 2740 3950 2750
rect 4250 2740 4300 2750
rect 7000 2740 7050 2750
rect 8100 2740 8150 2750
rect 8650 2740 8700 2750
rect 8950 2740 9050 2750
rect 9150 2740 9300 2750
rect 9600 2740 9700 2750
rect 9900 2740 9950 2750
rect 2000 2730 2050 2740
rect 3900 2730 3950 2740
rect 4250 2730 4300 2740
rect 7000 2730 7050 2740
rect 8100 2730 8150 2740
rect 8650 2730 8700 2740
rect 8950 2730 9050 2740
rect 9150 2730 9300 2740
rect 9600 2730 9700 2740
rect 9900 2730 9950 2740
rect 2000 2720 2050 2730
rect 3900 2720 3950 2730
rect 4250 2720 4300 2730
rect 7000 2720 7050 2730
rect 8100 2720 8150 2730
rect 8650 2720 8700 2730
rect 8950 2720 9050 2730
rect 9150 2720 9300 2730
rect 9600 2720 9700 2730
rect 9900 2720 9950 2730
rect 2000 2710 2050 2720
rect 3900 2710 3950 2720
rect 4250 2710 4300 2720
rect 7000 2710 7050 2720
rect 8100 2710 8150 2720
rect 8650 2710 8700 2720
rect 8950 2710 9050 2720
rect 9150 2710 9300 2720
rect 9600 2710 9700 2720
rect 9900 2710 9950 2720
rect 2000 2700 2050 2710
rect 3900 2700 3950 2710
rect 4250 2700 4300 2710
rect 7000 2700 7050 2710
rect 8100 2700 8150 2710
rect 8650 2700 8700 2710
rect 8950 2700 9050 2710
rect 9150 2700 9300 2710
rect 9600 2700 9700 2710
rect 9900 2700 9950 2710
rect 2200 2690 2450 2700
rect 2800 2690 3000 2700
rect 3100 2690 3150 2700
rect 4250 2690 4300 2700
rect 6000 2690 6100 2700
rect 8050 2690 8100 2700
rect 8650 2690 8900 2700
rect 9200 2690 9250 2700
rect 2200 2680 2450 2690
rect 2800 2680 3000 2690
rect 3100 2680 3150 2690
rect 4250 2680 4300 2690
rect 6000 2680 6100 2690
rect 8050 2680 8100 2690
rect 8650 2680 8900 2690
rect 9200 2680 9250 2690
rect 2200 2670 2450 2680
rect 2800 2670 3000 2680
rect 3100 2670 3150 2680
rect 4250 2670 4300 2680
rect 6000 2670 6100 2680
rect 8050 2670 8100 2680
rect 8650 2670 8900 2680
rect 9200 2670 9250 2680
rect 2200 2660 2450 2670
rect 2800 2660 3000 2670
rect 3100 2660 3150 2670
rect 4250 2660 4300 2670
rect 6000 2660 6100 2670
rect 8050 2660 8100 2670
rect 8650 2660 8900 2670
rect 9200 2660 9250 2670
rect 2200 2650 2450 2660
rect 2800 2650 3000 2660
rect 3100 2650 3150 2660
rect 4250 2650 4300 2660
rect 6000 2650 6100 2660
rect 8050 2650 8100 2660
rect 8650 2650 8900 2660
rect 9200 2650 9250 2660
rect 1950 2640 2000 2650
rect 2050 2640 2100 2650
rect 2400 2640 2450 2650
rect 2750 2640 2800 2650
rect 3000 2640 3050 2650
rect 3900 2640 3950 2650
rect 4200 2640 4300 2650
rect 5950 2640 6150 2650
rect 7700 2640 7750 2650
rect 8700 2640 8750 2650
rect 8850 2640 9000 2650
rect 9850 2640 9950 2650
rect 1950 2630 2000 2640
rect 2050 2630 2100 2640
rect 2400 2630 2450 2640
rect 2750 2630 2800 2640
rect 3000 2630 3050 2640
rect 3900 2630 3950 2640
rect 4200 2630 4300 2640
rect 5950 2630 6150 2640
rect 7700 2630 7750 2640
rect 8700 2630 8750 2640
rect 8850 2630 9000 2640
rect 9850 2630 9950 2640
rect 1950 2620 2000 2630
rect 2050 2620 2100 2630
rect 2400 2620 2450 2630
rect 2750 2620 2800 2630
rect 3000 2620 3050 2630
rect 3900 2620 3950 2630
rect 4200 2620 4300 2630
rect 5950 2620 6150 2630
rect 7700 2620 7750 2630
rect 8700 2620 8750 2630
rect 8850 2620 9000 2630
rect 9850 2620 9950 2630
rect 1950 2610 2000 2620
rect 2050 2610 2100 2620
rect 2400 2610 2450 2620
rect 2750 2610 2800 2620
rect 3000 2610 3050 2620
rect 3900 2610 3950 2620
rect 4200 2610 4300 2620
rect 5950 2610 6150 2620
rect 7700 2610 7750 2620
rect 8700 2610 8750 2620
rect 8850 2610 9000 2620
rect 9850 2610 9950 2620
rect 1950 2600 2000 2610
rect 2050 2600 2100 2610
rect 2400 2600 2450 2610
rect 2750 2600 2800 2610
rect 3000 2600 3050 2610
rect 3900 2600 3950 2610
rect 4200 2600 4300 2610
rect 5950 2600 6150 2610
rect 7700 2600 7750 2610
rect 8700 2600 8750 2610
rect 8850 2600 9000 2610
rect 9850 2600 9950 2610
rect 1950 2590 2050 2600
rect 2400 2590 2450 2600
rect 2800 2590 2850 2600
rect 3900 2590 3950 2600
rect 4200 2590 4250 2600
rect 5950 2590 6200 2600
rect 7200 2590 7300 2600
rect 7950 2590 8000 2600
rect 8850 2590 9000 2600
rect 9150 2590 9200 2600
rect 9850 2590 9900 2600
rect 1950 2580 2050 2590
rect 2400 2580 2450 2590
rect 2800 2580 2850 2590
rect 3900 2580 3950 2590
rect 4200 2580 4250 2590
rect 5950 2580 6200 2590
rect 7200 2580 7300 2590
rect 7950 2580 8000 2590
rect 8850 2580 9000 2590
rect 9150 2580 9200 2590
rect 9850 2580 9900 2590
rect 1950 2570 2050 2580
rect 2400 2570 2450 2580
rect 2800 2570 2850 2580
rect 3900 2570 3950 2580
rect 4200 2570 4250 2580
rect 5950 2570 6200 2580
rect 7200 2570 7300 2580
rect 7950 2570 8000 2580
rect 8850 2570 9000 2580
rect 9150 2570 9200 2580
rect 9850 2570 9900 2580
rect 1950 2560 2050 2570
rect 2400 2560 2450 2570
rect 2800 2560 2850 2570
rect 3900 2560 3950 2570
rect 4200 2560 4250 2570
rect 5950 2560 6200 2570
rect 7200 2560 7300 2570
rect 7950 2560 8000 2570
rect 8850 2560 9000 2570
rect 9150 2560 9200 2570
rect 9850 2560 9900 2570
rect 1950 2550 2050 2560
rect 2400 2550 2450 2560
rect 2800 2550 2850 2560
rect 3900 2550 3950 2560
rect 4200 2550 4250 2560
rect 5950 2550 6200 2560
rect 7200 2550 7300 2560
rect 7950 2550 8000 2560
rect 8850 2550 9000 2560
rect 9150 2550 9200 2560
rect 9850 2550 9900 2560
rect 1950 2540 2050 2550
rect 2100 2540 2200 2550
rect 2350 2540 2400 2550
rect 3100 2540 3200 2550
rect 3950 2540 4150 2550
rect 5850 2540 6200 2550
rect 7900 2540 7950 2550
rect 8850 2540 9050 2550
rect 9350 2540 9450 2550
rect 9550 2540 9600 2550
rect 9950 2540 9990 2550
rect 1950 2530 2050 2540
rect 2100 2530 2200 2540
rect 2350 2530 2400 2540
rect 3100 2530 3200 2540
rect 3950 2530 4150 2540
rect 5850 2530 6200 2540
rect 7900 2530 7950 2540
rect 8850 2530 9050 2540
rect 9350 2530 9450 2540
rect 9550 2530 9600 2540
rect 9950 2530 9990 2540
rect 1950 2520 2050 2530
rect 2100 2520 2200 2530
rect 2350 2520 2400 2530
rect 3100 2520 3200 2530
rect 3950 2520 4150 2530
rect 5850 2520 6200 2530
rect 7900 2520 7950 2530
rect 8850 2520 9050 2530
rect 9350 2520 9450 2530
rect 9550 2520 9600 2530
rect 9950 2520 9990 2530
rect 1950 2510 2050 2520
rect 2100 2510 2200 2520
rect 2350 2510 2400 2520
rect 3100 2510 3200 2520
rect 3950 2510 4150 2520
rect 5850 2510 6200 2520
rect 7900 2510 7950 2520
rect 8850 2510 9050 2520
rect 9350 2510 9450 2520
rect 9550 2510 9600 2520
rect 9950 2510 9990 2520
rect 1950 2500 2050 2510
rect 2100 2500 2200 2510
rect 2350 2500 2400 2510
rect 3100 2500 3200 2510
rect 3950 2500 4150 2510
rect 5850 2500 6200 2510
rect 7900 2500 7950 2510
rect 8850 2500 9050 2510
rect 9350 2500 9450 2510
rect 9550 2500 9600 2510
rect 9950 2500 9990 2510
rect 3200 2490 3250 2500
rect 5800 2490 6250 2500
rect 6750 2490 6800 2500
rect 7250 2490 7300 2500
rect 8950 2490 9150 2500
rect 9250 2490 9300 2500
rect 9650 2490 9700 2500
rect 3200 2480 3250 2490
rect 5800 2480 6250 2490
rect 6750 2480 6800 2490
rect 7250 2480 7300 2490
rect 8950 2480 9150 2490
rect 9250 2480 9300 2490
rect 9650 2480 9700 2490
rect 3200 2470 3250 2480
rect 5800 2470 6250 2480
rect 6750 2470 6800 2480
rect 7250 2470 7300 2480
rect 8950 2470 9150 2480
rect 9250 2470 9300 2480
rect 9650 2470 9700 2480
rect 3200 2460 3250 2470
rect 5800 2460 6250 2470
rect 6750 2460 6800 2470
rect 7250 2460 7300 2470
rect 8950 2460 9150 2470
rect 9250 2460 9300 2470
rect 9650 2460 9700 2470
rect 3200 2450 3250 2460
rect 5800 2450 6250 2460
rect 6750 2450 6800 2460
rect 7250 2450 7300 2460
rect 8950 2450 9150 2460
rect 9250 2450 9300 2460
rect 9650 2450 9700 2460
rect 1900 2440 1950 2450
rect 5800 2440 6300 2450
rect 6750 2440 6850 2450
rect 7300 2440 7450 2450
rect 9250 2440 9350 2450
rect 9500 2440 9550 2450
rect 9700 2440 9800 2450
rect 1900 2430 1950 2440
rect 5800 2430 6300 2440
rect 6750 2430 6850 2440
rect 7300 2430 7450 2440
rect 9250 2430 9350 2440
rect 9500 2430 9550 2440
rect 9700 2430 9800 2440
rect 1900 2420 1950 2430
rect 5800 2420 6300 2430
rect 6750 2420 6850 2430
rect 7300 2420 7450 2430
rect 9250 2420 9350 2430
rect 9500 2420 9550 2430
rect 9700 2420 9800 2430
rect 1900 2410 1950 2420
rect 5800 2410 6300 2420
rect 6750 2410 6850 2420
rect 7300 2410 7450 2420
rect 9250 2410 9350 2420
rect 9500 2410 9550 2420
rect 9700 2410 9800 2420
rect 1900 2400 1950 2410
rect 5800 2400 6300 2410
rect 6750 2400 6850 2410
rect 7300 2400 7450 2410
rect 9250 2400 9350 2410
rect 9500 2400 9550 2410
rect 9700 2400 9800 2410
rect 1900 2390 1950 2400
rect 5750 2390 6300 2400
rect 6850 2390 6950 2400
rect 7400 2390 7450 2400
rect 8400 2390 8500 2400
rect 9150 2390 9200 2400
rect 9250 2390 9400 2400
rect 9450 2390 9500 2400
rect 9550 2390 9600 2400
rect 1900 2380 1950 2390
rect 5750 2380 6300 2390
rect 6850 2380 6950 2390
rect 7400 2380 7450 2390
rect 8400 2380 8500 2390
rect 9150 2380 9200 2390
rect 9250 2380 9400 2390
rect 9450 2380 9500 2390
rect 9550 2380 9600 2390
rect 1900 2370 1950 2380
rect 5750 2370 6300 2380
rect 6850 2370 6950 2380
rect 7400 2370 7450 2380
rect 8400 2370 8500 2380
rect 9150 2370 9200 2380
rect 9250 2370 9400 2380
rect 9450 2370 9500 2380
rect 9550 2370 9600 2380
rect 1900 2360 1950 2370
rect 5750 2360 6300 2370
rect 6850 2360 6950 2370
rect 7400 2360 7450 2370
rect 8400 2360 8500 2370
rect 9150 2360 9200 2370
rect 9250 2360 9400 2370
rect 9450 2360 9500 2370
rect 9550 2360 9600 2370
rect 1900 2350 1950 2360
rect 5750 2350 6300 2360
rect 6850 2350 6950 2360
rect 7400 2350 7450 2360
rect 8400 2350 8500 2360
rect 9150 2350 9200 2360
rect 9250 2350 9400 2360
rect 9450 2350 9500 2360
rect 9550 2350 9600 2360
rect 3250 2340 3300 2350
rect 5750 2340 5900 2350
rect 6000 2340 6350 2350
rect 6950 2340 7100 2350
rect 7500 2340 7550 2350
rect 8550 2340 8600 2350
rect 9450 2340 9600 2350
rect 3250 2330 3300 2340
rect 5750 2330 5900 2340
rect 6000 2330 6350 2340
rect 6950 2330 7100 2340
rect 7500 2330 7550 2340
rect 8550 2330 8600 2340
rect 9450 2330 9600 2340
rect 3250 2320 3300 2330
rect 5750 2320 5900 2330
rect 6000 2320 6350 2330
rect 6950 2320 7100 2330
rect 7500 2320 7550 2330
rect 8550 2320 8600 2330
rect 9450 2320 9600 2330
rect 3250 2310 3300 2320
rect 5750 2310 5900 2320
rect 6000 2310 6350 2320
rect 6950 2310 7100 2320
rect 7500 2310 7550 2320
rect 8550 2310 8600 2320
rect 9450 2310 9600 2320
rect 3250 2300 3300 2310
rect 5750 2300 5900 2310
rect 6000 2300 6350 2310
rect 6950 2300 7100 2310
rect 7500 2300 7550 2310
rect 8550 2300 8600 2310
rect 9450 2300 9600 2310
rect 1850 2290 1900 2300
rect 3250 2290 3300 2300
rect 5700 2290 5900 2300
rect 6050 2290 6400 2300
rect 6750 2290 6800 2300
rect 7200 2290 7250 2300
rect 8350 2290 8400 2300
rect 8600 2290 8650 2300
rect 9100 2290 9150 2300
rect 9500 2290 9550 2300
rect 1850 2280 1900 2290
rect 3250 2280 3300 2290
rect 5700 2280 5900 2290
rect 6050 2280 6400 2290
rect 6750 2280 6800 2290
rect 7200 2280 7250 2290
rect 8350 2280 8400 2290
rect 8600 2280 8650 2290
rect 9100 2280 9150 2290
rect 9500 2280 9550 2290
rect 1850 2270 1900 2280
rect 3250 2270 3300 2280
rect 5700 2270 5900 2280
rect 6050 2270 6400 2280
rect 6750 2270 6800 2280
rect 7200 2270 7250 2280
rect 8350 2270 8400 2280
rect 8600 2270 8650 2280
rect 9100 2270 9150 2280
rect 9500 2270 9550 2280
rect 1850 2260 1900 2270
rect 3250 2260 3300 2270
rect 5700 2260 5900 2270
rect 6050 2260 6400 2270
rect 6750 2260 6800 2270
rect 7200 2260 7250 2270
rect 8350 2260 8400 2270
rect 8600 2260 8650 2270
rect 9100 2260 9150 2270
rect 9500 2260 9550 2270
rect 1850 2250 1900 2260
rect 3250 2250 3300 2260
rect 5700 2250 5900 2260
rect 6050 2250 6400 2260
rect 6750 2250 6800 2260
rect 7200 2250 7250 2260
rect 8350 2250 8400 2260
rect 8600 2250 8650 2260
rect 9100 2250 9150 2260
rect 9500 2250 9550 2260
rect 1850 2240 1900 2250
rect 3250 2240 3300 2250
rect 5700 2240 6450 2250
rect 6750 2240 6800 2250
rect 7350 2240 7400 2250
rect 8350 2240 8400 2250
rect 8800 2240 8850 2250
rect 9000 2240 9050 2250
rect 9300 2240 9400 2250
rect 9750 2240 9800 2250
rect 1850 2230 1900 2240
rect 3250 2230 3300 2240
rect 5700 2230 6450 2240
rect 6750 2230 6800 2240
rect 7350 2230 7400 2240
rect 8350 2230 8400 2240
rect 8800 2230 8850 2240
rect 9000 2230 9050 2240
rect 9300 2230 9400 2240
rect 9750 2230 9800 2240
rect 1850 2220 1900 2230
rect 3250 2220 3300 2230
rect 5700 2220 6450 2230
rect 6750 2220 6800 2230
rect 7350 2220 7400 2230
rect 8350 2220 8400 2230
rect 8800 2220 8850 2230
rect 9000 2220 9050 2230
rect 9300 2220 9400 2230
rect 9750 2220 9800 2230
rect 1850 2210 1900 2220
rect 3250 2210 3300 2220
rect 5700 2210 6450 2220
rect 6750 2210 6800 2220
rect 7350 2210 7400 2220
rect 8350 2210 8400 2220
rect 8800 2210 8850 2220
rect 9000 2210 9050 2220
rect 9300 2210 9400 2220
rect 9750 2210 9800 2220
rect 1850 2200 1900 2210
rect 3250 2200 3300 2210
rect 5700 2200 6450 2210
rect 6750 2200 6800 2210
rect 7350 2200 7400 2210
rect 8350 2200 8400 2210
rect 8800 2200 8850 2210
rect 9000 2200 9050 2210
rect 9300 2200 9400 2210
rect 9750 2200 9800 2210
rect 1850 2190 1900 2200
rect 2450 2190 2650 2200
rect 2750 2190 2800 2200
rect 3250 2190 3300 2200
rect 5650 2190 6400 2200
rect 6450 2190 6500 2200
rect 6750 2190 6900 2200
rect 7400 2190 7500 2200
rect 7700 2190 7750 2200
rect 8350 2190 8400 2200
rect 9450 2190 9500 2200
rect 9750 2190 9800 2200
rect 1850 2180 1900 2190
rect 2450 2180 2650 2190
rect 2750 2180 2800 2190
rect 3250 2180 3300 2190
rect 5650 2180 6400 2190
rect 6450 2180 6500 2190
rect 6750 2180 6900 2190
rect 7400 2180 7500 2190
rect 7700 2180 7750 2190
rect 8350 2180 8400 2190
rect 9450 2180 9500 2190
rect 9750 2180 9800 2190
rect 1850 2170 1900 2180
rect 2450 2170 2650 2180
rect 2750 2170 2800 2180
rect 3250 2170 3300 2180
rect 5650 2170 6400 2180
rect 6450 2170 6500 2180
rect 6750 2170 6900 2180
rect 7400 2170 7500 2180
rect 7700 2170 7750 2180
rect 8350 2170 8400 2180
rect 9450 2170 9500 2180
rect 9750 2170 9800 2180
rect 1850 2160 1900 2170
rect 2450 2160 2650 2170
rect 2750 2160 2800 2170
rect 3250 2160 3300 2170
rect 5650 2160 6400 2170
rect 6450 2160 6500 2170
rect 6750 2160 6900 2170
rect 7400 2160 7500 2170
rect 7700 2160 7750 2170
rect 8350 2160 8400 2170
rect 9450 2160 9500 2170
rect 9750 2160 9800 2170
rect 1850 2150 1900 2160
rect 2450 2150 2650 2160
rect 2750 2150 2800 2160
rect 3250 2150 3300 2160
rect 5650 2150 6400 2160
rect 6450 2150 6500 2160
rect 6750 2150 6900 2160
rect 7400 2150 7500 2160
rect 7700 2150 7750 2160
rect 8350 2150 8400 2160
rect 9450 2150 9500 2160
rect 9750 2150 9800 2160
rect 1850 2140 1900 2150
rect 2400 2140 2700 2150
rect 3250 2140 3300 2150
rect 5550 2140 6100 2150
rect 6200 2140 6400 2150
rect 6450 2140 6500 2150
rect 6750 2140 6950 2150
rect 7800 2140 7850 2150
rect 9250 2140 9300 2150
rect 9500 2140 9650 2150
rect 1850 2130 1900 2140
rect 2400 2130 2700 2140
rect 3250 2130 3300 2140
rect 5550 2130 6100 2140
rect 6200 2130 6400 2140
rect 6450 2130 6500 2140
rect 6750 2130 6950 2140
rect 7800 2130 7850 2140
rect 9250 2130 9300 2140
rect 9500 2130 9650 2140
rect 1850 2120 1900 2130
rect 2400 2120 2700 2130
rect 3250 2120 3300 2130
rect 5550 2120 6100 2130
rect 6200 2120 6400 2130
rect 6450 2120 6500 2130
rect 6750 2120 6950 2130
rect 7800 2120 7850 2130
rect 9250 2120 9300 2130
rect 9500 2120 9650 2130
rect 1850 2110 1900 2120
rect 2400 2110 2700 2120
rect 3250 2110 3300 2120
rect 5550 2110 6100 2120
rect 6200 2110 6400 2120
rect 6450 2110 6500 2120
rect 6750 2110 6950 2120
rect 7800 2110 7850 2120
rect 9250 2110 9300 2120
rect 9500 2110 9650 2120
rect 1850 2100 1900 2110
rect 2400 2100 2700 2110
rect 3250 2100 3300 2110
rect 5550 2100 6100 2110
rect 6200 2100 6400 2110
rect 6450 2100 6500 2110
rect 6750 2100 6950 2110
rect 7800 2100 7850 2110
rect 9250 2100 9300 2110
rect 9500 2100 9650 2110
rect 1850 2090 1900 2100
rect 3250 2090 3300 2100
rect 5350 2090 6100 2100
rect 6200 2090 6400 2100
rect 6450 2090 6500 2100
rect 6900 2090 7000 2100
rect 7850 2090 7900 2100
rect 9200 2090 9250 2100
rect 9300 2090 9600 2100
rect 9650 2090 9700 2100
rect 1850 2080 1900 2090
rect 3250 2080 3300 2090
rect 5350 2080 6100 2090
rect 6200 2080 6400 2090
rect 6450 2080 6500 2090
rect 6900 2080 7000 2090
rect 7850 2080 7900 2090
rect 9200 2080 9250 2090
rect 9300 2080 9600 2090
rect 9650 2080 9700 2090
rect 1850 2070 1900 2080
rect 3250 2070 3300 2080
rect 5350 2070 6100 2080
rect 6200 2070 6400 2080
rect 6450 2070 6500 2080
rect 6900 2070 7000 2080
rect 7850 2070 7900 2080
rect 9200 2070 9250 2080
rect 9300 2070 9600 2080
rect 9650 2070 9700 2080
rect 1850 2060 1900 2070
rect 3250 2060 3300 2070
rect 5350 2060 6100 2070
rect 6200 2060 6400 2070
rect 6450 2060 6500 2070
rect 6900 2060 7000 2070
rect 7850 2060 7900 2070
rect 9200 2060 9250 2070
rect 9300 2060 9600 2070
rect 9650 2060 9700 2070
rect 1850 2050 1900 2060
rect 3250 2050 3300 2060
rect 5350 2050 6100 2060
rect 6200 2050 6400 2060
rect 6450 2050 6500 2060
rect 6900 2050 7000 2060
rect 7850 2050 7900 2060
rect 9200 2050 9250 2060
rect 9300 2050 9600 2060
rect 9650 2050 9700 2060
rect 1850 2040 1900 2050
rect 3200 2040 3250 2050
rect 5300 2040 6100 2050
rect 6300 2040 6400 2050
rect 6450 2040 6500 2050
rect 6800 2040 6850 2050
rect 6950 2040 7050 2050
rect 7250 2040 7350 2050
rect 7950 2040 8000 2050
rect 8400 2040 8550 2050
rect 9100 2040 9450 2050
rect 1850 2030 1900 2040
rect 3200 2030 3250 2040
rect 5300 2030 6100 2040
rect 6300 2030 6400 2040
rect 6450 2030 6500 2040
rect 6800 2030 6850 2040
rect 6950 2030 7050 2040
rect 7250 2030 7350 2040
rect 7950 2030 8000 2040
rect 8400 2030 8550 2040
rect 9100 2030 9450 2040
rect 1850 2020 1900 2030
rect 3200 2020 3250 2030
rect 5300 2020 6100 2030
rect 6300 2020 6400 2030
rect 6450 2020 6500 2030
rect 6800 2020 6850 2030
rect 6950 2020 7050 2030
rect 7250 2020 7350 2030
rect 7950 2020 8000 2030
rect 8400 2020 8550 2030
rect 9100 2020 9450 2030
rect 1850 2010 1900 2020
rect 3200 2010 3250 2020
rect 5300 2010 6100 2020
rect 6300 2010 6400 2020
rect 6450 2010 6500 2020
rect 6800 2010 6850 2020
rect 6950 2010 7050 2020
rect 7250 2010 7350 2020
rect 7950 2010 8000 2020
rect 8400 2010 8550 2020
rect 9100 2010 9450 2020
rect 1850 2000 1900 2010
rect 3200 2000 3250 2010
rect 5300 2000 6100 2010
rect 6300 2000 6400 2010
rect 6450 2000 6500 2010
rect 6800 2000 6850 2010
rect 6950 2000 7050 2010
rect 7250 2000 7350 2010
rect 7950 2000 8000 2010
rect 8400 2000 8550 2010
rect 9100 2000 9450 2010
rect 1850 1990 1900 2000
rect 3200 1990 3250 2000
rect 5250 1990 6100 2000
rect 6350 1990 6400 2000
rect 6450 1990 6500 2000
rect 6800 1990 6850 2000
rect 7050 1990 7350 2000
rect 8400 1990 8450 2000
rect 8550 1990 8600 2000
rect 1850 1980 1900 1990
rect 3200 1980 3250 1990
rect 5250 1980 6100 1990
rect 6350 1980 6400 1990
rect 6450 1980 6500 1990
rect 6800 1980 6850 1990
rect 7050 1980 7350 1990
rect 8400 1980 8450 1990
rect 8550 1980 8600 1990
rect 1850 1970 1900 1980
rect 3200 1970 3250 1980
rect 5250 1970 6100 1980
rect 6350 1970 6400 1980
rect 6450 1970 6500 1980
rect 6800 1970 6850 1980
rect 7050 1970 7350 1980
rect 8400 1970 8450 1980
rect 8550 1970 8600 1980
rect 1850 1960 1900 1970
rect 3200 1960 3250 1970
rect 5250 1960 6100 1970
rect 6350 1960 6400 1970
rect 6450 1960 6500 1970
rect 6800 1960 6850 1970
rect 7050 1960 7350 1970
rect 8400 1960 8450 1970
rect 8550 1960 8600 1970
rect 1850 1950 1900 1960
rect 3200 1950 3250 1960
rect 5250 1950 6100 1960
rect 6350 1950 6400 1960
rect 6450 1950 6500 1960
rect 6800 1950 6850 1960
rect 7050 1950 7350 1960
rect 8400 1950 8450 1960
rect 8550 1950 8600 1960
rect 1850 1940 1900 1950
rect 3200 1940 3300 1950
rect 4500 1940 4550 1950
rect 4750 1940 4850 1950
rect 5000 1940 6100 1950
rect 6350 1940 6500 1950
rect 6800 1940 6850 1950
rect 7300 1940 7350 1950
rect 7800 1940 7850 1950
rect 8400 1940 8450 1950
rect 1850 1930 1900 1940
rect 3200 1930 3300 1940
rect 4500 1930 4550 1940
rect 4750 1930 4850 1940
rect 5000 1930 6100 1940
rect 6350 1930 6500 1940
rect 6800 1930 6850 1940
rect 7300 1930 7350 1940
rect 7800 1930 7850 1940
rect 8400 1930 8450 1940
rect 1850 1920 1900 1930
rect 3200 1920 3300 1930
rect 4500 1920 4550 1930
rect 4750 1920 4850 1930
rect 5000 1920 6100 1930
rect 6350 1920 6500 1930
rect 6800 1920 6850 1930
rect 7300 1920 7350 1930
rect 7800 1920 7850 1930
rect 8400 1920 8450 1930
rect 1850 1910 1900 1920
rect 3200 1910 3300 1920
rect 4500 1910 4550 1920
rect 4750 1910 4850 1920
rect 5000 1910 6100 1920
rect 6350 1910 6500 1920
rect 6800 1910 6850 1920
rect 7300 1910 7350 1920
rect 7800 1910 7850 1920
rect 8400 1910 8450 1920
rect 1850 1900 1900 1910
rect 3200 1900 3300 1910
rect 4500 1900 4550 1910
rect 4750 1900 4850 1910
rect 5000 1900 6100 1910
rect 6350 1900 6500 1910
rect 6800 1900 6850 1910
rect 7300 1900 7350 1910
rect 7800 1900 7850 1910
rect 8400 1900 8450 1910
rect 1850 1890 1900 1900
rect 2400 1890 2500 1900
rect 2750 1890 2850 1900
rect 3250 1890 3300 1900
rect 4450 1890 4500 1900
rect 4750 1890 4800 1900
rect 4850 1890 4900 1900
rect 4950 1890 6050 1900
rect 6400 1890 6450 1900
rect 6800 1890 6850 1900
rect 7300 1890 7350 1900
rect 7800 1890 7850 1900
rect 8400 1890 8450 1900
rect 9700 1890 9750 1900
rect 1850 1880 1900 1890
rect 2400 1880 2500 1890
rect 2750 1880 2850 1890
rect 3250 1880 3300 1890
rect 4450 1880 4500 1890
rect 4750 1880 4800 1890
rect 4850 1880 4900 1890
rect 4950 1880 6050 1890
rect 6400 1880 6450 1890
rect 6800 1880 6850 1890
rect 7300 1880 7350 1890
rect 7800 1880 7850 1890
rect 8400 1880 8450 1890
rect 9700 1880 9750 1890
rect 1850 1870 1900 1880
rect 2400 1870 2500 1880
rect 2750 1870 2850 1880
rect 3250 1870 3300 1880
rect 4450 1870 4500 1880
rect 4750 1870 4800 1880
rect 4850 1870 4900 1880
rect 4950 1870 6050 1880
rect 6400 1870 6450 1880
rect 6800 1870 6850 1880
rect 7300 1870 7350 1880
rect 7800 1870 7850 1880
rect 8400 1870 8450 1880
rect 9700 1870 9750 1880
rect 1850 1860 1900 1870
rect 2400 1860 2500 1870
rect 2750 1860 2850 1870
rect 3250 1860 3300 1870
rect 4450 1860 4500 1870
rect 4750 1860 4800 1870
rect 4850 1860 4900 1870
rect 4950 1860 6050 1870
rect 6400 1860 6450 1870
rect 6800 1860 6850 1870
rect 7300 1860 7350 1870
rect 7800 1860 7850 1870
rect 8400 1860 8450 1870
rect 9700 1860 9750 1870
rect 1850 1850 1900 1860
rect 2400 1850 2500 1860
rect 2750 1850 2850 1860
rect 3250 1850 3300 1860
rect 4450 1850 4500 1860
rect 4750 1850 4800 1860
rect 4850 1850 4900 1860
rect 4950 1850 6050 1860
rect 6400 1850 6450 1860
rect 6800 1850 6850 1860
rect 7300 1850 7350 1860
rect 7800 1850 7850 1860
rect 8400 1850 8450 1860
rect 9700 1850 9750 1860
rect 1850 1840 1900 1850
rect 2300 1840 2350 1850
rect 2850 1840 2900 1850
rect 3250 1840 3300 1850
rect 4450 1840 4500 1850
rect 4550 1840 4650 1850
rect 4750 1840 4900 1850
rect 4950 1840 6000 1850
rect 6350 1840 6450 1850
rect 6800 1840 6850 1850
rect 7300 1840 7350 1850
rect 7800 1840 7850 1850
rect 8350 1840 8500 1850
rect 9100 1840 9150 1850
rect 9700 1840 9750 1850
rect 9950 1840 9990 1850
rect 1850 1830 1900 1840
rect 2300 1830 2350 1840
rect 2850 1830 2900 1840
rect 3250 1830 3300 1840
rect 4450 1830 4500 1840
rect 4550 1830 4650 1840
rect 4750 1830 4900 1840
rect 4950 1830 6000 1840
rect 6350 1830 6450 1840
rect 6800 1830 6850 1840
rect 7300 1830 7350 1840
rect 7800 1830 7850 1840
rect 8350 1830 8500 1840
rect 9100 1830 9150 1840
rect 9700 1830 9750 1840
rect 9950 1830 9990 1840
rect 1850 1820 1900 1830
rect 2300 1820 2350 1830
rect 2850 1820 2900 1830
rect 3250 1820 3300 1830
rect 4450 1820 4500 1830
rect 4550 1820 4650 1830
rect 4750 1820 4900 1830
rect 4950 1820 6000 1830
rect 6350 1820 6450 1830
rect 6800 1820 6850 1830
rect 7300 1820 7350 1830
rect 7800 1820 7850 1830
rect 8350 1820 8500 1830
rect 9100 1820 9150 1830
rect 9700 1820 9750 1830
rect 9950 1820 9990 1830
rect 1850 1810 1900 1820
rect 2300 1810 2350 1820
rect 2850 1810 2900 1820
rect 3250 1810 3300 1820
rect 4450 1810 4500 1820
rect 4550 1810 4650 1820
rect 4750 1810 4900 1820
rect 4950 1810 6000 1820
rect 6350 1810 6450 1820
rect 6800 1810 6850 1820
rect 7300 1810 7350 1820
rect 7800 1810 7850 1820
rect 8350 1810 8500 1820
rect 9100 1810 9150 1820
rect 9700 1810 9750 1820
rect 9950 1810 9990 1820
rect 1850 1800 1900 1810
rect 2300 1800 2350 1810
rect 2850 1800 2900 1810
rect 3250 1800 3300 1810
rect 4450 1800 4500 1810
rect 4550 1800 4650 1810
rect 4750 1800 4900 1810
rect 4950 1800 6000 1810
rect 6350 1800 6450 1810
rect 6800 1800 6850 1810
rect 7300 1800 7350 1810
rect 7800 1800 7850 1810
rect 8350 1800 8500 1810
rect 9100 1800 9150 1810
rect 9700 1800 9750 1810
rect 9950 1800 9990 1810
rect 2350 1790 2450 1800
rect 2500 1790 2750 1800
rect 3250 1790 3300 1800
rect 4050 1790 4100 1800
rect 4450 1790 4500 1800
rect 4700 1790 4900 1800
rect 4950 1790 5200 1800
rect 5250 1790 5950 1800
rect 6350 1790 6450 1800
rect 6800 1790 6850 1800
rect 7300 1790 7350 1800
rect 7850 1790 7900 1800
rect 8350 1790 8400 1800
rect 8450 1790 8500 1800
rect 9700 1790 9750 1800
rect 2350 1780 2450 1790
rect 2500 1780 2750 1790
rect 3250 1780 3300 1790
rect 4050 1780 4100 1790
rect 4450 1780 4500 1790
rect 4700 1780 4900 1790
rect 4950 1780 5200 1790
rect 5250 1780 5950 1790
rect 6350 1780 6450 1790
rect 6800 1780 6850 1790
rect 7300 1780 7350 1790
rect 7850 1780 7900 1790
rect 8350 1780 8400 1790
rect 8450 1780 8500 1790
rect 9700 1780 9750 1790
rect 2350 1770 2450 1780
rect 2500 1770 2750 1780
rect 3250 1770 3300 1780
rect 4050 1770 4100 1780
rect 4450 1770 4500 1780
rect 4700 1770 4900 1780
rect 4950 1770 5200 1780
rect 5250 1770 5950 1780
rect 6350 1770 6450 1780
rect 6800 1770 6850 1780
rect 7300 1770 7350 1780
rect 7850 1770 7900 1780
rect 8350 1770 8400 1780
rect 8450 1770 8500 1780
rect 9700 1770 9750 1780
rect 2350 1760 2450 1770
rect 2500 1760 2750 1770
rect 3250 1760 3300 1770
rect 4050 1760 4100 1770
rect 4450 1760 4500 1770
rect 4700 1760 4900 1770
rect 4950 1760 5200 1770
rect 5250 1760 5950 1770
rect 6350 1760 6450 1770
rect 6800 1760 6850 1770
rect 7300 1760 7350 1770
rect 7850 1760 7900 1770
rect 8350 1760 8400 1770
rect 8450 1760 8500 1770
rect 9700 1760 9750 1770
rect 2350 1750 2450 1760
rect 2500 1750 2750 1760
rect 3250 1750 3300 1760
rect 4050 1750 4100 1760
rect 4450 1750 4500 1760
rect 4700 1750 4900 1760
rect 4950 1750 5200 1760
rect 5250 1750 5950 1760
rect 6350 1750 6450 1760
rect 6800 1750 6850 1760
rect 7300 1750 7350 1760
rect 7850 1750 7900 1760
rect 8350 1750 8400 1760
rect 8450 1750 8500 1760
rect 9700 1750 9750 1760
rect 1900 1740 1950 1750
rect 3200 1740 3250 1750
rect 4050 1740 4100 1750
rect 4200 1740 4250 1750
rect 4450 1740 4650 1750
rect 4700 1740 5150 1750
rect 5200 1740 5250 1750
rect 5300 1740 5950 1750
rect 6350 1740 6450 1750
rect 7300 1740 7350 1750
rect 7850 1740 7900 1750
rect 8350 1740 8400 1750
rect 8450 1740 8500 1750
rect 9100 1740 9150 1750
rect 9700 1740 9800 1750
rect 1900 1730 1950 1740
rect 3200 1730 3250 1740
rect 4050 1730 4100 1740
rect 4200 1730 4250 1740
rect 4450 1730 4650 1740
rect 4700 1730 5150 1740
rect 5200 1730 5250 1740
rect 5300 1730 5950 1740
rect 6350 1730 6450 1740
rect 7300 1730 7350 1740
rect 7850 1730 7900 1740
rect 8350 1730 8400 1740
rect 8450 1730 8500 1740
rect 9100 1730 9150 1740
rect 9700 1730 9800 1740
rect 1900 1720 1950 1730
rect 3200 1720 3250 1730
rect 4050 1720 4100 1730
rect 4200 1720 4250 1730
rect 4450 1720 4650 1730
rect 4700 1720 5150 1730
rect 5200 1720 5250 1730
rect 5300 1720 5950 1730
rect 6350 1720 6450 1730
rect 7300 1720 7350 1730
rect 7850 1720 7900 1730
rect 8350 1720 8400 1730
rect 8450 1720 8500 1730
rect 9100 1720 9150 1730
rect 9700 1720 9800 1730
rect 1900 1710 1950 1720
rect 3200 1710 3250 1720
rect 4050 1710 4100 1720
rect 4200 1710 4250 1720
rect 4450 1710 4650 1720
rect 4700 1710 5150 1720
rect 5200 1710 5250 1720
rect 5300 1710 5950 1720
rect 6350 1710 6450 1720
rect 7300 1710 7350 1720
rect 7850 1710 7900 1720
rect 8350 1710 8400 1720
rect 8450 1710 8500 1720
rect 9100 1710 9150 1720
rect 9700 1710 9800 1720
rect 1900 1700 1950 1710
rect 3200 1700 3250 1710
rect 4050 1700 4100 1710
rect 4200 1700 4250 1710
rect 4450 1700 4650 1710
rect 4700 1700 5150 1710
rect 5200 1700 5250 1710
rect 5300 1700 5950 1710
rect 6350 1700 6450 1710
rect 7300 1700 7350 1710
rect 7850 1700 7900 1710
rect 8350 1700 8400 1710
rect 8450 1700 8500 1710
rect 9100 1700 9150 1710
rect 9700 1700 9800 1710
rect 1900 1690 1950 1700
rect 3200 1690 3250 1700
rect 4050 1690 4100 1700
rect 4150 1690 4250 1700
rect 4450 1690 4500 1700
rect 4600 1690 5900 1700
rect 6400 1690 6450 1700
rect 7300 1690 7350 1700
rect 7850 1690 7900 1700
rect 8450 1690 8550 1700
rect 9100 1690 9150 1700
rect 1900 1680 1950 1690
rect 3200 1680 3250 1690
rect 4050 1680 4100 1690
rect 4150 1680 4250 1690
rect 4450 1680 4500 1690
rect 4600 1680 5900 1690
rect 6400 1680 6450 1690
rect 7300 1680 7350 1690
rect 7850 1680 7900 1690
rect 8450 1680 8550 1690
rect 9100 1680 9150 1690
rect 1900 1670 1950 1680
rect 3200 1670 3250 1680
rect 4050 1670 4100 1680
rect 4150 1670 4250 1680
rect 4450 1670 4500 1680
rect 4600 1670 5900 1680
rect 6400 1670 6450 1680
rect 7300 1670 7350 1680
rect 7850 1670 7900 1680
rect 8450 1670 8550 1680
rect 9100 1670 9150 1680
rect 1900 1660 1950 1670
rect 3200 1660 3250 1670
rect 4050 1660 4100 1670
rect 4150 1660 4250 1670
rect 4450 1660 4500 1670
rect 4600 1660 5900 1670
rect 6400 1660 6450 1670
rect 7300 1660 7350 1670
rect 7850 1660 7900 1670
rect 8450 1660 8550 1670
rect 9100 1660 9150 1670
rect 1900 1650 1950 1660
rect 3200 1650 3250 1660
rect 4050 1650 4100 1660
rect 4150 1650 4250 1660
rect 4450 1650 4500 1660
rect 4600 1650 5900 1660
rect 6400 1650 6450 1660
rect 7300 1650 7350 1660
rect 7850 1650 7900 1660
rect 8450 1650 8550 1660
rect 9100 1650 9150 1660
rect 1950 1640 2000 1650
rect 3150 1640 3200 1650
rect 4150 1640 4300 1650
rect 4950 1640 5450 1650
rect 5500 1640 5900 1650
rect 6800 1640 6850 1650
rect 7850 1640 7900 1650
rect 8400 1640 8500 1650
rect 9150 1640 9200 1650
rect 1950 1630 2000 1640
rect 3150 1630 3200 1640
rect 4150 1630 4300 1640
rect 4950 1630 5450 1640
rect 5500 1630 5900 1640
rect 6800 1630 6850 1640
rect 7850 1630 7900 1640
rect 8400 1630 8500 1640
rect 9150 1630 9200 1640
rect 1950 1620 2000 1630
rect 3150 1620 3200 1630
rect 4150 1620 4300 1630
rect 4950 1620 5450 1630
rect 5500 1620 5900 1630
rect 6800 1620 6850 1630
rect 7850 1620 7900 1630
rect 8400 1620 8500 1630
rect 9150 1620 9200 1630
rect 1950 1610 2000 1620
rect 3150 1610 3200 1620
rect 4150 1610 4300 1620
rect 4950 1610 5450 1620
rect 5500 1610 5900 1620
rect 6800 1610 6850 1620
rect 7850 1610 7900 1620
rect 8400 1610 8500 1620
rect 9150 1610 9200 1620
rect 1950 1600 2000 1610
rect 3150 1600 3200 1610
rect 4150 1600 4300 1610
rect 4950 1600 5450 1610
rect 5500 1600 5900 1610
rect 6800 1600 6850 1610
rect 7850 1600 7900 1610
rect 8400 1600 8500 1610
rect 9150 1600 9200 1610
rect 1950 1590 2000 1600
rect 3100 1590 3150 1600
rect 4150 1590 4250 1600
rect 4300 1590 4350 1600
rect 5100 1590 5650 1600
rect 5700 1590 5800 1600
rect 5850 1590 5900 1600
rect 6800 1590 6850 1600
rect 7850 1590 7900 1600
rect 8300 1590 8350 1600
rect 8400 1590 8450 1600
rect 9800 1590 9850 1600
rect 1950 1580 2000 1590
rect 3100 1580 3150 1590
rect 4150 1580 4250 1590
rect 4300 1580 4350 1590
rect 5100 1580 5650 1590
rect 5700 1580 5800 1590
rect 5850 1580 5900 1590
rect 6800 1580 6850 1590
rect 7850 1580 7900 1590
rect 8300 1580 8350 1590
rect 8400 1580 8450 1590
rect 9800 1580 9850 1590
rect 1950 1570 2000 1580
rect 3100 1570 3150 1580
rect 4150 1570 4250 1580
rect 4300 1570 4350 1580
rect 5100 1570 5650 1580
rect 5700 1570 5800 1580
rect 5850 1570 5900 1580
rect 6800 1570 6850 1580
rect 7850 1570 7900 1580
rect 8300 1570 8350 1580
rect 8400 1570 8450 1580
rect 9800 1570 9850 1580
rect 1950 1560 2000 1570
rect 3100 1560 3150 1570
rect 4150 1560 4250 1570
rect 4300 1560 4350 1570
rect 5100 1560 5650 1570
rect 5700 1560 5800 1570
rect 5850 1560 5900 1570
rect 6800 1560 6850 1570
rect 7850 1560 7900 1570
rect 8300 1560 8350 1570
rect 8400 1560 8450 1570
rect 9800 1560 9850 1570
rect 1950 1550 2000 1560
rect 3100 1550 3150 1560
rect 4150 1550 4250 1560
rect 4300 1550 4350 1560
rect 5100 1550 5650 1560
rect 5700 1550 5800 1560
rect 5850 1550 5900 1560
rect 6800 1550 6850 1560
rect 7850 1550 7900 1560
rect 8300 1550 8350 1560
rect 8400 1550 8450 1560
rect 9800 1550 9850 1560
rect 2000 1540 2050 1550
rect 3050 1540 3100 1550
rect 4150 1540 4250 1550
rect 5250 1540 5350 1550
rect 5400 1540 5800 1550
rect 6800 1540 6850 1550
rect 7850 1540 7900 1550
rect 8400 1540 8450 1550
rect 9700 1540 9750 1550
rect 9800 1540 9850 1550
rect 9950 1540 9990 1550
rect 2000 1530 2050 1540
rect 3050 1530 3100 1540
rect 4150 1530 4250 1540
rect 5250 1530 5350 1540
rect 5400 1530 5800 1540
rect 6800 1530 6850 1540
rect 7850 1530 7900 1540
rect 8400 1530 8450 1540
rect 9700 1530 9750 1540
rect 9800 1530 9850 1540
rect 9950 1530 9990 1540
rect 2000 1520 2050 1530
rect 3050 1520 3100 1530
rect 4150 1520 4250 1530
rect 5250 1520 5350 1530
rect 5400 1520 5800 1530
rect 6800 1520 6850 1530
rect 7850 1520 7900 1530
rect 8400 1520 8450 1530
rect 9700 1520 9750 1530
rect 9800 1520 9850 1530
rect 9950 1520 9990 1530
rect 2000 1510 2050 1520
rect 3050 1510 3100 1520
rect 4150 1510 4250 1520
rect 5250 1510 5350 1520
rect 5400 1510 5800 1520
rect 6800 1510 6850 1520
rect 7850 1510 7900 1520
rect 8400 1510 8450 1520
rect 9700 1510 9750 1520
rect 9800 1510 9850 1520
rect 9950 1510 9990 1520
rect 2000 1500 2050 1510
rect 3050 1500 3100 1510
rect 4150 1500 4250 1510
rect 5250 1500 5350 1510
rect 5400 1500 5800 1510
rect 6800 1500 6850 1510
rect 7850 1500 7900 1510
rect 8400 1500 8450 1510
rect 9700 1500 9750 1510
rect 9800 1500 9850 1510
rect 9950 1500 9990 1510
rect 2050 1490 2100 1500
rect 2950 1490 3050 1500
rect 4350 1490 4400 1500
rect 5400 1490 5800 1500
rect 6800 1490 6850 1500
rect 7350 1490 7400 1500
rect 7850 1490 7900 1500
rect 8400 1490 8450 1500
rect 9700 1490 9750 1500
rect 2050 1480 2100 1490
rect 2950 1480 3050 1490
rect 4350 1480 4400 1490
rect 5400 1480 5800 1490
rect 6800 1480 6850 1490
rect 7350 1480 7400 1490
rect 7850 1480 7900 1490
rect 8400 1480 8450 1490
rect 9700 1480 9750 1490
rect 2050 1470 2100 1480
rect 2950 1470 3050 1480
rect 4350 1470 4400 1480
rect 5400 1470 5800 1480
rect 6800 1470 6850 1480
rect 7350 1470 7400 1480
rect 7850 1470 7900 1480
rect 8400 1470 8450 1480
rect 9700 1470 9750 1480
rect 2050 1460 2100 1470
rect 2950 1460 3050 1470
rect 4350 1460 4400 1470
rect 5400 1460 5800 1470
rect 6800 1460 6850 1470
rect 7350 1460 7400 1470
rect 7850 1460 7900 1470
rect 8400 1460 8450 1470
rect 9700 1460 9750 1470
rect 2050 1450 2100 1460
rect 2950 1450 3050 1460
rect 4350 1450 4400 1460
rect 5400 1450 5800 1460
rect 6800 1450 6850 1460
rect 7350 1450 7400 1460
rect 7850 1450 7900 1460
rect 8400 1450 8450 1460
rect 9700 1450 9750 1460
rect 900 1440 950 1450
rect 2100 1440 2150 1450
rect 2900 1440 2950 1450
rect 4150 1440 4200 1450
rect 5400 1440 5850 1450
rect 6800 1440 6850 1450
rect 7350 1440 7400 1450
rect 7900 1440 7950 1450
rect 8250 1440 8300 1450
rect 8400 1440 8450 1450
rect 900 1430 950 1440
rect 2100 1430 2150 1440
rect 2900 1430 2950 1440
rect 4150 1430 4200 1440
rect 5400 1430 5850 1440
rect 6800 1430 6850 1440
rect 7350 1430 7400 1440
rect 7900 1430 7950 1440
rect 8250 1430 8300 1440
rect 8400 1430 8450 1440
rect 900 1420 950 1430
rect 2100 1420 2150 1430
rect 2900 1420 2950 1430
rect 4150 1420 4200 1430
rect 5400 1420 5850 1430
rect 6800 1420 6850 1430
rect 7350 1420 7400 1430
rect 7900 1420 7950 1430
rect 8250 1420 8300 1430
rect 8400 1420 8450 1430
rect 900 1410 950 1420
rect 2100 1410 2150 1420
rect 2900 1410 2950 1420
rect 4150 1410 4200 1420
rect 5400 1410 5850 1420
rect 6800 1410 6850 1420
rect 7350 1410 7400 1420
rect 7900 1410 7950 1420
rect 8250 1410 8300 1420
rect 8400 1410 8450 1420
rect 900 1400 950 1410
rect 2100 1400 2150 1410
rect 2900 1400 2950 1410
rect 4150 1400 4200 1410
rect 5400 1400 5850 1410
rect 6800 1400 6850 1410
rect 7350 1400 7400 1410
rect 7900 1400 7950 1410
rect 8250 1400 8300 1410
rect 8400 1400 8450 1410
rect 2150 1390 2200 1400
rect 2800 1390 2850 1400
rect 4200 1390 4250 1400
rect 5450 1390 5850 1400
rect 6800 1390 6850 1400
rect 7350 1390 7400 1400
rect 7900 1390 7950 1400
rect 8200 1390 8250 1400
rect 8400 1390 8450 1400
rect 9650 1390 9700 1400
rect 2150 1380 2200 1390
rect 2800 1380 2850 1390
rect 4200 1380 4250 1390
rect 5450 1380 5850 1390
rect 6800 1380 6850 1390
rect 7350 1380 7400 1390
rect 7900 1380 7950 1390
rect 8200 1380 8250 1390
rect 8400 1380 8450 1390
rect 9650 1380 9700 1390
rect 2150 1370 2200 1380
rect 2800 1370 2850 1380
rect 4200 1370 4250 1380
rect 5450 1370 5850 1380
rect 6800 1370 6850 1380
rect 7350 1370 7400 1380
rect 7900 1370 7950 1380
rect 8200 1370 8250 1380
rect 8400 1370 8450 1380
rect 9650 1370 9700 1380
rect 2150 1360 2200 1370
rect 2800 1360 2850 1370
rect 4200 1360 4250 1370
rect 5450 1360 5850 1370
rect 6800 1360 6850 1370
rect 7350 1360 7400 1370
rect 7900 1360 7950 1370
rect 8200 1360 8250 1370
rect 8400 1360 8450 1370
rect 9650 1360 9700 1370
rect 2150 1350 2200 1360
rect 2800 1350 2850 1360
rect 4200 1350 4250 1360
rect 5450 1350 5850 1360
rect 6800 1350 6850 1360
rect 7350 1350 7400 1360
rect 7900 1350 7950 1360
rect 8200 1350 8250 1360
rect 8400 1350 8450 1360
rect 9650 1350 9700 1360
rect 2200 1340 2350 1350
rect 2750 1340 2800 1350
rect 3500 1340 3550 1350
rect 3650 1340 3700 1350
rect 4200 1340 4250 1350
rect 4400 1340 4450 1350
rect 5700 1340 5850 1350
rect 6800 1340 6850 1350
rect 7350 1340 7400 1350
rect 7900 1340 7950 1350
rect 8150 1340 8250 1350
rect 8350 1340 8450 1350
rect 9150 1340 9250 1350
rect 9650 1340 9700 1350
rect 2200 1330 2350 1340
rect 2750 1330 2800 1340
rect 3500 1330 3550 1340
rect 3650 1330 3700 1340
rect 4200 1330 4250 1340
rect 4400 1330 4450 1340
rect 5700 1330 5850 1340
rect 6800 1330 6850 1340
rect 7350 1330 7400 1340
rect 7900 1330 7950 1340
rect 8150 1330 8250 1340
rect 8350 1330 8450 1340
rect 9150 1330 9250 1340
rect 9650 1330 9700 1340
rect 2200 1320 2350 1330
rect 2750 1320 2800 1330
rect 3500 1320 3550 1330
rect 3650 1320 3700 1330
rect 4200 1320 4250 1330
rect 4400 1320 4450 1330
rect 5700 1320 5850 1330
rect 6800 1320 6850 1330
rect 7350 1320 7400 1330
rect 7900 1320 7950 1330
rect 8150 1320 8250 1330
rect 8350 1320 8450 1330
rect 9150 1320 9250 1330
rect 9650 1320 9700 1330
rect 2200 1310 2350 1320
rect 2750 1310 2800 1320
rect 3500 1310 3550 1320
rect 3650 1310 3700 1320
rect 4200 1310 4250 1320
rect 4400 1310 4450 1320
rect 5700 1310 5850 1320
rect 6800 1310 6850 1320
rect 7350 1310 7400 1320
rect 7900 1310 7950 1320
rect 8150 1310 8250 1320
rect 8350 1310 8450 1320
rect 9150 1310 9250 1320
rect 9650 1310 9700 1320
rect 2200 1300 2350 1310
rect 2750 1300 2800 1310
rect 3500 1300 3550 1310
rect 3650 1300 3700 1310
rect 4200 1300 4250 1310
rect 4400 1300 4450 1310
rect 5700 1300 5850 1310
rect 6800 1300 6850 1310
rect 7350 1300 7400 1310
rect 7900 1300 7950 1310
rect 8150 1300 8250 1310
rect 8350 1300 8450 1310
rect 9150 1300 9250 1310
rect 9650 1300 9700 1310
rect 2250 1290 2700 1300
rect 3700 1290 3750 1300
rect 5250 1290 5450 1300
rect 5750 1290 5850 1300
rect 6800 1290 6850 1300
rect 7350 1290 7400 1300
rect 7900 1290 7950 1300
rect 8150 1290 8450 1300
rect 9050 1290 9150 1300
rect 9250 1290 9300 1300
rect 9650 1290 9700 1300
rect 9750 1290 9850 1300
rect 9950 1290 9990 1300
rect 2250 1280 2700 1290
rect 3700 1280 3750 1290
rect 5250 1280 5450 1290
rect 5750 1280 5850 1290
rect 6800 1280 6850 1290
rect 7350 1280 7400 1290
rect 7900 1280 7950 1290
rect 8150 1280 8450 1290
rect 9050 1280 9150 1290
rect 9250 1280 9300 1290
rect 9650 1280 9700 1290
rect 9750 1280 9850 1290
rect 9950 1280 9990 1290
rect 2250 1270 2700 1280
rect 3700 1270 3750 1280
rect 5250 1270 5450 1280
rect 5750 1270 5850 1280
rect 6800 1270 6850 1280
rect 7350 1270 7400 1280
rect 7900 1270 7950 1280
rect 8150 1270 8450 1280
rect 9050 1270 9150 1280
rect 9250 1270 9300 1280
rect 9650 1270 9700 1280
rect 9750 1270 9850 1280
rect 9950 1270 9990 1280
rect 2250 1260 2700 1270
rect 3700 1260 3750 1270
rect 5250 1260 5450 1270
rect 5750 1260 5850 1270
rect 6800 1260 6850 1270
rect 7350 1260 7400 1270
rect 7900 1260 7950 1270
rect 8150 1260 8450 1270
rect 9050 1260 9150 1270
rect 9250 1260 9300 1270
rect 9650 1260 9700 1270
rect 9750 1260 9850 1270
rect 9950 1260 9990 1270
rect 2250 1250 2700 1260
rect 3700 1250 3750 1260
rect 5250 1250 5450 1260
rect 5750 1250 5850 1260
rect 6800 1250 6850 1260
rect 7350 1250 7400 1260
rect 7900 1250 7950 1260
rect 8150 1250 8450 1260
rect 9050 1250 9150 1260
rect 9250 1250 9300 1260
rect 9650 1250 9700 1260
rect 9750 1250 9850 1260
rect 9950 1250 9990 1260
rect 3500 1240 3650 1250
rect 5000 1240 5250 1250
rect 5350 1240 5600 1250
rect 5750 1240 5850 1250
rect 6800 1240 6850 1250
rect 7350 1240 7400 1250
rect 7900 1240 7950 1250
rect 8150 1240 8450 1250
rect 8850 1240 9150 1250
rect 9250 1240 9300 1250
rect 9600 1240 9650 1250
rect 9950 1240 9990 1250
rect 3500 1230 3650 1240
rect 5000 1230 5250 1240
rect 5350 1230 5600 1240
rect 5750 1230 5850 1240
rect 6800 1230 6850 1240
rect 7350 1230 7400 1240
rect 7900 1230 7950 1240
rect 8150 1230 8450 1240
rect 8850 1230 9150 1240
rect 9250 1230 9300 1240
rect 9600 1230 9650 1240
rect 9950 1230 9990 1240
rect 3500 1220 3650 1230
rect 5000 1220 5250 1230
rect 5350 1220 5600 1230
rect 5750 1220 5850 1230
rect 6800 1220 6850 1230
rect 7350 1220 7400 1230
rect 7900 1220 7950 1230
rect 8150 1220 8450 1230
rect 8850 1220 9150 1230
rect 9250 1220 9300 1230
rect 9600 1220 9650 1230
rect 9950 1220 9990 1230
rect 3500 1210 3650 1220
rect 5000 1210 5250 1220
rect 5350 1210 5600 1220
rect 5750 1210 5850 1220
rect 6800 1210 6850 1220
rect 7350 1210 7400 1220
rect 7900 1210 7950 1220
rect 8150 1210 8450 1220
rect 8850 1210 9150 1220
rect 9250 1210 9300 1220
rect 9600 1210 9650 1220
rect 9950 1210 9990 1220
rect 3500 1200 3650 1210
rect 5000 1200 5250 1210
rect 5350 1200 5600 1210
rect 5750 1200 5850 1210
rect 6800 1200 6850 1210
rect 7350 1200 7400 1210
rect 7900 1200 7950 1210
rect 8150 1200 8450 1210
rect 8850 1200 9150 1210
rect 9250 1200 9300 1210
rect 9600 1200 9650 1210
rect 9950 1200 9990 1210
rect 800 1190 850 1200
rect 3600 1190 3700 1200
rect 3850 1190 3900 1200
rect 4700 1190 4900 1200
rect 5000 1190 5050 1200
rect 5400 1190 5600 1200
rect 6650 1190 6700 1200
rect 6800 1190 6850 1200
rect 7350 1190 7400 1200
rect 8150 1190 8450 1200
rect 8700 1190 9100 1200
rect 9250 1190 9300 1200
rect 9600 1190 9650 1200
rect 9700 1190 9750 1200
rect 800 1180 850 1190
rect 3600 1180 3700 1190
rect 3850 1180 3900 1190
rect 4700 1180 4900 1190
rect 5000 1180 5050 1190
rect 5400 1180 5600 1190
rect 6650 1180 6700 1190
rect 6800 1180 6850 1190
rect 7350 1180 7400 1190
rect 8150 1180 8450 1190
rect 8700 1180 9100 1190
rect 9250 1180 9300 1190
rect 9600 1180 9650 1190
rect 9700 1180 9750 1190
rect 800 1170 850 1180
rect 3600 1170 3700 1180
rect 3850 1170 3900 1180
rect 4700 1170 4900 1180
rect 5000 1170 5050 1180
rect 5400 1170 5600 1180
rect 6650 1170 6700 1180
rect 6800 1170 6850 1180
rect 7350 1170 7400 1180
rect 8150 1170 8450 1180
rect 8700 1170 9100 1180
rect 9250 1170 9300 1180
rect 9600 1170 9650 1180
rect 9700 1170 9750 1180
rect 800 1160 850 1170
rect 3600 1160 3700 1170
rect 3850 1160 3900 1170
rect 4700 1160 4900 1170
rect 5000 1160 5050 1170
rect 5400 1160 5600 1170
rect 6650 1160 6700 1170
rect 6800 1160 6850 1170
rect 7350 1160 7400 1170
rect 8150 1160 8450 1170
rect 8700 1160 9100 1170
rect 9250 1160 9300 1170
rect 9600 1160 9650 1170
rect 9700 1160 9750 1170
rect 800 1150 850 1160
rect 3600 1150 3700 1160
rect 3850 1150 3900 1160
rect 4700 1150 4900 1160
rect 5000 1150 5050 1160
rect 5400 1150 5600 1160
rect 6650 1150 6700 1160
rect 6800 1150 6850 1160
rect 7350 1150 7400 1160
rect 8150 1150 8450 1160
rect 8700 1150 9100 1160
rect 9250 1150 9300 1160
rect 9600 1150 9650 1160
rect 9700 1150 9750 1160
rect 750 1140 850 1150
rect 2100 1140 2250 1150
rect 3650 1140 3750 1150
rect 4200 1140 4250 1150
rect 4450 1140 4500 1150
rect 6800 1140 6850 1150
rect 7350 1140 7400 1150
rect 7950 1140 8000 1150
rect 8150 1140 8450 1150
rect 8650 1140 9100 1150
rect 9150 1140 9300 1150
rect 9550 1140 9600 1150
rect 9700 1140 9750 1150
rect 9800 1140 9850 1150
rect 750 1130 850 1140
rect 2100 1130 2250 1140
rect 3650 1130 3750 1140
rect 4200 1130 4250 1140
rect 4450 1130 4500 1140
rect 6800 1130 6850 1140
rect 7350 1130 7400 1140
rect 7950 1130 8000 1140
rect 8150 1130 8450 1140
rect 8650 1130 9100 1140
rect 9150 1130 9300 1140
rect 9550 1130 9600 1140
rect 9700 1130 9750 1140
rect 9800 1130 9850 1140
rect 750 1120 850 1130
rect 2100 1120 2250 1130
rect 3650 1120 3750 1130
rect 4200 1120 4250 1130
rect 4450 1120 4500 1130
rect 6800 1120 6850 1130
rect 7350 1120 7400 1130
rect 7950 1120 8000 1130
rect 8150 1120 8450 1130
rect 8650 1120 9100 1130
rect 9150 1120 9300 1130
rect 9550 1120 9600 1130
rect 9700 1120 9750 1130
rect 9800 1120 9850 1130
rect 750 1110 850 1120
rect 2100 1110 2250 1120
rect 3650 1110 3750 1120
rect 4200 1110 4250 1120
rect 4450 1110 4500 1120
rect 6800 1110 6850 1120
rect 7350 1110 7400 1120
rect 7950 1110 8000 1120
rect 8150 1110 8450 1120
rect 8650 1110 9100 1120
rect 9150 1110 9300 1120
rect 9550 1110 9600 1120
rect 9700 1110 9750 1120
rect 9800 1110 9850 1120
rect 750 1100 850 1110
rect 2100 1100 2250 1110
rect 3650 1100 3750 1110
rect 4200 1100 4250 1110
rect 4450 1100 4500 1110
rect 6800 1100 6850 1110
rect 7350 1100 7400 1110
rect 7950 1100 8000 1110
rect 8150 1100 8450 1110
rect 8650 1100 9100 1110
rect 9150 1100 9300 1110
rect 9550 1100 9600 1110
rect 9700 1100 9750 1110
rect 9800 1100 9850 1110
rect 750 1090 850 1100
rect 1500 1090 1600 1100
rect 2050 1090 2300 1100
rect 3650 1090 3750 1100
rect 4000 1090 4050 1100
rect 4200 1090 4250 1100
rect 6500 1090 6550 1100
rect 6800 1090 6850 1100
rect 7350 1090 7400 1100
rect 7950 1090 8000 1100
rect 8150 1090 8500 1100
rect 8550 1090 9000 1100
rect 9050 1090 9100 1100
rect 9800 1090 9850 1100
rect 9950 1090 9990 1100
rect 750 1080 850 1090
rect 1500 1080 1600 1090
rect 2050 1080 2300 1090
rect 3650 1080 3750 1090
rect 4000 1080 4050 1090
rect 4200 1080 4250 1090
rect 6500 1080 6550 1090
rect 6800 1080 6850 1090
rect 7350 1080 7400 1090
rect 7950 1080 8000 1090
rect 8150 1080 8500 1090
rect 8550 1080 9000 1090
rect 9050 1080 9100 1090
rect 9800 1080 9850 1090
rect 9950 1080 9990 1090
rect 750 1070 850 1080
rect 1500 1070 1600 1080
rect 2050 1070 2300 1080
rect 3650 1070 3750 1080
rect 4000 1070 4050 1080
rect 4200 1070 4250 1080
rect 6500 1070 6550 1080
rect 6800 1070 6850 1080
rect 7350 1070 7400 1080
rect 7950 1070 8000 1080
rect 8150 1070 8500 1080
rect 8550 1070 9000 1080
rect 9050 1070 9100 1080
rect 9800 1070 9850 1080
rect 9950 1070 9990 1080
rect 750 1060 850 1070
rect 1500 1060 1600 1070
rect 2050 1060 2300 1070
rect 3650 1060 3750 1070
rect 4000 1060 4050 1070
rect 4200 1060 4250 1070
rect 6500 1060 6550 1070
rect 6800 1060 6850 1070
rect 7350 1060 7400 1070
rect 7950 1060 8000 1070
rect 8150 1060 8500 1070
rect 8550 1060 9000 1070
rect 9050 1060 9100 1070
rect 9800 1060 9850 1070
rect 9950 1060 9990 1070
rect 750 1050 850 1060
rect 1500 1050 1600 1060
rect 2050 1050 2300 1060
rect 3650 1050 3750 1060
rect 4000 1050 4050 1060
rect 4200 1050 4250 1060
rect 6500 1050 6550 1060
rect 6800 1050 6850 1060
rect 7350 1050 7400 1060
rect 7950 1050 8000 1060
rect 8150 1050 8500 1060
rect 8550 1050 9000 1060
rect 9050 1050 9100 1060
rect 9800 1050 9850 1060
rect 9950 1050 9990 1060
rect 750 1040 850 1050
rect 1450 1040 1550 1050
rect 2050 1040 2100 1050
rect 2200 1040 2800 1050
rect 3700 1040 3850 1050
rect 4650 1040 4700 1050
rect 6450 1040 6500 1050
rect 6800 1040 6850 1050
rect 7350 1040 7400 1050
rect 7950 1040 8000 1050
rect 8100 1040 8150 1050
rect 8250 1040 8400 1050
rect 8500 1040 8900 1050
rect 9100 1040 9150 1050
rect 9750 1040 9850 1050
rect 750 1030 850 1040
rect 1450 1030 1550 1040
rect 2050 1030 2100 1040
rect 2200 1030 2800 1040
rect 3700 1030 3850 1040
rect 4650 1030 4700 1040
rect 6450 1030 6500 1040
rect 6800 1030 6850 1040
rect 7350 1030 7400 1040
rect 7950 1030 8000 1040
rect 8100 1030 8150 1040
rect 8250 1030 8400 1040
rect 8500 1030 8900 1040
rect 9100 1030 9150 1040
rect 9750 1030 9850 1040
rect 750 1020 850 1030
rect 1450 1020 1550 1030
rect 2050 1020 2100 1030
rect 2200 1020 2800 1030
rect 3700 1020 3850 1030
rect 4650 1020 4700 1030
rect 6450 1020 6500 1030
rect 6800 1020 6850 1030
rect 7350 1020 7400 1030
rect 7950 1020 8000 1030
rect 8100 1020 8150 1030
rect 8250 1020 8400 1030
rect 8500 1020 8900 1030
rect 9100 1020 9150 1030
rect 9750 1020 9850 1030
rect 750 1010 850 1020
rect 1450 1010 1550 1020
rect 2050 1010 2100 1020
rect 2200 1010 2800 1020
rect 3700 1010 3850 1020
rect 4650 1010 4700 1020
rect 6450 1010 6500 1020
rect 6800 1010 6850 1020
rect 7350 1010 7400 1020
rect 7950 1010 8000 1020
rect 8100 1010 8150 1020
rect 8250 1010 8400 1020
rect 8500 1010 8900 1020
rect 9100 1010 9150 1020
rect 9750 1010 9850 1020
rect 750 1000 850 1010
rect 1450 1000 1550 1010
rect 2050 1000 2100 1010
rect 2200 1000 2800 1010
rect 3700 1000 3850 1010
rect 4650 1000 4700 1010
rect 6450 1000 6500 1010
rect 6800 1000 6850 1010
rect 7350 1000 7400 1010
rect 7950 1000 8000 1010
rect 8100 1000 8150 1010
rect 8250 1000 8400 1010
rect 8500 1000 8900 1010
rect 9100 1000 9150 1010
rect 9750 1000 9850 1010
rect 700 990 800 1000
rect 1400 990 1500 1000
rect 2000 990 2050 1000
rect 2300 990 2750 1000
rect 3750 990 3850 1000
rect 4750 990 4800 1000
rect 5450 990 5500 1000
rect 6450 990 6500 1000
rect 6800 990 6850 1000
rect 7350 990 7400 1000
rect 7950 990 8000 1000
rect 8100 990 8150 1000
rect 8250 990 8400 1000
rect 8550 990 8900 1000
rect 9100 990 9150 1000
rect 700 980 800 990
rect 1400 980 1500 990
rect 2000 980 2050 990
rect 2300 980 2750 990
rect 3750 980 3850 990
rect 4750 980 4800 990
rect 5450 980 5500 990
rect 6450 980 6500 990
rect 6800 980 6850 990
rect 7350 980 7400 990
rect 7950 980 8000 990
rect 8100 980 8150 990
rect 8250 980 8400 990
rect 8550 980 8900 990
rect 9100 980 9150 990
rect 700 970 800 980
rect 1400 970 1500 980
rect 2000 970 2050 980
rect 2300 970 2750 980
rect 3750 970 3850 980
rect 4750 970 4800 980
rect 5450 970 5500 980
rect 6450 970 6500 980
rect 6800 970 6850 980
rect 7350 970 7400 980
rect 7950 970 8000 980
rect 8100 970 8150 980
rect 8250 970 8400 980
rect 8550 970 8900 980
rect 9100 970 9150 980
rect 700 960 800 970
rect 1400 960 1500 970
rect 2000 960 2050 970
rect 2300 960 2750 970
rect 3750 960 3850 970
rect 4750 960 4800 970
rect 5450 960 5500 970
rect 6450 960 6500 970
rect 6800 960 6850 970
rect 7350 960 7400 970
rect 7950 960 8000 970
rect 8100 960 8150 970
rect 8250 960 8400 970
rect 8550 960 8900 970
rect 9100 960 9150 970
rect 700 950 800 960
rect 1400 950 1500 960
rect 2000 950 2050 960
rect 2300 950 2750 960
rect 3750 950 3850 960
rect 4750 950 4800 960
rect 5450 950 5500 960
rect 6450 950 6500 960
rect 6800 950 6850 960
rect 7350 950 7400 960
rect 7950 950 8000 960
rect 8100 950 8150 960
rect 8250 950 8400 960
rect 8550 950 8900 960
rect 9100 950 9150 960
rect 700 940 800 950
rect 1350 940 1450 950
rect 2000 940 2050 950
rect 2700 940 2750 950
rect 3800 940 3850 950
rect 5350 940 5800 950
rect 6450 940 6500 950
rect 7350 940 7400 950
rect 7950 940 8000 950
rect 8100 940 8150 950
rect 8250 940 8450 950
rect 8550 940 8850 950
rect 9100 940 9150 950
rect 9450 940 9500 950
rect 700 930 800 940
rect 1350 930 1450 940
rect 2000 930 2050 940
rect 2700 930 2750 940
rect 3800 930 3850 940
rect 5350 930 5800 940
rect 6450 930 6500 940
rect 7350 930 7400 940
rect 7950 930 8000 940
rect 8100 930 8150 940
rect 8250 930 8450 940
rect 8550 930 8850 940
rect 9100 930 9150 940
rect 9450 930 9500 940
rect 700 920 800 930
rect 1350 920 1450 930
rect 2000 920 2050 930
rect 2700 920 2750 930
rect 3800 920 3850 930
rect 5350 920 5800 930
rect 6450 920 6500 930
rect 7350 920 7400 930
rect 7950 920 8000 930
rect 8100 920 8150 930
rect 8250 920 8450 930
rect 8550 920 8850 930
rect 9100 920 9150 930
rect 9450 920 9500 930
rect 700 910 800 920
rect 1350 910 1450 920
rect 2000 910 2050 920
rect 2700 910 2750 920
rect 3800 910 3850 920
rect 5350 910 5800 920
rect 6450 910 6500 920
rect 7350 910 7400 920
rect 7950 910 8000 920
rect 8100 910 8150 920
rect 8250 910 8450 920
rect 8550 910 8850 920
rect 9100 910 9150 920
rect 9450 910 9500 920
rect 700 900 800 910
rect 1350 900 1450 910
rect 2000 900 2050 910
rect 2700 900 2750 910
rect 3800 900 3850 910
rect 5350 900 5800 910
rect 6450 900 6500 910
rect 7350 900 7400 910
rect 7950 900 8000 910
rect 8100 900 8150 910
rect 8250 900 8450 910
rect 8550 900 8850 910
rect 9100 900 9150 910
rect 9450 900 9500 910
rect 650 890 700 900
rect 750 890 800 900
rect 1300 890 1400 900
rect 2000 890 2050 900
rect 2650 890 2700 900
rect 3850 890 3900 900
rect 4850 890 4900 900
rect 5350 890 5500 900
rect 6450 890 6500 900
rect 7350 890 7400 900
rect 7950 890 8000 900
rect 8100 890 8150 900
rect 8250 890 8450 900
rect 8600 890 8800 900
rect 650 880 700 890
rect 750 880 800 890
rect 1300 880 1400 890
rect 2000 880 2050 890
rect 2650 880 2700 890
rect 3850 880 3900 890
rect 4850 880 4900 890
rect 5350 880 5500 890
rect 6450 880 6500 890
rect 7350 880 7400 890
rect 7950 880 8000 890
rect 8100 880 8150 890
rect 8250 880 8450 890
rect 8600 880 8800 890
rect 650 870 700 880
rect 750 870 800 880
rect 1300 870 1400 880
rect 2000 870 2050 880
rect 2650 870 2700 880
rect 3850 870 3900 880
rect 4850 870 4900 880
rect 5350 870 5500 880
rect 6450 870 6500 880
rect 7350 870 7400 880
rect 7950 870 8000 880
rect 8100 870 8150 880
rect 8250 870 8450 880
rect 8600 870 8800 880
rect 650 860 700 870
rect 750 860 800 870
rect 1300 860 1400 870
rect 2000 860 2050 870
rect 2650 860 2700 870
rect 3850 860 3900 870
rect 4850 860 4900 870
rect 5350 860 5500 870
rect 6450 860 6500 870
rect 7350 860 7400 870
rect 7950 860 8000 870
rect 8100 860 8150 870
rect 8250 860 8450 870
rect 8600 860 8800 870
rect 650 850 700 860
rect 750 850 800 860
rect 1300 850 1400 860
rect 2000 850 2050 860
rect 2650 850 2700 860
rect 3850 850 3900 860
rect 4850 850 4900 860
rect 5350 850 5500 860
rect 6450 850 6500 860
rect 7350 850 7400 860
rect 7950 850 8000 860
rect 8100 850 8150 860
rect 8250 850 8450 860
rect 8600 850 8800 860
rect 650 840 700 850
rect 750 840 800 850
rect 1200 840 1350 850
rect 2050 840 2100 850
rect 2600 840 2650 850
rect 3900 840 4000 850
rect 6450 840 6500 850
rect 7350 840 7400 850
rect 8100 840 8150 850
rect 8300 840 8750 850
rect 9150 840 9200 850
rect 9400 840 9450 850
rect 650 830 700 840
rect 750 830 800 840
rect 1200 830 1350 840
rect 2050 830 2100 840
rect 2600 830 2650 840
rect 3900 830 4000 840
rect 6450 830 6500 840
rect 7350 830 7400 840
rect 8100 830 8150 840
rect 8300 830 8750 840
rect 9150 830 9200 840
rect 9400 830 9450 840
rect 650 820 700 830
rect 750 820 800 830
rect 1200 820 1350 830
rect 2050 820 2100 830
rect 2600 820 2650 830
rect 3900 820 4000 830
rect 6450 820 6500 830
rect 7350 820 7400 830
rect 8100 820 8150 830
rect 8300 820 8750 830
rect 9150 820 9200 830
rect 9400 820 9450 830
rect 650 810 700 820
rect 750 810 800 820
rect 1200 810 1350 820
rect 2050 810 2100 820
rect 2600 810 2650 820
rect 3900 810 4000 820
rect 6450 810 6500 820
rect 7350 810 7400 820
rect 8100 810 8150 820
rect 8300 810 8750 820
rect 9150 810 9200 820
rect 9400 810 9450 820
rect 650 800 700 810
rect 750 800 800 810
rect 1200 800 1350 810
rect 2050 800 2100 810
rect 2600 800 2650 810
rect 3900 800 4000 810
rect 6450 800 6500 810
rect 7350 800 7400 810
rect 8100 800 8150 810
rect 8300 800 8750 810
rect 9150 800 9200 810
rect 9400 800 9450 810
rect 700 790 750 800
rect 1150 790 1300 800
rect 2050 790 2100 800
rect 3600 790 3850 800
rect 6500 790 6550 800
rect 7350 790 7400 800
rect 8000 790 8050 800
rect 8100 790 8150 800
rect 8300 790 8750 800
rect 9150 790 9200 800
rect 700 780 750 790
rect 1150 780 1300 790
rect 2050 780 2100 790
rect 3600 780 3850 790
rect 6500 780 6550 790
rect 7350 780 7400 790
rect 8000 780 8050 790
rect 8100 780 8150 790
rect 8300 780 8750 790
rect 9150 780 9200 790
rect 700 770 750 780
rect 1150 770 1300 780
rect 2050 770 2100 780
rect 3600 770 3850 780
rect 6500 770 6550 780
rect 7350 770 7400 780
rect 8000 770 8050 780
rect 8100 770 8150 780
rect 8300 770 8750 780
rect 9150 770 9200 780
rect 700 760 750 770
rect 1150 760 1300 770
rect 2050 760 2100 770
rect 3600 760 3850 770
rect 6500 760 6550 770
rect 7350 760 7400 770
rect 8000 760 8050 770
rect 8100 760 8150 770
rect 8300 760 8750 770
rect 9150 760 9200 770
rect 700 750 750 760
rect 1150 750 1300 760
rect 2050 750 2100 760
rect 3600 750 3850 760
rect 6500 750 6550 760
rect 7350 750 7400 760
rect 8000 750 8050 760
rect 8100 750 8150 760
rect 8300 750 8750 760
rect 9150 750 9200 760
rect 600 740 650 750
rect 700 740 750 750
rect 1100 740 1150 750
rect 1200 740 1250 750
rect 3400 740 3450 750
rect 3900 740 3950 750
rect 4900 740 4950 750
rect 6200 740 6250 750
rect 6500 740 6550 750
rect 6850 740 6900 750
rect 7350 740 7400 750
rect 8000 740 8050 750
rect 8100 740 8150 750
rect 8350 740 8700 750
rect 9350 740 9400 750
rect 600 730 650 740
rect 700 730 750 740
rect 1100 730 1150 740
rect 1200 730 1250 740
rect 3400 730 3450 740
rect 3900 730 3950 740
rect 4900 730 4950 740
rect 6200 730 6250 740
rect 6500 730 6550 740
rect 6850 730 6900 740
rect 7350 730 7400 740
rect 8000 730 8050 740
rect 8100 730 8150 740
rect 8350 730 8700 740
rect 9350 730 9400 740
rect 600 720 650 730
rect 700 720 750 730
rect 1100 720 1150 730
rect 1200 720 1250 730
rect 3400 720 3450 730
rect 3900 720 3950 730
rect 4900 720 4950 730
rect 6200 720 6250 730
rect 6500 720 6550 730
rect 6850 720 6900 730
rect 7350 720 7400 730
rect 8000 720 8050 730
rect 8100 720 8150 730
rect 8350 720 8700 730
rect 9350 720 9400 730
rect 600 710 650 720
rect 700 710 750 720
rect 1100 710 1150 720
rect 1200 710 1250 720
rect 3400 710 3450 720
rect 3900 710 3950 720
rect 4900 710 4950 720
rect 6200 710 6250 720
rect 6500 710 6550 720
rect 6850 710 6900 720
rect 7350 710 7400 720
rect 8000 710 8050 720
rect 8100 710 8150 720
rect 8350 710 8700 720
rect 9350 710 9400 720
rect 600 700 650 710
rect 700 700 750 710
rect 1100 700 1150 710
rect 1200 700 1250 710
rect 3400 700 3450 710
rect 3900 700 3950 710
rect 4900 700 4950 710
rect 6200 700 6250 710
rect 6500 700 6550 710
rect 6850 700 6900 710
rect 7350 700 7400 710
rect 8000 700 8050 710
rect 8100 700 8150 710
rect 8350 700 8700 710
rect 9350 700 9400 710
rect 600 690 700 700
rect 1050 690 1100 700
rect 1150 690 1250 700
rect 2100 690 2150 700
rect 2350 690 2400 700
rect 4100 690 4150 700
rect 4700 690 4750 700
rect 4900 690 4950 700
rect 6050 690 6150 700
rect 6550 690 6600 700
rect 6850 690 6900 700
rect 7300 690 7350 700
rect 8000 690 8050 700
rect 8100 690 8150 700
rect 8400 690 8650 700
rect 9150 690 9200 700
rect 600 680 700 690
rect 1050 680 1100 690
rect 1150 680 1250 690
rect 2100 680 2150 690
rect 2350 680 2400 690
rect 4100 680 4150 690
rect 4700 680 4750 690
rect 4900 680 4950 690
rect 6050 680 6150 690
rect 6550 680 6600 690
rect 6850 680 6900 690
rect 7300 680 7350 690
rect 8000 680 8050 690
rect 8100 680 8150 690
rect 8400 680 8650 690
rect 9150 680 9200 690
rect 600 670 700 680
rect 1050 670 1100 680
rect 1150 670 1250 680
rect 2100 670 2150 680
rect 2350 670 2400 680
rect 4100 670 4150 680
rect 4700 670 4750 680
rect 4900 670 4950 680
rect 6050 670 6150 680
rect 6550 670 6600 680
rect 6850 670 6900 680
rect 7300 670 7350 680
rect 8000 670 8050 680
rect 8100 670 8150 680
rect 8400 670 8650 680
rect 9150 670 9200 680
rect 600 660 700 670
rect 1050 660 1100 670
rect 1150 660 1250 670
rect 2100 660 2150 670
rect 2350 660 2400 670
rect 4100 660 4150 670
rect 4700 660 4750 670
rect 4900 660 4950 670
rect 6050 660 6150 670
rect 6550 660 6600 670
rect 6850 660 6900 670
rect 7300 660 7350 670
rect 8000 660 8050 670
rect 8100 660 8150 670
rect 8400 660 8650 670
rect 9150 660 9200 670
rect 600 650 700 660
rect 1050 650 1100 660
rect 1150 650 1250 660
rect 2100 650 2150 660
rect 2350 650 2400 660
rect 4100 650 4150 660
rect 4700 650 4750 660
rect 4900 650 4950 660
rect 6050 650 6150 660
rect 6550 650 6600 660
rect 6850 650 6900 660
rect 7300 650 7350 660
rect 8000 650 8050 660
rect 8100 650 8150 660
rect 8400 650 8650 660
rect 9150 650 9200 660
rect 450 640 800 650
rect 900 640 1200 650
rect 2100 640 2150 650
rect 2200 640 2300 650
rect 3150 640 3250 650
rect 5950 640 6250 650
rect 6550 640 6600 650
rect 7300 640 7350 650
rect 8050 640 8150 650
rect 8450 640 8550 650
rect 9150 640 9200 650
rect 450 630 800 640
rect 900 630 1200 640
rect 2100 630 2150 640
rect 2200 630 2300 640
rect 3150 630 3250 640
rect 5950 630 6250 640
rect 6550 630 6600 640
rect 7300 630 7350 640
rect 8050 630 8150 640
rect 8450 630 8550 640
rect 9150 630 9200 640
rect 450 620 800 630
rect 900 620 1200 630
rect 2100 620 2150 630
rect 2200 620 2300 630
rect 3150 620 3250 630
rect 5950 620 6250 630
rect 6550 620 6600 630
rect 7300 620 7350 630
rect 8050 620 8150 630
rect 8450 620 8550 630
rect 9150 620 9200 630
rect 450 610 800 620
rect 900 610 1200 620
rect 2100 610 2150 620
rect 2200 610 2300 620
rect 3150 610 3250 620
rect 5950 610 6250 620
rect 6550 610 6600 620
rect 7300 610 7350 620
rect 8050 610 8150 620
rect 8450 610 8550 620
rect 9150 610 9200 620
rect 450 600 800 610
rect 900 600 1200 610
rect 2100 600 2150 610
rect 2200 600 2300 610
rect 3150 600 3250 610
rect 5950 600 6250 610
rect 6550 600 6600 610
rect 7300 600 7350 610
rect 8050 600 8150 610
rect 8450 600 8550 610
rect 9150 600 9200 610
rect 650 590 800 600
rect 850 590 950 600
rect 1050 590 1100 600
rect 1250 590 1450 600
rect 3050 590 3100 600
rect 4500 590 4550 600
rect 4650 590 4700 600
rect 4750 590 4800 600
rect 6000 590 6250 600
rect 6600 590 6650 600
rect 6900 590 6950 600
rect 7300 590 7350 600
rect 9150 590 9200 600
rect 9250 590 9300 600
rect 650 580 800 590
rect 850 580 950 590
rect 1050 580 1100 590
rect 1250 580 1450 590
rect 3050 580 3100 590
rect 4500 580 4550 590
rect 4650 580 4700 590
rect 4750 580 4800 590
rect 6000 580 6250 590
rect 6600 580 6650 590
rect 6900 580 6950 590
rect 7300 580 7350 590
rect 9150 580 9200 590
rect 9250 580 9300 590
rect 650 570 800 580
rect 850 570 950 580
rect 1050 570 1100 580
rect 1250 570 1450 580
rect 3050 570 3100 580
rect 4500 570 4550 580
rect 4650 570 4700 580
rect 4750 570 4800 580
rect 6000 570 6250 580
rect 6600 570 6650 580
rect 6900 570 6950 580
rect 7300 570 7350 580
rect 9150 570 9200 580
rect 9250 570 9300 580
rect 650 560 800 570
rect 850 560 950 570
rect 1050 560 1100 570
rect 1250 560 1450 570
rect 3050 560 3100 570
rect 4500 560 4550 570
rect 4650 560 4700 570
rect 4750 560 4800 570
rect 6000 560 6250 570
rect 6600 560 6650 570
rect 6900 560 6950 570
rect 7300 560 7350 570
rect 9150 560 9200 570
rect 9250 560 9300 570
rect 650 550 800 560
rect 850 550 950 560
rect 1050 550 1100 560
rect 1250 550 1450 560
rect 3050 550 3100 560
rect 4500 550 4550 560
rect 4650 550 4700 560
rect 4750 550 4800 560
rect 6000 550 6250 560
rect 6600 550 6650 560
rect 6900 550 6950 560
rect 7300 550 7350 560
rect 9150 550 9200 560
rect 9250 550 9300 560
rect 300 540 350 550
rect 600 540 650 550
rect 900 540 1050 550
rect 1200 540 1250 550
rect 4300 540 4450 550
rect 4550 540 4650 550
rect 6050 540 6250 550
rect 6650 540 6700 550
rect 6900 540 6950 550
rect 7250 540 7350 550
rect 9150 540 9250 550
rect 300 530 350 540
rect 600 530 650 540
rect 900 530 1050 540
rect 1200 530 1250 540
rect 4300 530 4450 540
rect 4550 530 4650 540
rect 6050 530 6250 540
rect 6650 530 6700 540
rect 6900 530 6950 540
rect 7250 530 7350 540
rect 9150 530 9250 540
rect 300 520 350 530
rect 600 520 650 530
rect 900 520 1050 530
rect 1200 520 1250 530
rect 4300 520 4450 530
rect 4550 520 4650 530
rect 6050 520 6250 530
rect 6650 520 6700 530
rect 6900 520 6950 530
rect 7250 520 7350 530
rect 9150 520 9250 530
rect 300 510 350 520
rect 600 510 650 520
rect 900 510 1050 520
rect 1200 510 1250 520
rect 4300 510 4450 520
rect 4550 510 4650 520
rect 6050 510 6250 520
rect 6650 510 6700 520
rect 6900 510 6950 520
rect 7250 510 7350 520
rect 9150 510 9250 520
rect 300 500 350 510
rect 600 500 650 510
rect 900 500 1050 510
rect 1200 500 1250 510
rect 4300 500 4450 510
rect 4550 500 4650 510
rect 6050 500 6250 510
rect 6650 500 6700 510
rect 6900 500 6950 510
rect 7250 500 7350 510
rect 9150 500 9250 510
rect 300 490 400 500
rect 500 490 550 500
rect 2100 490 2200 500
rect 2750 490 2800 500
rect 4950 490 5000 500
rect 6050 490 6200 500
rect 6650 490 6700 500
rect 7250 490 7300 500
rect 9100 490 9250 500
rect 300 480 400 490
rect 500 480 550 490
rect 2100 480 2200 490
rect 2750 480 2800 490
rect 4950 480 5000 490
rect 6050 480 6200 490
rect 6650 480 6700 490
rect 7250 480 7300 490
rect 9100 480 9250 490
rect 300 470 400 480
rect 500 470 550 480
rect 2100 470 2200 480
rect 2750 470 2800 480
rect 4950 470 5000 480
rect 6050 470 6200 480
rect 6650 470 6700 480
rect 7250 470 7300 480
rect 9100 470 9250 480
rect 300 460 400 470
rect 500 460 550 470
rect 2100 460 2200 470
rect 2750 460 2800 470
rect 4950 460 5000 470
rect 6050 460 6200 470
rect 6650 460 6700 470
rect 7250 460 7300 470
rect 9100 460 9250 470
rect 300 450 400 460
rect 500 450 550 460
rect 2100 450 2200 460
rect 2750 450 2800 460
rect 4950 450 5000 460
rect 6050 450 6200 460
rect 6650 450 6700 460
rect 7250 450 7300 460
rect 9100 450 9250 460
rect 350 440 500 450
rect 1700 440 1800 450
rect 2300 440 2550 450
rect 4200 440 4250 450
rect 4950 440 5000 450
rect 6050 440 6200 450
rect 6700 440 6750 450
rect 7200 440 7300 450
rect 9100 440 9200 450
rect 350 430 500 440
rect 1700 430 1800 440
rect 2300 430 2550 440
rect 4200 430 4250 440
rect 4950 430 5000 440
rect 6050 430 6200 440
rect 6700 430 6750 440
rect 7200 430 7300 440
rect 9100 430 9200 440
rect 350 420 500 430
rect 1700 420 1800 430
rect 2300 420 2550 430
rect 4200 420 4250 430
rect 4950 420 5000 430
rect 6050 420 6200 430
rect 6700 420 6750 430
rect 7200 420 7300 430
rect 9100 420 9200 430
rect 350 410 500 420
rect 1700 410 1800 420
rect 2300 410 2550 420
rect 4200 410 4250 420
rect 4950 410 5000 420
rect 6050 410 6200 420
rect 6700 410 6750 420
rect 7200 410 7300 420
rect 9100 410 9200 420
rect 350 400 500 410
rect 1700 400 1800 410
rect 2300 400 2550 410
rect 4200 400 4250 410
rect 4950 400 5000 410
rect 6050 400 6200 410
rect 6700 400 6750 410
rect 7200 400 7300 410
rect 9100 400 9200 410
rect 350 390 400 400
rect 450 390 500 400
rect 1050 390 1100 400
rect 4200 390 4250 400
rect 4300 390 4350 400
rect 4700 390 4750 400
rect 4950 390 5000 400
rect 6050 390 6200 400
rect 6750 390 6800 400
rect 7200 390 7300 400
rect 9100 390 9200 400
rect 9250 390 9400 400
rect 350 380 400 390
rect 450 380 500 390
rect 1050 380 1100 390
rect 4200 380 4250 390
rect 4300 380 4350 390
rect 4700 380 4750 390
rect 4950 380 5000 390
rect 6050 380 6200 390
rect 6750 380 6800 390
rect 7200 380 7300 390
rect 9100 380 9200 390
rect 9250 380 9400 390
rect 350 370 400 380
rect 450 370 500 380
rect 1050 370 1100 380
rect 4200 370 4250 380
rect 4300 370 4350 380
rect 4700 370 4750 380
rect 4950 370 5000 380
rect 6050 370 6200 380
rect 6750 370 6800 380
rect 7200 370 7300 380
rect 9100 370 9200 380
rect 9250 370 9400 380
rect 350 360 400 370
rect 450 360 500 370
rect 1050 360 1100 370
rect 4200 360 4250 370
rect 4300 360 4350 370
rect 4700 360 4750 370
rect 4950 360 5000 370
rect 6050 360 6200 370
rect 6750 360 6800 370
rect 7200 360 7300 370
rect 9100 360 9200 370
rect 9250 360 9400 370
rect 350 350 400 360
rect 450 350 500 360
rect 1050 350 1100 360
rect 4200 350 4250 360
rect 4300 350 4350 360
rect 4700 350 4750 360
rect 4950 350 5000 360
rect 6050 350 6200 360
rect 6750 350 6800 360
rect 7200 350 7300 360
rect 9100 350 9200 360
rect 9250 350 9400 360
rect 0 340 50 350
rect 350 340 400 350
rect 450 340 700 350
rect 4150 340 4300 350
rect 4350 340 4450 350
rect 4700 340 4750 350
rect 4950 340 5000 350
rect 6150 340 6200 350
rect 6750 340 6850 350
rect 7100 340 7250 350
rect 9050 340 9150 350
rect 0 330 50 340
rect 350 330 400 340
rect 450 330 700 340
rect 4150 330 4300 340
rect 4350 330 4450 340
rect 4700 330 4750 340
rect 4950 330 5000 340
rect 6150 330 6200 340
rect 6750 330 6850 340
rect 7100 330 7250 340
rect 9050 330 9150 340
rect 0 320 50 330
rect 350 320 400 330
rect 450 320 700 330
rect 4150 320 4300 330
rect 4350 320 4450 330
rect 4700 320 4750 330
rect 4950 320 5000 330
rect 6150 320 6200 330
rect 6750 320 6850 330
rect 7100 320 7250 330
rect 9050 320 9150 330
rect 0 310 50 320
rect 350 310 400 320
rect 450 310 700 320
rect 4150 310 4300 320
rect 4350 310 4450 320
rect 4700 310 4750 320
rect 4950 310 5000 320
rect 6150 310 6200 320
rect 6750 310 6850 320
rect 7100 310 7250 320
rect 9050 310 9150 320
rect 0 300 50 310
rect 350 300 400 310
rect 450 300 700 310
rect 4150 300 4300 310
rect 4350 300 4450 310
rect 4700 300 4750 310
rect 4950 300 5000 310
rect 6150 300 6200 310
rect 6750 300 6850 310
rect 7100 300 7250 310
rect 9050 300 9150 310
rect 0 290 50 300
rect 350 290 500 300
rect 600 290 700 300
rect 800 290 900 300
rect 1000 290 1050 300
rect 4100 290 4250 300
rect 4500 290 4550 300
rect 4650 290 4700 300
rect 6850 290 7250 300
rect 9050 290 9100 300
rect 9200 290 9250 300
rect 9400 290 9450 300
rect 0 280 50 290
rect 350 280 500 290
rect 600 280 700 290
rect 800 280 900 290
rect 1000 280 1050 290
rect 4100 280 4250 290
rect 4500 280 4550 290
rect 4650 280 4700 290
rect 6850 280 7250 290
rect 9050 280 9100 290
rect 9200 280 9250 290
rect 9400 280 9450 290
rect 0 270 50 280
rect 350 270 500 280
rect 600 270 700 280
rect 800 270 900 280
rect 1000 270 1050 280
rect 4100 270 4250 280
rect 4500 270 4550 280
rect 4650 270 4700 280
rect 6850 270 7250 280
rect 9050 270 9100 280
rect 9200 270 9250 280
rect 9400 270 9450 280
rect 0 260 50 270
rect 350 260 500 270
rect 600 260 700 270
rect 800 260 900 270
rect 1000 260 1050 270
rect 4100 260 4250 270
rect 4500 260 4550 270
rect 4650 260 4700 270
rect 6850 260 7250 270
rect 9050 260 9100 270
rect 9200 260 9250 270
rect 9400 260 9450 270
rect 0 250 50 260
rect 350 250 500 260
rect 600 250 700 260
rect 800 250 900 260
rect 1000 250 1050 260
rect 4100 250 4250 260
rect 4500 250 4550 260
rect 4650 250 4700 260
rect 6850 250 7250 260
rect 9050 250 9100 260
rect 9200 250 9250 260
rect 9400 250 9450 260
rect 0 240 150 250
rect 200 240 250 250
rect 350 240 450 250
rect 600 240 700 250
rect 850 240 1000 250
rect 4150 240 4250 250
rect 4300 240 4400 250
rect 4500 240 4650 250
rect 4850 240 4900 250
rect 6950 240 7250 250
rect 8850 240 8950 250
rect 9000 240 9100 250
rect 9250 240 9350 250
rect 0 230 150 240
rect 200 230 250 240
rect 350 230 450 240
rect 600 230 700 240
rect 850 230 1000 240
rect 4150 230 4250 240
rect 4300 230 4400 240
rect 4500 230 4650 240
rect 4850 230 4900 240
rect 6950 230 7250 240
rect 8850 230 8950 240
rect 9000 230 9100 240
rect 9250 230 9350 240
rect 0 220 150 230
rect 200 220 250 230
rect 350 220 450 230
rect 600 220 700 230
rect 850 220 1000 230
rect 4150 220 4250 230
rect 4300 220 4400 230
rect 4500 220 4650 230
rect 4850 220 4900 230
rect 6950 220 7250 230
rect 8850 220 8950 230
rect 9000 220 9100 230
rect 9250 220 9350 230
rect 0 210 150 220
rect 200 210 250 220
rect 350 210 450 220
rect 600 210 700 220
rect 850 210 1000 220
rect 4150 210 4250 220
rect 4300 210 4400 220
rect 4500 210 4650 220
rect 4850 210 4900 220
rect 6950 210 7250 220
rect 8850 210 8950 220
rect 9000 210 9100 220
rect 9250 210 9350 220
rect 0 200 150 210
rect 200 200 250 210
rect 350 200 450 210
rect 600 200 700 210
rect 850 200 1000 210
rect 4150 200 4250 210
rect 4300 200 4400 210
rect 4500 200 4650 210
rect 4850 200 4900 210
rect 6950 200 7250 210
rect 8850 200 8950 210
rect 9000 200 9100 210
rect 9250 200 9350 210
rect 0 190 100 200
rect 200 190 350 200
rect 450 190 1000 200
rect 4150 190 4600 200
rect 4800 190 4900 200
rect 6150 190 6250 200
rect 7050 190 7250 200
rect 8850 190 8900 200
rect 9000 190 9100 200
rect 9150 190 9200 200
rect 9300 190 9350 200
rect 9750 190 9800 200
rect 9850 190 9990 200
rect 0 180 100 190
rect 200 180 350 190
rect 450 180 1000 190
rect 4150 180 4600 190
rect 4800 180 4900 190
rect 6150 180 6250 190
rect 7050 180 7250 190
rect 8850 180 8900 190
rect 9000 180 9100 190
rect 9150 180 9200 190
rect 9300 180 9350 190
rect 9750 180 9800 190
rect 9850 180 9990 190
rect 0 170 100 180
rect 200 170 350 180
rect 450 170 1000 180
rect 4150 170 4600 180
rect 4800 170 4900 180
rect 6150 170 6250 180
rect 7050 170 7250 180
rect 8850 170 8900 180
rect 9000 170 9100 180
rect 9150 170 9200 180
rect 9300 170 9350 180
rect 9750 170 9800 180
rect 9850 170 9990 180
rect 0 160 100 170
rect 200 160 350 170
rect 450 160 1000 170
rect 4150 160 4600 170
rect 4800 160 4900 170
rect 6150 160 6250 170
rect 7050 160 7250 170
rect 8850 160 8900 170
rect 9000 160 9100 170
rect 9150 160 9200 170
rect 9300 160 9350 170
rect 9750 160 9800 170
rect 9850 160 9990 170
rect 0 150 100 160
rect 200 150 350 160
rect 450 150 1000 160
rect 4150 150 4600 160
rect 4800 150 4900 160
rect 6150 150 6250 160
rect 7050 150 7250 160
rect 8850 150 8900 160
rect 9000 150 9100 160
rect 9150 150 9200 160
rect 9300 150 9350 160
rect 9750 150 9800 160
rect 9850 150 9990 160
rect 100 140 150 150
rect 700 140 750 150
rect 900 140 1000 150
rect 4500 140 4850 150
rect 4900 140 4950 150
rect 5000 140 5050 150
rect 6150 140 6250 150
rect 7100 140 7250 150
rect 8800 140 8850 150
rect 8900 140 8950 150
rect 9150 140 9200 150
rect 9900 140 9990 150
rect 100 130 150 140
rect 700 130 750 140
rect 900 130 1000 140
rect 4500 130 4850 140
rect 4900 130 4950 140
rect 5000 130 5050 140
rect 6150 130 6250 140
rect 7100 130 7250 140
rect 8800 130 8850 140
rect 8900 130 8950 140
rect 9150 130 9200 140
rect 9900 130 9990 140
rect 100 120 150 130
rect 700 120 750 130
rect 900 120 1000 130
rect 4500 120 4850 130
rect 4900 120 4950 130
rect 5000 120 5050 130
rect 6150 120 6250 130
rect 7100 120 7250 130
rect 8800 120 8850 130
rect 8900 120 8950 130
rect 9150 120 9200 130
rect 9900 120 9990 130
rect 100 110 150 120
rect 700 110 750 120
rect 900 110 1000 120
rect 4500 110 4850 120
rect 4900 110 4950 120
rect 5000 110 5050 120
rect 6150 110 6250 120
rect 7100 110 7250 120
rect 8800 110 8850 120
rect 8900 110 8950 120
rect 9150 110 9200 120
rect 9900 110 9990 120
rect 100 100 150 110
rect 700 100 750 110
rect 900 100 1000 110
rect 4500 100 4850 110
rect 4900 100 4950 110
rect 5000 100 5050 110
rect 6150 100 6250 110
rect 7100 100 7250 110
rect 8800 100 8850 110
rect 8900 100 8950 110
rect 9150 100 9200 110
rect 9900 100 9990 110
rect 100 90 150 100
rect 950 90 1000 100
rect 4600 90 4800 100
rect 4900 90 4950 100
rect 6150 90 6300 100
rect 7200 90 7250 100
rect 8750 90 8800 100
rect 9000 90 9050 100
rect 9150 90 9200 100
rect 9400 90 9450 100
rect 9900 90 9990 100
rect 100 80 150 90
rect 950 80 1000 90
rect 4600 80 4800 90
rect 4900 80 4950 90
rect 6150 80 6300 90
rect 7200 80 7250 90
rect 8750 80 8800 90
rect 9000 80 9050 90
rect 9150 80 9200 90
rect 9400 80 9450 90
rect 9900 80 9990 90
rect 100 70 150 80
rect 950 70 1000 80
rect 4600 70 4800 80
rect 4900 70 4950 80
rect 6150 70 6300 80
rect 7200 70 7250 80
rect 8750 70 8800 80
rect 9000 70 9050 80
rect 9150 70 9200 80
rect 9400 70 9450 80
rect 9900 70 9990 80
rect 100 60 150 70
rect 950 60 1000 70
rect 4600 60 4800 70
rect 4900 60 4950 70
rect 6150 60 6300 70
rect 7200 60 7250 70
rect 8750 60 8800 70
rect 9000 60 9050 70
rect 9150 60 9200 70
rect 9400 60 9450 70
rect 9900 60 9990 70
rect 100 50 150 60
rect 950 50 1000 60
rect 4600 50 4800 60
rect 4900 50 4950 60
rect 6150 50 6300 60
rect 7200 50 7250 60
rect 8750 50 8800 60
rect 9000 50 9050 60
rect 9150 50 9200 60
rect 9400 50 9450 60
rect 9900 50 9990 60
rect 100 40 150 50
rect 950 40 1000 50
rect 4350 40 4400 50
rect 4650 40 4750 50
rect 4900 40 4950 50
rect 6150 40 6350 50
rect 7200 40 7250 50
rect 8600 40 8650 50
rect 8700 40 8750 50
rect 8900 40 8950 50
rect 9000 40 9050 50
rect 9150 40 9200 50
rect 9450 40 9500 50
rect 9750 40 9800 50
rect 9900 40 9950 50
rect 100 30 150 40
rect 950 30 1000 40
rect 4350 30 4400 40
rect 4650 30 4750 40
rect 4900 30 4950 40
rect 6150 30 6350 40
rect 7200 30 7250 40
rect 8600 30 8650 40
rect 8700 30 8750 40
rect 8900 30 8950 40
rect 9000 30 9050 40
rect 9150 30 9200 40
rect 9450 30 9500 40
rect 9750 30 9800 40
rect 9900 30 9950 40
rect 100 20 150 30
rect 950 20 1000 30
rect 4350 20 4400 30
rect 4650 20 4750 30
rect 4900 20 4950 30
rect 6150 20 6350 30
rect 7200 20 7250 30
rect 8600 20 8650 30
rect 8700 20 8750 30
rect 8900 20 8950 30
rect 9000 20 9050 30
rect 9150 20 9200 30
rect 9450 20 9500 30
rect 9750 20 9800 30
rect 9900 20 9950 30
rect 100 10 150 20
rect 950 10 1000 20
rect 4350 10 4400 20
rect 4650 10 4750 20
rect 4900 10 4950 20
rect 6150 10 6350 20
rect 7200 10 7250 20
rect 8600 10 8650 20
rect 8700 10 8750 20
rect 8900 10 8950 20
rect 9000 10 9050 20
rect 9150 10 9200 20
rect 9450 10 9500 20
rect 9750 10 9800 20
rect 9900 10 9950 20
rect 100 0 150 10
rect 950 0 1000 10
rect 4350 0 4400 10
rect 4650 0 4750 10
rect 4900 0 4950 10
rect 6150 0 6350 10
rect 7200 0 7250 10
rect 8600 0 8650 10
rect 8700 0 8750 10
rect 8900 0 8950 10
rect 9000 0 9050 10
rect 9150 0 9200 10
rect 9450 0 9500 10
rect 9750 0 9800 10
rect 9900 0 9950 10
<< metal4 >>
rect 2100 7490 2150 7500
rect 3700 7490 3850 7500
rect 9550 7490 9650 7500
rect 2100 7480 2150 7490
rect 3700 7480 3850 7490
rect 9550 7480 9650 7490
rect 2100 7470 2150 7480
rect 3700 7470 3850 7480
rect 9550 7470 9650 7480
rect 2100 7460 2150 7470
rect 3700 7460 3850 7470
rect 9550 7460 9650 7470
rect 2100 7450 2150 7460
rect 3700 7450 3850 7460
rect 9550 7450 9650 7460
rect 2050 7440 2100 7450
rect 3550 7440 3600 7450
rect 3650 7440 3700 7450
rect 3800 7440 3850 7450
rect 9550 7440 9600 7450
rect 2050 7430 2100 7440
rect 3550 7430 3600 7440
rect 3650 7430 3700 7440
rect 3800 7430 3850 7440
rect 9550 7430 9600 7440
rect 2050 7420 2100 7430
rect 3550 7420 3600 7430
rect 3650 7420 3700 7430
rect 3800 7420 3850 7430
rect 9550 7420 9600 7430
rect 2050 7410 2100 7420
rect 3550 7410 3600 7420
rect 3650 7410 3700 7420
rect 3800 7410 3850 7420
rect 9550 7410 9600 7420
rect 2050 7400 2100 7410
rect 3550 7400 3600 7410
rect 3650 7400 3700 7410
rect 3800 7400 3850 7410
rect 9550 7400 9600 7410
rect 3600 7390 3650 7400
rect 3850 7390 3900 7400
rect 9550 7390 9600 7400
rect 3600 7380 3650 7390
rect 3850 7380 3900 7390
rect 9550 7380 9600 7390
rect 3600 7370 3650 7380
rect 3850 7370 3900 7380
rect 9550 7370 9600 7380
rect 3600 7360 3650 7370
rect 3850 7360 3900 7370
rect 9550 7360 9600 7370
rect 3600 7350 3650 7360
rect 3850 7350 3900 7360
rect 9550 7350 9600 7360
rect 2000 7340 2050 7350
rect 3350 7340 3400 7350
rect 3850 7340 3900 7350
rect 9550 7340 9600 7350
rect 2000 7330 2050 7340
rect 3350 7330 3400 7340
rect 3850 7330 3900 7340
rect 9550 7330 9600 7340
rect 2000 7320 2050 7330
rect 3350 7320 3400 7330
rect 3850 7320 3900 7330
rect 9550 7320 9600 7330
rect 2000 7310 2050 7320
rect 3350 7310 3400 7320
rect 3850 7310 3900 7320
rect 9550 7310 9600 7320
rect 2000 7300 2050 7310
rect 3350 7300 3400 7310
rect 3850 7300 3900 7310
rect 9550 7300 9600 7310
rect 1950 7290 2000 7300
rect 3400 7290 3450 7300
rect 3800 7290 3900 7300
rect 9550 7290 9600 7300
rect 1950 7280 2000 7290
rect 3400 7280 3450 7290
rect 3800 7280 3900 7290
rect 9550 7280 9600 7290
rect 1950 7270 2000 7280
rect 3400 7270 3450 7280
rect 3800 7270 3900 7280
rect 9550 7270 9600 7280
rect 1950 7260 2000 7270
rect 3400 7260 3450 7270
rect 3800 7260 3900 7270
rect 9550 7260 9600 7270
rect 1950 7250 2000 7260
rect 3400 7250 3450 7260
rect 3800 7250 3900 7260
rect 9550 7250 9600 7260
rect 3800 7240 3850 7250
rect 3900 7240 3950 7250
rect 9550 7240 9600 7250
rect 3800 7230 3850 7240
rect 3900 7230 3950 7240
rect 9550 7230 9600 7240
rect 3800 7220 3850 7230
rect 3900 7220 3950 7230
rect 9550 7220 9600 7230
rect 3800 7210 3850 7220
rect 3900 7210 3950 7220
rect 9550 7210 9600 7220
rect 3800 7200 3850 7210
rect 3900 7200 3950 7210
rect 9550 7200 9600 7210
rect 1900 7190 1950 7200
rect 3400 7190 3450 7200
rect 3900 7190 3950 7200
rect 9550 7190 9600 7200
rect 1900 7180 1950 7190
rect 3400 7180 3450 7190
rect 3900 7180 3950 7190
rect 9550 7180 9600 7190
rect 1900 7170 1950 7180
rect 3400 7170 3450 7180
rect 3900 7170 3950 7180
rect 9550 7170 9600 7180
rect 1900 7160 1950 7170
rect 3400 7160 3450 7170
rect 3900 7160 3950 7170
rect 9550 7160 9600 7170
rect 1900 7150 1950 7160
rect 3400 7150 3450 7160
rect 3900 7150 3950 7160
rect 9550 7150 9600 7160
rect 3450 7140 3550 7150
rect 3700 7140 3800 7150
rect 9550 7140 9600 7150
rect 3450 7130 3550 7140
rect 3700 7130 3800 7140
rect 9550 7130 9600 7140
rect 3450 7120 3550 7130
rect 3700 7120 3800 7130
rect 9550 7120 9600 7130
rect 3450 7110 3550 7120
rect 3700 7110 3800 7120
rect 9550 7110 9600 7120
rect 3450 7100 3550 7110
rect 3700 7100 3800 7110
rect 9550 7100 9600 7110
rect 3550 7090 3650 7100
rect 3950 7090 4000 7100
rect 9550 7090 9600 7100
rect 3550 7080 3650 7090
rect 3950 7080 4000 7090
rect 9550 7080 9600 7090
rect 3550 7070 3650 7080
rect 3950 7070 4000 7080
rect 9550 7070 9600 7080
rect 3550 7060 3650 7070
rect 3950 7060 4000 7070
rect 9550 7060 9600 7070
rect 3550 7050 3650 7060
rect 3950 7050 4000 7060
rect 9550 7050 9600 7060
rect 3550 7040 3650 7050
rect 3750 7040 3800 7050
rect 3950 7040 4000 7050
rect 9550 7040 9600 7050
rect 3550 7030 3650 7040
rect 3750 7030 3800 7040
rect 3950 7030 4000 7040
rect 9550 7030 9600 7040
rect 3550 7020 3650 7030
rect 3750 7020 3800 7030
rect 3950 7020 4000 7030
rect 9550 7020 9600 7030
rect 3550 7010 3650 7020
rect 3750 7010 3800 7020
rect 3950 7010 4000 7020
rect 9550 7010 9600 7020
rect 3550 7000 3650 7010
rect 3750 7000 3800 7010
rect 3950 7000 4000 7010
rect 9550 7000 9600 7010
rect 1900 6990 1950 7000
rect 3700 6990 3850 7000
rect 3950 6990 4000 7000
rect 9550 6990 9600 7000
rect 1900 6980 1950 6990
rect 3700 6980 3850 6990
rect 3950 6980 4000 6990
rect 9550 6980 9600 6990
rect 1900 6970 1950 6980
rect 3700 6970 3850 6980
rect 3950 6970 4000 6980
rect 9550 6970 9600 6980
rect 1900 6960 1950 6970
rect 3700 6960 3850 6970
rect 3950 6960 4000 6970
rect 9550 6960 9600 6970
rect 1900 6950 1950 6960
rect 3700 6950 3850 6960
rect 3950 6950 4000 6960
rect 9550 6950 9600 6960
rect 1850 6940 1900 6950
rect 3250 6940 3400 6950
rect 3900 6940 4000 6950
rect 1850 6930 1900 6940
rect 3250 6930 3400 6940
rect 3900 6930 4000 6940
rect 1850 6920 1900 6930
rect 3250 6920 3400 6930
rect 3900 6920 4000 6930
rect 1850 6910 1900 6920
rect 3250 6910 3400 6920
rect 3900 6910 4000 6920
rect 1850 6900 1900 6910
rect 3250 6900 3400 6910
rect 3900 6900 4000 6910
rect 1850 6890 1900 6900
rect 3250 6890 3400 6900
rect 3450 6890 3500 6900
rect 3900 6890 4000 6900
rect 9550 6890 9600 6900
rect 1850 6880 1900 6890
rect 3250 6880 3400 6890
rect 3450 6880 3500 6890
rect 3900 6880 4000 6890
rect 9550 6880 9600 6890
rect 1850 6870 1900 6880
rect 3250 6870 3400 6880
rect 3450 6870 3500 6880
rect 3900 6870 4000 6880
rect 9550 6870 9600 6880
rect 1850 6860 1900 6870
rect 3250 6860 3400 6870
rect 3450 6860 3500 6870
rect 3900 6860 4000 6870
rect 9550 6860 9600 6870
rect 1850 6850 1900 6860
rect 3250 6850 3400 6860
rect 3450 6850 3500 6860
rect 3900 6850 4000 6860
rect 9550 6850 9600 6860
rect 1850 6840 1900 6850
rect 3100 6840 3450 6850
rect 3550 6840 3600 6850
rect 3900 6840 4000 6850
rect 9550 6840 9600 6850
rect 1850 6830 1900 6840
rect 3100 6830 3450 6840
rect 3550 6830 3600 6840
rect 3900 6830 4000 6840
rect 9550 6830 9600 6840
rect 1850 6820 1900 6830
rect 3100 6820 3450 6830
rect 3550 6820 3600 6830
rect 3900 6820 4000 6830
rect 9550 6820 9600 6830
rect 1850 6810 1900 6820
rect 3100 6810 3450 6820
rect 3550 6810 3600 6820
rect 3900 6810 4000 6820
rect 9550 6810 9600 6820
rect 1850 6800 1900 6810
rect 3100 6800 3450 6810
rect 3550 6800 3600 6810
rect 3900 6800 4000 6810
rect 9550 6800 9600 6810
rect 3050 6790 3350 6800
rect 3650 6790 3700 6800
rect 9550 6790 9600 6800
rect 3050 6780 3350 6790
rect 3650 6780 3700 6790
rect 9550 6780 9600 6790
rect 3050 6770 3350 6780
rect 3650 6770 3700 6780
rect 9550 6770 9600 6780
rect 3050 6760 3350 6770
rect 3650 6760 3700 6770
rect 9550 6760 9600 6770
rect 3050 6750 3350 6760
rect 3650 6750 3700 6760
rect 9550 6750 9600 6760
rect 2350 6740 2450 6750
rect 3300 6740 3450 6750
rect 3700 6740 3750 6750
rect 3950 6740 4000 6750
rect 9500 6740 9550 6750
rect 2350 6730 2450 6740
rect 3300 6730 3450 6740
rect 3700 6730 3750 6740
rect 3950 6730 4000 6740
rect 9500 6730 9550 6740
rect 2350 6720 2450 6730
rect 3300 6720 3450 6730
rect 3700 6720 3750 6730
rect 3950 6720 4000 6730
rect 9500 6720 9550 6730
rect 2350 6710 2450 6720
rect 3300 6710 3450 6720
rect 3700 6710 3750 6720
rect 3950 6710 4000 6720
rect 9500 6710 9550 6720
rect 2350 6700 2450 6710
rect 3300 6700 3450 6710
rect 3700 6700 3750 6710
rect 3950 6700 4000 6710
rect 9500 6700 9550 6710
rect 1800 6690 1850 6700
rect 2250 6690 2300 6700
rect 2450 6690 2500 6700
rect 3500 6690 3550 6700
rect 3950 6690 4000 6700
rect 9550 6690 9600 6700
rect 9950 6690 9990 6700
rect 1800 6680 1850 6690
rect 2250 6680 2300 6690
rect 2450 6680 2500 6690
rect 3500 6680 3550 6690
rect 3950 6680 4000 6690
rect 9550 6680 9600 6690
rect 9950 6680 9990 6690
rect 1800 6670 1850 6680
rect 2250 6670 2300 6680
rect 2450 6670 2500 6680
rect 3500 6670 3550 6680
rect 3950 6670 4000 6680
rect 9550 6670 9600 6680
rect 9950 6670 9990 6680
rect 1800 6660 1850 6670
rect 2250 6660 2300 6670
rect 2450 6660 2500 6670
rect 3500 6660 3550 6670
rect 3950 6660 4000 6670
rect 9550 6660 9600 6670
rect 9950 6660 9990 6670
rect 1800 6650 1850 6660
rect 2250 6650 2300 6660
rect 2450 6650 2500 6660
rect 3500 6650 3550 6660
rect 3950 6650 4000 6660
rect 9550 6650 9600 6660
rect 9950 6650 9990 6660
rect 1600 6640 1650 6650
rect 1700 6640 1750 6650
rect 2500 6640 2550 6650
rect 3650 6640 3700 6650
rect 3950 6640 4000 6650
rect 9450 6640 9500 6650
rect 9550 6640 9600 6650
rect 9800 6640 9850 6650
rect 1600 6630 1650 6640
rect 1700 6630 1750 6640
rect 2500 6630 2550 6640
rect 3650 6630 3700 6640
rect 3950 6630 4000 6640
rect 9450 6630 9500 6640
rect 9550 6630 9600 6640
rect 9800 6630 9850 6640
rect 1600 6620 1650 6630
rect 1700 6620 1750 6630
rect 2500 6620 2550 6630
rect 3650 6620 3700 6630
rect 3950 6620 4000 6630
rect 9450 6620 9500 6630
rect 9550 6620 9600 6630
rect 9800 6620 9850 6630
rect 1600 6610 1650 6620
rect 1700 6610 1750 6620
rect 2500 6610 2550 6620
rect 3650 6610 3700 6620
rect 3950 6610 4000 6620
rect 9450 6610 9500 6620
rect 9550 6610 9600 6620
rect 9800 6610 9850 6620
rect 1600 6600 1650 6610
rect 1700 6600 1750 6610
rect 2500 6600 2550 6610
rect 3650 6600 3700 6610
rect 3950 6600 4000 6610
rect 9450 6600 9500 6610
rect 9550 6600 9600 6610
rect 9800 6600 9850 6610
rect 1500 6590 1550 6600
rect 1650 6590 1750 6600
rect 2150 6590 2250 6600
rect 2550 6590 2600 6600
rect 3750 6590 3800 6600
rect 6000 6590 6450 6600
rect 9450 6590 9700 6600
rect 1500 6580 1550 6590
rect 1650 6580 1750 6590
rect 2150 6580 2250 6590
rect 2550 6580 2600 6590
rect 3750 6580 3800 6590
rect 6000 6580 6450 6590
rect 9450 6580 9700 6590
rect 1500 6570 1550 6580
rect 1650 6570 1750 6580
rect 2150 6570 2250 6580
rect 2550 6570 2600 6580
rect 3750 6570 3800 6580
rect 6000 6570 6450 6580
rect 9450 6570 9700 6580
rect 1500 6560 1550 6570
rect 1650 6560 1750 6570
rect 2150 6560 2250 6570
rect 2550 6560 2600 6570
rect 3750 6560 3800 6570
rect 6000 6560 6450 6570
rect 9450 6560 9700 6570
rect 1500 6550 1550 6560
rect 1650 6550 1750 6560
rect 2150 6550 2250 6560
rect 2550 6550 2600 6560
rect 3750 6550 3800 6560
rect 6000 6550 6450 6560
rect 9450 6550 9700 6560
rect 1300 6540 1350 6550
rect 2500 6540 2550 6550
rect 3850 6540 3900 6550
rect 4000 6540 4050 6550
rect 5950 6540 6150 6550
rect 6600 6540 6650 6550
rect 9900 6540 9990 6550
rect 1300 6530 1350 6540
rect 2500 6530 2550 6540
rect 3850 6530 3900 6540
rect 4000 6530 4050 6540
rect 5950 6530 6150 6540
rect 6600 6530 6650 6540
rect 9900 6530 9990 6540
rect 1300 6520 1350 6530
rect 2500 6520 2550 6530
rect 3850 6520 3900 6530
rect 4000 6520 4050 6530
rect 5950 6520 6150 6530
rect 6600 6520 6650 6530
rect 9900 6520 9990 6530
rect 1300 6510 1350 6520
rect 2500 6510 2550 6520
rect 3850 6510 3900 6520
rect 4000 6510 4050 6520
rect 5950 6510 6150 6520
rect 6600 6510 6650 6520
rect 9900 6510 9990 6520
rect 1300 6500 1350 6510
rect 2500 6500 2550 6510
rect 3850 6500 3900 6510
rect 4000 6500 4050 6510
rect 5950 6500 6150 6510
rect 6600 6500 6650 6510
rect 9900 6500 9990 6510
rect 1200 6490 1250 6500
rect 2250 6490 2300 6500
rect 2350 6490 2400 6500
rect 3900 6490 4050 6500
rect 5800 6490 6050 6500
rect 6650 6490 6750 6500
rect 9700 6490 9800 6500
rect 1200 6480 1250 6490
rect 2250 6480 2300 6490
rect 2350 6480 2400 6490
rect 3900 6480 4050 6490
rect 5800 6480 6050 6490
rect 6650 6480 6750 6490
rect 9700 6480 9800 6490
rect 1200 6470 1250 6480
rect 2250 6470 2300 6480
rect 2350 6470 2400 6480
rect 3900 6470 4050 6480
rect 5800 6470 6050 6480
rect 6650 6470 6750 6480
rect 9700 6470 9800 6480
rect 1200 6460 1250 6470
rect 2250 6460 2300 6470
rect 2350 6460 2400 6470
rect 3900 6460 4050 6470
rect 5800 6460 6050 6470
rect 6650 6460 6750 6470
rect 9700 6460 9800 6470
rect 1200 6450 1250 6460
rect 2250 6450 2300 6460
rect 2350 6450 2400 6460
rect 3900 6450 4050 6460
rect 5800 6450 6050 6460
rect 6650 6450 6750 6460
rect 9700 6450 9800 6460
rect 1200 6440 1250 6450
rect 1650 6440 1750 6450
rect 2100 6440 2150 6450
rect 2300 6440 2400 6450
rect 4000 6440 4050 6450
rect 5700 6440 6050 6450
rect 6700 6440 6800 6450
rect 9600 6440 9650 6450
rect 1200 6430 1250 6440
rect 1650 6430 1750 6440
rect 2100 6430 2150 6440
rect 2300 6430 2400 6440
rect 4000 6430 4050 6440
rect 5700 6430 6050 6440
rect 6700 6430 6800 6440
rect 9600 6430 9650 6440
rect 1200 6420 1250 6430
rect 1650 6420 1750 6430
rect 2100 6420 2150 6430
rect 2300 6420 2400 6430
rect 4000 6420 4050 6430
rect 5700 6420 6050 6430
rect 6700 6420 6800 6430
rect 9600 6420 9650 6430
rect 1200 6410 1250 6420
rect 1650 6410 1750 6420
rect 2100 6410 2150 6420
rect 2300 6410 2400 6420
rect 4000 6410 4050 6420
rect 5700 6410 6050 6420
rect 6700 6410 6800 6420
rect 9600 6410 9650 6420
rect 1200 6400 1250 6410
rect 1650 6400 1750 6410
rect 2100 6400 2150 6410
rect 2300 6400 2400 6410
rect 4000 6400 4050 6410
rect 5700 6400 6050 6410
rect 6700 6400 6800 6410
rect 9600 6400 9650 6410
rect 1200 6390 1400 6400
rect 1650 6390 1700 6400
rect 1850 6390 2100 6400
rect 2350 6390 2400 6400
rect 4050 6390 4100 6400
rect 5650 6390 5800 6400
rect 5850 6390 6150 6400
rect 6250 6390 6350 6400
rect 6800 6390 6850 6400
rect 9600 6390 9650 6400
rect 1200 6380 1400 6390
rect 1650 6380 1700 6390
rect 1850 6380 2100 6390
rect 2350 6380 2400 6390
rect 4050 6380 4100 6390
rect 5650 6380 5800 6390
rect 5850 6380 6150 6390
rect 6250 6380 6350 6390
rect 6800 6380 6850 6390
rect 9600 6380 9650 6390
rect 1200 6370 1400 6380
rect 1650 6370 1700 6380
rect 1850 6370 2100 6380
rect 2350 6370 2400 6380
rect 4050 6370 4100 6380
rect 5650 6370 5800 6380
rect 5850 6370 6150 6380
rect 6250 6370 6350 6380
rect 6800 6370 6850 6380
rect 9600 6370 9650 6380
rect 1200 6360 1400 6370
rect 1650 6360 1700 6370
rect 1850 6360 2100 6370
rect 2350 6360 2400 6370
rect 4050 6360 4100 6370
rect 5650 6360 5800 6370
rect 5850 6360 6150 6370
rect 6250 6360 6350 6370
rect 6800 6360 6850 6370
rect 9600 6360 9650 6370
rect 1200 6350 1400 6360
rect 1650 6350 1700 6360
rect 1850 6350 2100 6360
rect 2350 6350 2400 6360
rect 4050 6350 4100 6360
rect 5650 6350 5800 6360
rect 5850 6350 6150 6360
rect 6250 6350 6350 6360
rect 6800 6350 6850 6360
rect 9600 6350 9650 6360
rect 1200 6340 1300 6350
rect 1850 6340 1900 6350
rect 5400 6340 5500 6350
rect 5800 6340 5900 6350
rect 6350 6340 6400 6350
rect 6800 6340 6850 6350
rect 9350 6340 9500 6350
rect 9600 6340 9650 6350
rect 1200 6330 1300 6340
rect 1850 6330 1900 6340
rect 5400 6330 5500 6340
rect 5800 6330 5900 6340
rect 6350 6330 6400 6340
rect 6800 6330 6850 6340
rect 9350 6330 9500 6340
rect 9600 6330 9650 6340
rect 1200 6320 1300 6330
rect 1850 6320 1900 6330
rect 5400 6320 5500 6330
rect 5800 6320 5900 6330
rect 6350 6320 6400 6330
rect 6800 6320 6850 6330
rect 9350 6320 9500 6330
rect 9600 6320 9650 6330
rect 1200 6310 1300 6320
rect 1850 6310 1900 6320
rect 5400 6310 5500 6320
rect 5800 6310 5900 6320
rect 6350 6310 6400 6320
rect 6800 6310 6850 6320
rect 9350 6310 9500 6320
rect 9600 6310 9650 6320
rect 1200 6300 1300 6310
rect 1850 6300 1900 6310
rect 5400 6300 5500 6310
rect 5800 6300 5900 6310
rect 6350 6300 6400 6310
rect 6800 6300 6850 6310
rect 9350 6300 9500 6310
rect 9600 6300 9650 6310
rect 1200 6290 1250 6300
rect 1300 6290 1400 6300
rect 5300 6290 5350 6300
rect 5650 6290 5800 6300
rect 6450 6290 6500 6300
rect 9250 6290 9350 6300
rect 9400 6290 9650 6300
rect 1200 6280 1250 6290
rect 1300 6280 1400 6290
rect 5300 6280 5350 6290
rect 5650 6280 5800 6290
rect 6450 6280 6500 6290
rect 9250 6280 9350 6290
rect 9400 6280 9650 6290
rect 1200 6270 1250 6280
rect 1300 6270 1400 6280
rect 5300 6270 5350 6280
rect 5650 6270 5800 6280
rect 6450 6270 6500 6280
rect 9250 6270 9350 6280
rect 9400 6270 9650 6280
rect 1200 6260 1250 6270
rect 1300 6260 1400 6270
rect 5300 6260 5350 6270
rect 5650 6260 5800 6270
rect 6450 6260 6500 6270
rect 9250 6260 9350 6270
rect 9400 6260 9650 6270
rect 1200 6250 1250 6260
rect 1300 6250 1400 6260
rect 5300 6250 5350 6260
rect 5650 6250 5800 6260
rect 6450 6250 6500 6260
rect 9250 6250 9350 6260
rect 9400 6250 9650 6260
rect 1150 6240 1250 6250
rect 5550 6240 5600 6250
rect 6500 6240 6550 6250
rect 6850 6240 6900 6250
rect 9250 6240 9400 6250
rect 9800 6240 9850 6250
rect 9900 6240 9950 6250
rect 1150 6230 1250 6240
rect 5550 6230 5600 6240
rect 6500 6230 6550 6240
rect 6850 6230 6900 6240
rect 9250 6230 9400 6240
rect 9800 6230 9850 6240
rect 9900 6230 9950 6240
rect 1150 6220 1250 6230
rect 5550 6220 5600 6230
rect 6500 6220 6550 6230
rect 6850 6220 6900 6230
rect 9250 6220 9400 6230
rect 9800 6220 9850 6230
rect 9900 6220 9950 6230
rect 1150 6210 1250 6220
rect 5550 6210 5600 6220
rect 6500 6210 6550 6220
rect 6850 6210 6900 6220
rect 9250 6210 9400 6220
rect 9800 6210 9850 6220
rect 9900 6210 9950 6220
rect 1150 6200 1250 6210
rect 5550 6200 5600 6210
rect 6500 6200 6550 6210
rect 6850 6200 6900 6210
rect 9250 6200 9400 6210
rect 9800 6200 9850 6210
rect 9900 6200 9950 6210
rect 1150 6190 1250 6200
rect 1750 6190 1800 6200
rect 4250 6190 4300 6200
rect 5250 6190 5300 6200
rect 5500 6190 5550 6200
rect 6600 6190 6650 6200
rect 6900 6190 6950 6200
rect 9200 6190 9250 6200
rect 9800 6190 9850 6200
rect 1150 6180 1250 6190
rect 1750 6180 1800 6190
rect 4250 6180 4300 6190
rect 5250 6180 5300 6190
rect 5500 6180 5550 6190
rect 6600 6180 6650 6190
rect 6900 6180 6950 6190
rect 9200 6180 9250 6190
rect 9800 6180 9850 6190
rect 1150 6170 1250 6180
rect 1750 6170 1800 6180
rect 4250 6170 4300 6180
rect 5250 6170 5300 6180
rect 5500 6170 5550 6180
rect 6600 6170 6650 6180
rect 6900 6170 6950 6180
rect 9200 6170 9250 6180
rect 9800 6170 9850 6180
rect 1150 6160 1250 6170
rect 1750 6160 1800 6170
rect 4250 6160 4300 6170
rect 5250 6160 5300 6170
rect 5500 6160 5550 6170
rect 6600 6160 6650 6170
rect 6900 6160 6950 6170
rect 9200 6160 9250 6170
rect 9800 6160 9850 6170
rect 1150 6150 1250 6160
rect 1750 6150 1800 6160
rect 4250 6150 4300 6160
rect 5250 6150 5300 6160
rect 5500 6150 5550 6160
rect 6600 6150 6650 6160
rect 6900 6150 6950 6160
rect 9200 6150 9250 6160
rect 9800 6150 9850 6160
rect 1100 6140 1250 6150
rect 1700 6140 1800 6150
rect 2400 6140 2450 6150
rect 5200 6140 5250 6150
rect 6650 6140 6700 6150
rect 6950 6140 7000 6150
rect 9100 6140 9150 6150
rect 9850 6140 9950 6150
rect 1100 6130 1250 6140
rect 1700 6130 1800 6140
rect 2400 6130 2450 6140
rect 5200 6130 5250 6140
rect 6650 6130 6700 6140
rect 6950 6130 7000 6140
rect 9100 6130 9150 6140
rect 9850 6130 9950 6140
rect 1100 6120 1250 6130
rect 1700 6120 1800 6130
rect 2400 6120 2450 6130
rect 5200 6120 5250 6130
rect 6650 6120 6700 6130
rect 6950 6120 7000 6130
rect 9100 6120 9150 6130
rect 9850 6120 9950 6130
rect 1100 6110 1250 6120
rect 1700 6110 1800 6120
rect 2400 6110 2450 6120
rect 5200 6110 5250 6120
rect 6650 6110 6700 6120
rect 6950 6110 7000 6120
rect 9100 6110 9150 6120
rect 9850 6110 9950 6120
rect 1100 6100 1250 6110
rect 1700 6100 1800 6110
rect 2400 6100 2450 6110
rect 5200 6100 5250 6110
rect 6650 6100 6700 6110
rect 6950 6100 7000 6110
rect 9100 6100 9150 6110
rect 9850 6100 9950 6110
rect 1100 6090 1250 6100
rect 1700 6090 1800 6100
rect 3850 6090 3900 6100
rect 4300 6090 4350 6100
rect 5200 6090 5250 6100
rect 5400 6090 5450 6100
rect 6650 6090 6700 6100
rect 6950 6090 7000 6100
rect 8950 6090 9050 6100
rect 9350 6090 9500 6100
rect 9850 6090 9950 6100
rect 1100 6080 1250 6090
rect 1700 6080 1800 6090
rect 3850 6080 3900 6090
rect 4300 6080 4350 6090
rect 5200 6080 5250 6090
rect 5400 6080 5450 6090
rect 6650 6080 6700 6090
rect 6950 6080 7000 6090
rect 8950 6080 9050 6090
rect 9350 6080 9500 6090
rect 9850 6080 9950 6090
rect 1100 6070 1250 6080
rect 1700 6070 1800 6080
rect 3850 6070 3900 6080
rect 4300 6070 4350 6080
rect 5200 6070 5250 6080
rect 5400 6070 5450 6080
rect 6650 6070 6700 6080
rect 6950 6070 7000 6080
rect 8950 6070 9050 6080
rect 9350 6070 9500 6080
rect 9850 6070 9950 6080
rect 1100 6060 1250 6070
rect 1700 6060 1800 6070
rect 3850 6060 3900 6070
rect 4300 6060 4350 6070
rect 5200 6060 5250 6070
rect 5400 6060 5450 6070
rect 6650 6060 6700 6070
rect 6950 6060 7000 6070
rect 8950 6060 9050 6070
rect 9350 6060 9500 6070
rect 9850 6060 9950 6070
rect 1100 6050 1250 6060
rect 1700 6050 1800 6060
rect 3850 6050 3900 6060
rect 4300 6050 4350 6060
rect 5200 6050 5250 6060
rect 5400 6050 5450 6060
rect 6650 6050 6700 6060
rect 6950 6050 7000 6060
rect 8950 6050 9050 6060
rect 9350 6050 9500 6060
rect 9850 6050 9950 6060
rect 750 6040 850 6050
rect 900 6040 1150 6050
rect 1750 6040 1800 6050
rect 2450 6040 2500 6050
rect 3800 6040 3850 6050
rect 5150 6040 5200 6050
rect 6700 6040 6750 6050
rect 8750 6040 8850 6050
rect 9200 6040 9250 6050
rect 9350 6040 9500 6050
rect 9900 6040 9950 6050
rect 750 6030 850 6040
rect 900 6030 1150 6040
rect 1750 6030 1800 6040
rect 2450 6030 2500 6040
rect 3800 6030 3850 6040
rect 5150 6030 5200 6040
rect 6700 6030 6750 6040
rect 8750 6030 8850 6040
rect 9200 6030 9250 6040
rect 9350 6030 9500 6040
rect 9900 6030 9950 6040
rect 750 6020 850 6030
rect 900 6020 1150 6030
rect 1750 6020 1800 6030
rect 2450 6020 2500 6030
rect 3800 6020 3850 6030
rect 5150 6020 5200 6030
rect 6700 6020 6750 6030
rect 8750 6020 8850 6030
rect 9200 6020 9250 6030
rect 9350 6020 9500 6030
rect 9900 6020 9950 6030
rect 750 6010 850 6020
rect 900 6010 1150 6020
rect 1750 6010 1800 6020
rect 2450 6010 2500 6020
rect 3800 6010 3850 6020
rect 5150 6010 5200 6020
rect 6700 6010 6750 6020
rect 8750 6010 8850 6020
rect 9200 6010 9250 6020
rect 9350 6010 9500 6020
rect 9900 6010 9950 6020
rect 750 6000 850 6010
rect 900 6000 1150 6010
rect 1750 6000 1800 6010
rect 2450 6000 2500 6010
rect 3800 6000 3850 6010
rect 5150 6000 5200 6010
rect 6700 6000 6750 6010
rect 8750 6000 8850 6010
rect 9200 6000 9250 6010
rect 9350 6000 9500 6010
rect 9900 6000 9950 6010
rect 700 5990 800 6000
rect 1000 5990 1100 6000
rect 1750 5990 1800 6000
rect 4050 5990 4100 6000
rect 5350 5990 5400 6000
rect 6700 5990 6750 6000
rect 8600 5990 8700 6000
rect 9050 5990 9150 6000
rect 9200 5990 9250 6000
rect 9350 5990 9500 6000
rect 9900 5990 9990 6000
rect 700 5980 800 5990
rect 1000 5980 1100 5990
rect 1750 5980 1800 5990
rect 4050 5980 4100 5990
rect 5350 5980 5400 5990
rect 6700 5980 6750 5990
rect 8600 5980 8700 5990
rect 9050 5980 9150 5990
rect 9200 5980 9250 5990
rect 9350 5980 9500 5990
rect 9900 5980 9990 5990
rect 700 5970 800 5980
rect 1000 5970 1100 5980
rect 1750 5970 1800 5980
rect 4050 5970 4100 5980
rect 5350 5970 5400 5980
rect 6700 5970 6750 5980
rect 8600 5970 8700 5980
rect 9050 5970 9150 5980
rect 9200 5970 9250 5980
rect 9350 5970 9500 5980
rect 9900 5970 9990 5980
rect 700 5960 800 5970
rect 1000 5960 1100 5970
rect 1750 5960 1800 5970
rect 4050 5960 4100 5970
rect 5350 5960 5400 5970
rect 6700 5960 6750 5970
rect 8600 5960 8700 5970
rect 9050 5960 9150 5970
rect 9200 5960 9250 5970
rect 9350 5960 9500 5970
rect 9900 5960 9990 5970
rect 700 5950 800 5960
rect 1000 5950 1100 5960
rect 1750 5950 1800 5960
rect 4050 5950 4100 5960
rect 5350 5950 5400 5960
rect 6700 5950 6750 5960
rect 8600 5950 8700 5960
rect 9050 5950 9150 5960
rect 9200 5950 9250 5960
rect 9350 5950 9500 5960
rect 9900 5950 9990 5960
rect 650 5940 700 5950
rect 800 5940 850 5950
rect 900 5940 950 5950
rect 1750 5940 1800 5950
rect 2450 5940 2500 5950
rect 3750 5940 3800 5950
rect 3850 5940 3900 5950
rect 4150 5940 4200 5950
rect 5100 5940 5150 5950
rect 6750 5940 6800 5950
rect 7000 5940 7050 5950
rect 8450 5940 8550 5950
rect 8850 5940 8900 5950
rect 8950 5940 9000 5950
rect 9200 5940 9250 5950
rect 9900 5940 9950 5950
rect 650 5930 700 5940
rect 800 5930 850 5940
rect 900 5930 950 5940
rect 1750 5930 1800 5940
rect 2450 5930 2500 5940
rect 3750 5930 3800 5940
rect 3850 5930 3900 5940
rect 4150 5930 4200 5940
rect 5100 5930 5150 5940
rect 6750 5930 6800 5940
rect 7000 5930 7050 5940
rect 8450 5930 8550 5940
rect 8850 5930 8900 5940
rect 8950 5930 9000 5940
rect 9200 5930 9250 5940
rect 9900 5930 9950 5940
rect 650 5920 700 5930
rect 800 5920 850 5930
rect 900 5920 950 5930
rect 1750 5920 1800 5930
rect 2450 5920 2500 5930
rect 3750 5920 3800 5930
rect 3850 5920 3900 5930
rect 4150 5920 4200 5930
rect 5100 5920 5150 5930
rect 6750 5920 6800 5930
rect 7000 5920 7050 5930
rect 8450 5920 8550 5930
rect 8850 5920 8900 5930
rect 8950 5920 9000 5930
rect 9200 5920 9250 5930
rect 9900 5920 9950 5930
rect 650 5910 700 5920
rect 800 5910 850 5920
rect 900 5910 950 5920
rect 1750 5910 1800 5920
rect 2450 5910 2500 5920
rect 3750 5910 3800 5920
rect 3850 5910 3900 5920
rect 4150 5910 4200 5920
rect 5100 5910 5150 5920
rect 6750 5910 6800 5920
rect 7000 5910 7050 5920
rect 8450 5910 8550 5920
rect 8850 5910 8900 5920
rect 8950 5910 9000 5920
rect 9200 5910 9250 5920
rect 9900 5910 9950 5920
rect 650 5900 700 5910
rect 800 5900 850 5910
rect 900 5900 950 5910
rect 1750 5900 1800 5910
rect 2450 5900 2500 5910
rect 3750 5900 3800 5910
rect 3850 5900 3900 5910
rect 4150 5900 4200 5910
rect 5100 5900 5150 5910
rect 6750 5900 6800 5910
rect 7000 5900 7050 5910
rect 8450 5900 8550 5910
rect 8850 5900 8900 5910
rect 8950 5900 9000 5910
rect 9200 5900 9250 5910
rect 9900 5900 9950 5910
rect 600 5890 650 5900
rect 800 5890 950 5900
rect 1850 5890 1900 5900
rect 2300 5890 2550 5900
rect 3150 5890 3200 5900
rect 3750 5890 3800 5900
rect 3900 5890 3950 5900
rect 4250 5890 4300 5900
rect 6750 5890 6800 5900
rect 7000 5890 7050 5900
rect 8250 5890 8350 5900
rect 8650 5890 8750 5900
rect 8800 5890 8850 5900
rect 8900 5890 9000 5900
rect 9050 5890 9100 5900
rect 9200 5890 9300 5900
rect 9900 5890 9950 5900
rect 600 5880 650 5890
rect 800 5880 950 5890
rect 1850 5880 1900 5890
rect 2300 5880 2550 5890
rect 3150 5880 3200 5890
rect 3750 5880 3800 5890
rect 3900 5880 3950 5890
rect 4250 5880 4300 5890
rect 6750 5880 6800 5890
rect 7000 5880 7050 5890
rect 8250 5880 8350 5890
rect 8650 5880 8750 5890
rect 8800 5880 8850 5890
rect 8900 5880 9000 5890
rect 9050 5880 9100 5890
rect 9200 5880 9300 5890
rect 9900 5880 9950 5890
rect 600 5870 650 5880
rect 800 5870 950 5880
rect 1850 5870 1900 5880
rect 2300 5870 2550 5880
rect 3150 5870 3200 5880
rect 3750 5870 3800 5880
rect 3900 5870 3950 5880
rect 4250 5870 4300 5880
rect 6750 5870 6800 5880
rect 7000 5870 7050 5880
rect 8250 5870 8350 5880
rect 8650 5870 8750 5880
rect 8800 5870 8850 5880
rect 8900 5870 9000 5880
rect 9050 5870 9100 5880
rect 9200 5870 9300 5880
rect 9900 5870 9950 5880
rect 600 5860 650 5870
rect 800 5860 950 5870
rect 1850 5860 1900 5870
rect 2300 5860 2550 5870
rect 3150 5860 3200 5870
rect 3750 5860 3800 5870
rect 3900 5860 3950 5870
rect 4250 5860 4300 5870
rect 6750 5860 6800 5870
rect 7000 5860 7050 5870
rect 8250 5860 8350 5870
rect 8650 5860 8750 5870
rect 8800 5860 8850 5870
rect 8900 5860 9000 5870
rect 9050 5860 9100 5870
rect 9200 5860 9300 5870
rect 9900 5860 9950 5870
rect 600 5850 650 5860
rect 800 5850 950 5860
rect 1850 5850 1900 5860
rect 2300 5850 2550 5860
rect 3150 5850 3200 5860
rect 3750 5850 3800 5860
rect 3900 5850 3950 5860
rect 4250 5850 4300 5860
rect 6750 5850 6800 5860
rect 7000 5850 7050 5860
rect 8250 5850 8350 5860
rect 8650 5850 8750 5860
rect 8800 5850 8850 5860
rect 8900 5850 9000 5860
rect 9050 5850 9100 5860
rect 9200 5850 9300 5860
rect 9900 5850 9950 5860
rect 550 5840 600 5850
rect 750 5840 800 5850
rect 1850 5840 1900 5850
rect 2250 5840 2300 5850
rect 2350 5840 2600 5850
rect 3050 5840 3200 5850
rect 3850 5840 3950 5850
rect 6750 5840 6800 5850
rect 8100 5840 8200 5850
rect 8650 5840 8700 5850
rect 8800 5840 8850 5850
rect 8900 5840 8950 5850
rect 9000 5840 9050 5850
rect 550 5830 600 5840
rect 750 5830 800 5840
rect 1850 5830 1900 5840
rect 2250 5830 2300 5840
rect 2350 5830 2600 5840
rect 3050 5830 3200 5840
rect 3850 5830 3950 5840
rect 6750 5830 6800 5840
rect 8100 5830 8200 5840
rect 8650 5830 8700 5840
rect 8800 5830 8850 5840
rect 8900 5830 8950 5840
rect 9000 5830 9050 5840
rect 550 5820 600 5830
rect 750 5820 800 5830
rect 1850 5820 1900 5830
rect 2250 5820 2300 5830
rect 2350 5820 2600 5830
rect 3050 5820 3200 5830
rect 3850 5820 3950 5830
rect 6750 5820 6800 5830
rect 8100 5820 8200 5830
rect 8650 5820 8700 5830
rect 8800 5820 8850 5830
rect 8900 5820 8950 5830
rect 9000 5820 9050 5830
rect 550 5810 600 5820
rect 750 5810 800 5820
rect 1850 5810 1900 5820
rect 2250 5810 2300 5820
rect 2350 5810 2600 5820
rect 3050 5810 3200 5820
rect 3850 5810 3950 5820
rect 6750 5810 6800 5820
rect 8100 5810 8200 5820
rect 8650 5810 8700 5820
rect 8800 5810 8850 5820
rect 8900 5810 8950 5820
rect 9000 5810 9050 5820
rect 550 5800 600 5810
rect 750 5800 800 5810
rect 1850 5800 1900 5810
rect 2250 5800 2300 5810
rect 2350 5800 2600 5810
rect 3050 5800 3200 5810
rect 3850 5800 3950 5810
rect 6750 5800 6800 5810
rect 8100 5800 8200 5810
rect 8650 5800 8700 5810
rect 8800 5800 8850 5810
rect 8900 5800 8950 5810
rect 9000 5800 9050 5810
rect 550 5790 650 5800
rect 700 5790 800 5800
rect 1900 5790 1950 5800
rect 2200 5790 2250 5800
rect 2350 5790 2550 5800
rect 3000 5790 3100 5800
rect 3150 5790 3200 5800
rect 3900 5790 4000 5800
rect 5050 5790 5100 5800
rect 5300 5790 5350 5800
rect 7950 5790 8050 5800
rect 8700 5790 8750 5800
rect 8850 5790 8950 5800
rect 550 5780 650 5790
rect 700 5780 800 5790
rect 1900 5780 1950 5790
rect 2200 5780 2250 5790
rect 2350 5780 2550 5790
rect 3000 5780 3100 5790
rect 3150 5780 3200 5790
rect 3900 5780 4000 5790
rect 5050 5780 5100 5790
rect 5300 5780 5350 5790
rect 7950 5780 8050 5790
rect 8700 5780 8750 5790
rect 8850 5780 8950 5790
rect 550 5770 650 5780
rect 700 5770 800 5780
rect 1900 5770 1950 5780
rect 2200 5770 2250 5780
rect 2350 5770 2550 5780
rect 3000 5770 3100 5780
rect 3150 5770 3200 5780
rect 3900 5770 4000 5780
rect 5050 5770 5100 5780
rect 5300 5770 5350 5780
rect 7950 5770 8050 5780
rect 8700 5770 8750 5780
rect 8850 5770 8950 5780
rect 550 5760 650 5770
rect 700 5760 800 5770
rect 1900 5760 1950 5770
rect 2200 5760 2250 5770
rect 2350 5760 2550 5770
rect 3000 5760 3100 5770
rect 3150 5760 3200 5770
rect 3900 5760 4000 5770
rect 5050 5760 5100 5770
rect 5300 5760 5350 5770
rect 7950 5760 8050 5770
rect 8700 5760 8750 5770
rect 8850 5760 8950 5770
rect 550 5750 650 5760
rect 700 5750 800 5760
rect 1900 5750 1950 5760
rect 2200 5750 2250 5760
rect 2350 5750 2550 5760
rect 3000 5750 3100 5760
rect 3150 5750 3200 5760
rect 3900 5750 4000 5760
rect 5050 5750 5100 5760
rect 5300 5750 5350 5760
rect 7950 5750 8050 5760
rect 8700 5750 8750 5760
rect 8850 5750 8950 5760
rect 600 5740 800 5750
rect 1900 5740 1950 5750
rect 2300 5740 2500 5750
rect 2950 5740 3050 5750
rect 3150 5740 3200 5750
rect 4000 5740 4050 5750
rect 5050 5740 5100 5750
rect 5300 5740 5350 5750
rect 7750 5740 7900 5750
rect 8400 5740 8450 5750
rect 8700 5740 8750 5750
rect 9950 5740 9990 5750
rect 600 5730 800 5740
rect 1900 5730 1950 5740
rect 2300 5730 2500 5740
rect 2950 5730 3050 5740
rect 3150 5730 3200 5740
rect 4000 5730 4050 5740
rect 5050 5730 5100 5740
rect 5300 5730 5350 5740
rect 7750 5730 7900 5740
rect 8400 5730 8450 5740
rect 8700 5730 8750 5740
rect 9950 5730 9990 5740
rect 600 5720 800 5730
rect 1900 5720 1950 5730
rect 2300 5720 2500 5730
rect 2950 5720 3050 5730
rect 3150 5720 3200 5730
rect 4000 5720 4050 5730
rect 5050 5720 5100 5730
rect 5300 5720 5350 5730
rect 7750 5720 7900 5730
rect 8400 5720 8450 5730
rect 8700 5720 8750 5730
rect 9950 5720 9990 5730
rect 600 5710 800 5720
rect 1900 5710 1950 5720
rect 2300 5710 2500 5720
rect 2950 5710 3050 5720
rect 3150 5710 3200 5720
rect 4000 5710 4050 5720
rect 5050 5710 5100 5720
rect 5300 5710 5350 5720
rect 7750 5710 7900 5720
rect 8400 5710 8450 5720
rect 8700 5710 8750 5720
rect 9950 5710 9990 5720
rect 600 5700 800 5710
rect 1900 5700 1950 5710
rect 2300 5700 2500 5710
rect 2950 5700 3050 5710
rect 3150 5700 3200 5710
rect 4000 5700 4050 5710
rect 5050 5700 5100 5710
rect 5300 5700 5350 5710
rect 7750 5700 7900 5710
rect 8400 5700 8450 5710
rect 8700 5700 8750 5710
rect 9950 5700 9990 5710
rect 600 5690 650 5700
rect 750 5690 800 5700
rect 1950 5690 2000 5700
rect 2150 5690 2200 5700
rect 2300 5690 2450 5700
rect 2800 5690 2850 5700
rect 2900 5690 3000 5700
rect 3150 5690 3200 5700
rect 5050 5690 5100 5700
rect 6800 5690 6850 5700
rect 6950 5690 7000 5700
rect 7650 5690 7700 5700
rect 8100 5690 8300 5700
rect 8400 5690 8450 5700
rect 600 5680 650 5690
rect 750 5680 800 5690
rect 1950 5680 2000 5690
rect 2150 5680 2200 5690
rect 2300 5680 2450 5690
rect 2800 5680 2850 5690
rect 2900 5680 3000 5690
rect 3150 5680 3200 5690
rect 5050 5680 5100 5690
rect 6800 5680 6850 5690
rect 6950 5680 7000 5690
rect 7650 5680 7700 5690
rect 8100 5680 8300 5690
rect 8400 5680 8450 5690
rect 600 5670 650 5680
rect 750 5670 800 5680
rect 1950 5670 2000 5680
rect 2150 5670 2200 5680
rect 2300 5670 2450 5680
rect 2800 5670 2850 5680
rect 2900 5670 3000 5680
rect 3150 5670 3200 5680
rect 5050 5670 5100 5680
rect 6800 5670 6850 5680
rect 6950 5670 7000 5680
rect 7650 5670 7700 5680
rect 8100 5670 8300 5680
rect 8400 5670 8450 5680
rect 600 5660 650 5670
rect 750 5660 800 5670
rect 1950 5660 2000 5670
rect 2150 5660 2200 5670
rect 2300 5660 2450 5670
rect 2800 5660 2850 5670
rect 2900 5660 3000 5670
rect 3150 5660 3200 5670
rect 5050 5660 5100 5670
rect 6800 5660 6850 5670
rect 6950 5660 7000 5670
rect 7650 5660 7700 5670
rect 8100 5660 8300 5670
rect 8400 5660 8450 5670
rect 600 5650 650 5660
rect 750 5650 800 5660
rect 1950 5650 2000 5660
rect 2150 5650 2200 5660
rect 2300 5650 2450 5660
rect 2800 5650 2850 5660
rect 2900 5650 3000 5660
rect 3150 5650 3200 5660
rect 5050 5650 5100 5660
rect 6800 5650 6850 5660
rect 6950 5650 7000 5660
rect 7650 5650 7700 5660
rect 8100 5650 8300 5660
rect 8400 5650 8450 5660
rect 500 5640 750 5650
rect 1950 5640 2050 5650
rect 2100 5640 2150 5650
rect 2250 5640 2350 5650
rect 2400 5640 2450 5650
rect 2800 5640 2900 5650
rect 3150 5640 3200 5650
rect 3800 5640 3950 5650
rect 5050 5640 5100 5650
rect 5500 5640 5600 5650
rect 5800 5640 5950 5650
rect 6300 5640 6450 5650
rect 6950 5640 7000 5650
rect 7450 5640 7550 5650
rect 7850 5640 7900 5650
rect 8050 5640 8300 5650
rect 8400 5640 8500 5650
rect 500 5630 750 5640
rect 1950 5630 2050 5640
rect 2100 5630 2150 5640
rect 2250 5630 2350 5640
rect 2400 5630 2450 5640
rect 2800 5630 2900 5640
rect 3150 5630 3200 5640
rect 3800 5630 3950 5640
rect 5050 5630 5100 5640
rect 5500 5630 5600 5640
rect 5800 5630 5950 5640
rect 6300 5630 6450 5640
rect 6950 5630 7000 5640
rect 7450 5630 7550 5640
rect 7850 5630 7900 5640
rect 8050 5630 8300 5640
rect 8400 5630 8500 5640
rect 500 5620 750 5630
rect 1950 5620 2050 5630
rect 2100 5620 2150 5630
rect 2250 5620 2350 5630
rect 2400 5620 2450 5630
rect 2800 5620 2900 5630
rect 3150 5620 3200 5630
rect 3800 5620 3950 5630
rect 5050 5620 5100 5630
rect 5500 5620 5600 5630
rect 5800 5620 5950 5630
rect 6300 5620 6450 5630
rect 6950 5620 7000 5630
rect 7450 5620 7550 5630
rect 7850 5620 7900 5630
rect 8050 5620 8300 5630
rect 8400 5620 8500 5630
rect 500 5610 750 5620
rect 1950 5610 2050 5620
rect 2100 5610 2150 5620
rect 2250 5610 2350 5620
rect 2400 5610 2450 5620
rect 2800 5610 2900 5620
rect 3150 5610 3200 5620
rect 3800 5610 3950 5620
rect 5050 5610 5100 5620
rect 5500 5610 5600 5620
rect 5800 5610 5950 5620
rect 6300 5610 6450 5620
rect 6950 5610 7000 5620
rect 7450 5610 7550 5620
rect 7850 5610 7900 5620
rect 8050 5610 8300 5620
rect 8400 5610 8500 5620
rect 500 5600 750 5610
rect 1950 5600 2050 5610
rect 2100 5600 2150 5610
rect 2250 5600 2350 5610
rect 2400 5600 2450 5610
rect 2800 5600 2900 5610
rect 3150 5600 3200 5610
rect 3800 5600 3950 5610
rect 5050 5600 5100 5610
rect 5500 5600 5600 5610
rect 5800 5600 5950 5610
rect 6300 5600 6450 5610
rect 6950 5600 7000 5610
rect 7450 5600 7550 5610
rect 7850 5600 7900 5610
rect 8050 5600 8300 5610
rect 8400 5600 8500 5610
rect 500 5590 650 5600
rect 2000 5590 2150 5600
rect 2250 5590 2400 5600
rect 2700 5590 2850 5600
rect 2950 5590 3000 5600
rect 3150 5590 3200 5600
rect 5250 5590 5300 5600
rect 5450 5590 5500 5600
rect 5950 5590 6200 5600
rect 6550 5590 6650 5600
rect 6850 5590 6900 5600
rect 6950 5590 7000 5600
rect 7350 5590 7400 5600
rect 7700 5590 7750 5600
rect 7800 5590 7950 5600
rect 8050 5590 8250 5600
rect 8950 5590 9050 5600
rect 500 5580 650 5590
rect 2000 5580 2150 5590
rect 2250 5580 2400 5590
rect 2700 5580 2850 5590
rect 2950 5580 3000 5590
rect 3150 5580 3200 5590
rect 5250 5580 5300 5590
rect 5450 5580 5500 5590
rect 5950 5580 6200 5590
rect 6550 5580 6650 5590
rect 6850 5580 6900 5590
rect 6950 5580 7000 5590
rect 7350 5580 7400 5590
rect 7700 5580 7750 5590
rect 7800 5580 7950 5590
rect 8050 5580 8250 5590
rect 8950 5580 9050 5590
rect 500 5570 650 5580
rect 2000 5570 2150 5580
rect 2250 5570 2400 5580
rect 2700 5570 2850 5580
rect 2950 5570 3000 5580
rect 3150 5570 3200 5580
rect 5250 5570 5300 5580
rect 5450 5570 5500 5580
rect 5950 5570 6200 5580
rect 6550 5570 6650 5580
rect 6850 5570 6900 5580
rect 6950 5570 7000 5580
rect 7350 5570 7400 5580
rect 7700 5570 7750 5580
rect 7800 5570 7950 5580
rect 8050 5570 8250 5580
rect 8950 5570 9050 5580
rect 500 5560 650 5570
rect 2000 5560 2150 5570
rect 2250 5560 2400 5570
rect 2700 5560 2850 5570
rect 2950 5560 3000 5570
rect 3150 5560 3200 5570
rect 5250 5560 5300 5570
rect 5450 5560 5500 5570
rect 5950 5560 6200 5570
rect 6550 5560 6650 5570
rect 6850 5560 6900 5570
rect 6950 5560 7000 5570
rect 7350 5560 7400 5570
rect 7700 5560 7750 5570
rect 7800 5560 7950 5570
rect 8050 5560 8250 5570
rect 8950 5560 9050 5570
rect 500 5550 650 5560
rect 2000 5550 2150 5560
rect 2250 5550 2400 5560
rect 2700 5550 2850 5560
rect 2950 5550 3000 5560
rect 3150 5550 3200 5560
rect 5250 5550 5300 5560
rect 5450 5550 5500 5560
rect 5950 5550 6200 5560
rect 6550 5550 6650 5560
rect 6850 5550 6900 5560
rect 6950 5550 7000 5560
rect 7350 5550 7400 5560
rect 7700 5550 7750 5560
rect 7800 5550 7950 5560
rect 8050 5550 8250 5560
rect 8950 5550 9050 5560
rect 450 5540 500 5550
rect 2000 5540 2150 5550
rect 2250 5540 2350 5550
rect 2700 5540 2800 5550
rect 3000 5540 3050 5550
rect 3150 5540 3200 5550
rect 3650 5540 3700 5550
rect 3750 5540 3800 5550
rect 5250 5540 5300 5550
rect 5400 5540 5500 5550
rect 6000 5540 6150 5550
rect 6600 5540 6700 5550
rect 6850 5540 6900 5550
rect 6950 5540 7000 5550
rect 7250 5540 7350 5550
rect 7550 5540 7700 5550
rect 7800 5540 7950 5550
rect 8050 5540 8100 5550
rect 8850 5540 8900 5550
rect 8950 5540 9000 5550
rect 450 5530 500 5540
rect 2000 5530 2150 5540
rect 2250 5530 2350 5540
rect 2700 5530 2800 5540
rect 3000 5530 3050 5540
rect 3150 5530 3200 5540
rect 3650 5530 3700 5540
rect 3750 5530 3800 5540
rect 5250 5530 5300 5540
rect 5400 5530 5500 5540
rect 6000 5530 6150 5540
rect 6600 5530 6700 5540
rect 6850 5530 6900 5540
rect 6950 5530 7000 5540
rect 7250 5530 7350 5540
rect 7550 5530 7700 5540
rect 7800 5530 7950 5540
rect 8050 5530 8100 5540
rect 8850 5530 8900 5540
rect 8950 5530 9000 5540
rect 450 5520 500 5530
rect 2000 5520 2150 5530
rect 2250 5520 2350 5530
rect 2700 5520 2800 5530
rect 3000 5520 3050 5530
rect 3150 5520 3200 5530
rect 3650 5520 3700 5530
rect 3750 5520 3800 5530
rect 5250 5520 5300 5530
rect 5400 5520 5500 5530
rect 6000 5520 6150 5530
rect 6600 5520 6700 5530
rect 6850 5520 6900 5530
rect 6950 5520 7000 5530
rect 7250 5520 7350 5530
rect 7550 5520 7700 5530
rect 7800 5520 7950 5530
rect 8050 5520 8100 5530
rect 8850 5520 8900 5530
rect 8950 5520 9000 5530
rect 450 5510 500 5520
rect 2000 5510 2150 5520
rect 2250 5510 2350 5520
rect 2700 5510 2800 5520
rect 3000 5510 3050 5520
rect 3150 5510 3200 5520
rect 3650 5510 3700 5520
rect 3750 5510 3800 5520
rect 5250 5510 5300 5520
rect 5400 5510 5500 5520
rect 6000 5510 6150 5520
rect 6600 5510 6700 5520
rect 6850 5510 6900 5520
rect 6950 5510 7000 5520
rect 7250 5510 7350 5520
rect 7550 5510 7700 5520
rect 7800 5510 7950 5520
rect 8050 5510 8100 5520
rect 8850 5510 8900 5520
rect 8950 5510 9000 5520
rect 450 5500 500 5510
rect 2000 5500 2150 5510
rect 2250 5500 2350 5510
rect 2700 5500 2800 5510
rect 3000 5500 3050 5510
rect 3150 5500 3200 5510
rect 3650 5500 3700 5510
rect 3750 5500 3800 5510
rect 5250 5500 5300 5510
rect 5400 5500 5500 5510
rect 6000 5500 6150 5510
rect 6600 5500 6700 5510
rect 6850 5500 6900 5510
rect 6950 5500 7000 5510
rect 7250 5500 7350 5510
rect 7550 5500 7700 5510
rect 7800 5500 7950 5510
rect 8050 5500 8100 5510
rect 8850 5500 8900 5510
rect 8950 5500 9000 5510
rect 400 5490 450 5500
rect 2000 5490 2150 5500
rect 2250 5490 2350 5500
rect 3050 5490 3150 5500
rect 3650 5490 3700 5500
rect 5400 5490 5450 5500
rect 5950 5490 6000 5500
rect 6100 5490 6150 5500
rect 6600 5490 6750 5500
rect 6950 5490 7000 5500
rect 7200 5490 7350 5500
rect 7500 5490 7750 5500
rect 7800 5490 7950 5500
rect 8700 5490 9000 5500
rect 9050 5490 9100 5500
rect 400 5480 450 5490
rect 2000 5480 2150 5490
rect 2250 5480 2350 5490
rect 3050 5480 3150 5490
rect 3650 5480 3700 5490
rect 5400 5480 5450 5490
rect 5950 5480 6000 5490
rect 6100 5480 6150 5490
rect 6600 5480 6750 5490
rect 6950 5480 7000 5490
rect 7200 5480 7350 5490
rect 7500 5480 7750 5490
rect 7800 5480 7950 5490
rect 8700 5480 9000 5490
rect 9050 5480 9100 5490
rect 400 5470 450 5480
rect 2000 5470 2150 5480
rect 2250 5470 2350 5480
rect 3050 5470 3150 5480
rect 3650 5470 3700 5480
rect 5400 5470 5450 5480
rect 5950 5470 6000 5480
rect 6100 5470 6150 5480
rect 6600 5470 6750 5480
rect 6950 5470 7000 5480
rect 7200 5470 7350 5480
rect 7500 5470 7750 5480
rect 7800 5470 7950 5480
rect 8700 5470 9000 5480
rect 9050 5470 9100 5480
rect 400 5460 450 5470
rect 2000 5460 2150 5470
rect 2250 5460 2350 5470
rect 3050 5460 3150 5470
rect 3650 5460 3700 5470
rect 5400 5460 5450 5470
rect 5950 5460 6000 5470
rect 6100 5460 6150 5470
rect 6600 5460 6750 5470
rect 6950 5460 7000 5470
rect 7200 5460 7350 5470
rect 7500 5460 7750 5470
rect 7800 5460 7950 5470
rect 8700 5460 9000 5470
rect 9050 5460 9100 5470
rect 400 5450 450 5460
rect 2000 5450 2150 5460
rect 2250 5450 2350 5460
rect 3050 5450 3150 5460
rect 3650 5450 3700 5460
rect 5400 5450 5450 5460
rect 5950 5450 6000 5460
rect 6100 5450 6150 5460
rect 6600 5450 6750 5460
rect 6950 5450 7000 5460
rect 7200 5450 7350 5460
rect 7500 5450 7750 5460
rect 7800 5450 7950 5460
rect 8700 5450 9000 5460
rect 9050 5450 9100 5460
rect 400 5440 450 5450
rect 500 5440 550 5450
rect 2050 5440 2150 5450
rect 2250 5440 2350 5450
rect 5050 5440 5100 5450
rect 5400 5440 5450 5450
rect 5950 5440 6000 5450
rect 6100 5440 6150 5450
rect 6650 5440 6750 5450
rect 6900 5440 6950 5450
rect 7200 5440 7250 5450
rect 7500 5440 7550 5450
rect 7600 5440 7750 5450
rect 8400 5440 8450 5450
rect 8500 5440 8950 5450
rect 9000 5440 9100 5450
rect 400 5430 450 5440
rect 500 5430 550 5440
rect 2050 5430 2150 5440
rect 2250 5430 2350 5440
rect 5050 5430 5100 5440
rect 5400 5430 5450 5440
rect 5950 5430 6000 5440
rect 6100 5430 6150 5440
rect 6650 5430 6750 5440
rect 6900 5430 6950 5440
rect 7200 5430 7250 5440
rect 7500 5430 7550 5440
rect 7600 5430 7750 5440
rect 8400 5430 8450 5440
rect 8500 5430 8950 5440
rect 9000 5430 9100 5440
rect 400 5420 450 5430
rect 500 5420 550 5430
rect 2050 5420 2150 5430
rect 2250 5420 2350 5430
rect 5050 5420 5100 5430
rect 5400 5420 5450 5430
rect 5950 5420 6000 5430
rect 6100 5420 6150 5430
rect 6650 5420 6750 5430
rect 6900 5420 6950 5430
rect 7200 5420 7250 5430
rect 7500 5420 7550 5430
rect 7600 5420 7750 5430
rect 8400 5420 8450 5430
rect 8500 5420 8950 5430
rect 9000 5420 9100 5430
rect 400 5410 450 5420
rect 500 5410 550 5420
rect 2050 5410 2150 5420
rect 2250 5410 2350 5420
rect 5050 5410 5100 5420
rect 5400 5410 5450 5420
rect 5950 5410 6000 5420
rect 6100 5410 6150 5420
rect 6650 5410 6750 5420
rect 6900 5410 6950 5420
rect 7200 5410 7250 5420
rect 7500 5410 7550 5420
rect 7600 5410 7750 5420
rect 8400 5410 8450 5420
rect 8500 5410 8950 5420
rect 9000 5410 9100 5420
rect 400 5400 450 5410
rect 500 5400 550 5410
rect 2050 5400 2150 5410
rect 2250 5400 2350 5410
rect 5050 5400 5100 5410
rect 5400 5400 5450 5410
rect 5950 5400 6000 5410
rect 6100 5400 6150 5410
rect 6650 5400 6750 5410
rect 6900 5400 6950 5410
rect 7200 5400 7250 5410
rect 7500 5400 7550 5410
rect 7600 5400 7750 5410
rect 8400 5400 8450 5410
rect 8500 5400 8950 5410
rect 9000 5400 9100 5410
rect 300 5390 350 5400
rect 500 5390 550 5400
rect 2250 5390 2350 5400
rect 3550 5390 3600 5400
rect 5050 5390 5100 5400
rect 5350 5390 5400 5400
rect 5950 5390 6000 5400
rect 6700 5390 6750 5400
rect 6900 5390 6950 5400
rect 7200 5390 7300 5400
rect 7550 5390 7600 5400
rect 8350 5390 8500 5400
rect 8550 5390 8850 5400
rect 9500 5390 9550 5400
rect 300 5380 350 5390
rect 500 5380 550 5390
rect 2250 5380 2350 5390
rect 3550 5380 3600 5390
rect 5050 5380 5100 5390
rect 5350 5380 5400 5390
rect 5950 5380 6000 5390
rect 6700 5380 6750 5390
rect 6900 5380 6950 5390
rect 7200 5380 7300 5390
rect 7550 5380 7600 5390
rect 8350 5380 8500 5390
rect 8550 5380 8850 5390
rect 9500 5380 9550 5390
rect 300 5370 350 5380
rect 500 5370 550 5380
rect 2250 5370 2350 5380
rect 3550 5370 3600 5380
rect 5050 5370 5100 5380
rect 5350 5370 5400 5380
rect 5950 5370 6000 5380
rect 6700 5370 6750 5380
rect 6900 5370 6950 5380
rect 7200 5370 7300 5380
rect 7550 5370 7600 5380
rect 8350 5370 8500 5380
rect 8550 5370 8850 5380
rect 9500 5370 9550 5380
rect 300 5360 350 5370
rect 500 5360 550 5370
rect 2250 5360 2350 5370
rect 3550 5360 3600 5370
rect 5050 5360 5100 5370
rect 5350 5360 5400 5370
rect 5950 5360 6000 5370
rect 6700 5360 6750 5370
rect 6900 5360 6950 5370
rect 7200 5360 7300 5370
rect 7550 5360 7600 5370
rect 8350 5360 8500 5370
rect 8550 5360 8850 5370
rect 9500 5360 9550 5370
rect 300 5350 350 5360
rect 500 5350 550 5360
rect 2250 5350 2350 5360
rect 3550 5350 3600 5360
rect 5050 5350 5100 5360
rect 5350 5350 5400 5360
rect 5950 5350 6000 5360
rect 6700 5350 6750 5360
rect 6900 5350 6950 5360
rect 7200 5350 7300 5360
rect 7550 5350 7600 5360
rect 8350 5350 8500 5360
rect 8550 5350 8850 5360
rect 9500 5350 9550 5360
rect 200 5340 250 5350
rect 450 5340 550 5350
rect 2250 5340 2350 5350
rect 3550 5340 3600 5350
rect 5050 5340 5100 5350
rect 5400 5340 5650 5350
rect 5900 5340 5950 5350
rect 6750 5340 6800 5350
rect 7250 5340 7300 5350
rect 8100 5340 8150 5350
rect 8250 5340 8300 5350
rect 8350 5340 8500 5350
rect 8550 5340 8700 5350
rect 9250 5340 9300 5350
rect 9550 5340 9600 5350
rect 200 5330 250 5340
rect 450 5330 550 5340
rect 2250 5330 2350 5340
rect 3550 5330 3600 5340
rect 5050 5330 5100 5340
rect 5400 5330 5650 5340
rect 5900 5330 5950 5340
rect 6750 5330 6800 5340
rect 7250 5330 7300 5340
rect 8100 5330 8150 5340
rect 8250 5330 8300 5340
rect 8350 5330 8500 5340
rect 8550 5330 8700 5340
rect 9250 5330 9300 5340
rect 9550 5330 9600 5340
rect 200 5320 250 5330
rect 450 5320 550 5330
rect 2250 5320 2350 5330
rect 3550 5320 3600 5330
rect 5050 5320 5100 5330
rect 5400 5320 5650 5330
rect 5900 5320 5950 5330
rect 6750 5320 6800 5330
rect 7250 5320 7300 5330
rect 8100 5320 8150 5330
rect 8250 5320 8300 5330
rect 8350 5320 8500 5330
rect 8550 5320 8700 5330
rect 9250 5320 9300 5330
rect 9550 5320 9600 5330
rect 200 5310 250 5320
rect 450 5310 550 5320
rect 2250 5310 2350 5320
rect 3550 5310 3600 5320
rect 5050 5310 5100 5320
rect 5400 5310 5650 5320
rect 5900 5310 5950 5320
rect 6750 5310 6800 5320
rect 7250 5310 7300 5320
rect 8100 5310 8150 5320
rect 8250 5310 8300 5320
rect 8350 5310 8500 5320
rect 8550 5310 8700 5320
rect 9250 5310 9300 5320
rect 9550 5310 9600 5320
rect 200 5300 250 5310
rect 450 5300 550 5310
rect 2250 5300 2350 5310
rect 3550 5300 3600 5310
rect 5050 5300 5100 5310
rect 5400 5300 5650 5310
rect 5900 5300 5950 5310
rect 6750 5300 6800 5310
rect 7250 5300 7300 5310
rect 8100 5300 8150 5310
rect 8250 5300 8300 5310
rect 8350 5300 8500 5310
rect 8550 5300 8700 5310
rect 9250 5300 9300 5310
rect 9550 5300 9600 5310
rect 150 5290 300 5300
rect 350 5290 550 5300
rect 2250 5290 2350 5300
rect 5050 5290 5100 5300
rect 5200 5290 5250 5300
rect 5550 5290 5650 5300
rect 5850 5290 5900 5300
rect 6150 5290 6200 5300
rect 6500 5290 6800 5300
rect 8000 5290 8050 5300
rect 8150 5290 8350 5300
rect 8400 5290 8500 5300
rect 150 5280 300 5290
rect 350 5280 550 5290
rect 2250 5280 2350 5290
rect 5050 5280 5100 5290
rect 5200 5280 5250 5290
rect 5550 5280 5650 5290
rect 5850 5280 5900 5290
rect 6150 5280 6200 5290
rect 6500 5280 6800 5290
rect 8000 5280 8050 5290
rect 8150 5280 8350 5290
rect 8400 5280 8500 5290
rect 150 5270 300 5280
rect 350 5270 550 5280
rect 2250 5270 2350 5280
rect 5050 5270 5100 5280
rect 5200 5270 5250 5280
rect 5550 5270 5650 5280
rect 5850 5270 5900 5280
rect 6150 5270 6200 5280
rect 6500 5270 6800 5280
rect 8000 5270 8050 5280
rect 8150 5270 8350 5280
rect 8400 5270 8500 5280
rect 150 5260 300 5270
rect 350 5260 550 5270
rect 2250 5260 2350 5270
rect 5050 5260 5100 5270
rect 5200 5260 5250 5270
rect 5550 5260 5650 5270
rect 5850 5260 5900 5270
rect 6150 5260 6200 5270
rect 6500 5260 6800 5270
rect 8000 5260 8050 5270
rect 8150 5260 8350 5270
rect 8400 5260 8500 5270
rect 150 5250 300 5260
rect 350 5250 550 5260
rect 2250 5250 2350 5260
rect 5050 5250 5100 5260
rect 5200 5250 5250 5260
rect 5550 5250 5650 5260
rect 5850 5250 5900 5260
rect 6150 5250 6200 5260
rect 6500 5250 6800 5260
rect 8000 5250 8050 5260
rect 8150 5250 8350 5260
rect 8400 5250 8500 5260
rect 100 5240 600 5250
rect 2250 5240 2350 5250
rect 2500 5240 2650 5250
rect 3500 5240 3550 5250
rect 5200 5240 5250 5250
rect 5600 5240 5800 5250
rect 6200 5240 6350 5250
rect 6550 5240 6600 5250
rect 7200 5240 7300 5250
rect 8000 5240 8050 5250
rect 8150 5240 8350 5250
rect 8950 5240 9000 5250
rect 9050 5240 9200 5250
rect 9750 5240 9800 5250
rect 9850 5240 9900 5250
rect 9950 5240 9990 5250
rect 100 5230 600 5240
rect 2250 5230 2350 5240
rect 2500 5230 2650 5240
rect 3500 5230 3550 5240
rect 5200 5230 5250 5240
rect 5600 5230 5800 5240
rect 6200 5230 6350 5240
rect 6550 5230 6600 5240
rect 7200 5230 7300 5240
rect 8000 5230 8050 5240
rect 8150 5230 8350 5240
rect 8950 5230 9000 5240
rect 9050 5230 9200 5240
rect 9750 5230 9800 5240
rect 9850 5230 9900 5240
rect 9950 5230 9990 5240
rect 100 5220 600 5230
rect 2250 5220 2350 5230
rect 2500 5220 2650 5230
rect 3500 5220 3550 5230
rect 5200 5220 5250 5230
rect 5600 5220 5800 5230
rect 6200 5220 6350 5230
rect 6550 5220 6600 5230
rect 7200 5220 7300 5230
rect 8000 5220 8050 5230
rect 8150 5220 8350 5230
rect 8950 5220 9000 5230
rect 9050 5220 9200 5230
rect 9750 5220 9800 5230
rect 9850 5220 9900 5230
rect 9950 5220 9990 5230
rect 100 5210 600 5220
rect 2250 5210 2350 5220
rect 2500 5210 2650 5220
rect 3500 5210 3550 5220
rect 5200 5210 5250 5220
rect 5600 5210 5800 5220
rect 6200 5210 6350 5220
rect 6550 5210 6600 5220
rect 7200 5210 7300 5220
rect 8000 5210 8050 5220
rect 8150 5210 8350 5220
rect 8950 5210 9000 5220
rect 9050 5210 9200 5220
rect 9750 5210 9800 5220
rect 9850 5210 9900 5220
rect 9950 5210 9990 5220
rect 100 5200 600 5210
rect 2250 5200 2350 5210
rect 2500 5200 2650 5210
rect 3500 5200 3550 5210
rect 5200 5200 5250 5210
rect 5600 5200 5800 5210
rect 6200 5200 6350 5210
rect 6550 5200 6600 5210
rect 7200 5200 7300 5210
rect 8000 5200 8050 5210
rect 8150 5200 8350 5210
rect 8950 5200 9000 5210
rect 9050 5200 9200 5210
rect 9750 5200 9800 5210
rect 9850 5200 9900 5210
rect 9950 5200 9990 5210
rect 50 5190 600 5200
rect 2250 5190 2350 5200
rect 2500 5190 2550 5200
rect 2650 5190 2700 5200
rect 5050 5190 5100 5200
rect 5200 5190 5250 5200
rect 7250 5190 7300 5200
rect 8050 5190 8200 5200
rect 8650 5190 8700 5200
rect 8750 5190 8800 5200
rect 8950 5190 9000 5200
rect 9700 5190 9750 5200
rect 9950 5190 9990 5200
rect 50 5180 600 5190
rect 2250 5180 2350 5190
rect 2500 5180 2550 5190
rect 2650 5180 2700 5190
rect 5050 5180 5100 5190
rect 5200 5180 5250 5190
rect 7250 5180 7300 5190
rect 8050 5180 8200 5190
rect 8650 5180 8700 5190
rect 8750 5180 8800 5190
rect 8950 5180 9000 5190
rect 9700 5180 9750 5190
rect 9950 5180 9990 5190
rect 50 5170 600 5180
rect 2250 5170 2350 5180
rect 2500 5170 2550 5180
rect 2650 5170 2700 5180
rect 5050 5170 5100 5180
rect 5200 5170 5250 5180
rect 7250 5170 7300 5180
rect 8050 5170 8200 5180
rect 8650 5170 8700 5180
rect 8750 5170 8800 5180
rect 8950 5170 9000 5180
rect 9700 5170 9750 5180
rect 9950 5170 9990 5180
rect 50 5160 600 5170
rect 2250 5160 2350 5170
rect 2500 5160 2550 5170
rect 2650 5160 2700 5170
rect 5050 5160 5100 5170
rect 5200 5160 5250 5170
rect 7250 5160 7300 5170
rect 8050 5160 8200 5170
rect 8650 5160 8700 5170
rect 8750 5160 8800 5170
rect 8950 5160 9000 5170
rect 9700 5160 9750 5170
rect 9950 5160 9990 5170
rect 50 5150 600 5160
rect 2250 5150 2350 5160
rect 2500 5150 2550 5160
rect 2650 5150 2700 5160
rect 5050 5150 5100 5160
rect 5200 5150 5250 5160
rect 7250 5150 7300 5160
rect 8050 5150 8200 5160
rect 8650 5150 8700 5160
rect 8750 5150 8800 5160
rect 8950 5150 9000 5160
rect 9700 5150 9750 5160
rect 9950 5150 9990 5160
rect 0 5140 500 5150
rect 2300 5140 2400 5150
rect 2500 5140 2550 5150
rect 2600 5140 2700 5150
rect 5100 5140 5150 5150
rect 5200 5140 5250 5150
rect 8650 5140 8700 5150
rect 8850 5140 8900 5150
rect 9400 5140 9450 5150
rect 9800 5140 9850 5150
rect 0 5130 500 5140
rect 2300 5130 2400 5140
rect 2500 5130 2550 5140
rect 2600 5130 2700 5140
rect 5100 5130 5150 5140
rect 5200 5130 5250 5140
rect 8650 5130 8700 5140
rect 8850 5130 8900 5140
rect 9400 5130 9450 5140
rect 9800 5130 9850 5140
rect 0 5120 500 5130
rect 2300 5120 2400 5130
rect 2500 5120 2550 5130
rect 2600 5120 2700 5130
rect 5100 5120 5150 5130
rect 5200 5120 5250 5130
rect 8650 5120 8700 5130
rect 8850 5120 8900 5130
rect 9400 5120 9450 5130
rect 9800 5120 9850 5130
rect 0 5110 500 5120
rect 2300 5110 2400 5120
rect 2500 5110 2550 5120
rect 2600 5110 2700 5120
rect 5100 5110 5150 5120
rect 5200 5110 5250 5120
rect 8650 5110 8700 5120
rect 8850 5110 8900 5120
rect 9400 5110 9450 5120
rect 9800 5110 9850 5120
rect 0 5100 500 5110
rect 2300 5100 2400 5110
rect 2500 5100 2550 5110
rect 2600 5100 2700 5110
rect 5100 5100 5150 5110
rect 5200 5100 5250 5110
rect 8650 5100 8700 5110
rect 8850 5100 8900 5110
rect 9400 5100 9450 5110
rect 9800 5100 9850 5110
rect 0 5090 350 5100
rect 2300 5090 2400 5100
rect 2500 5090 2650 5100
rect 3400 5090 3450 5100
rect 5200 5090 5250 5100
rect 8300 5090 8400 5100
rect 8450 5090 8500 5100
rect 9150 5090 9200 5100
rect 9250 5090 9300 5100
rect 9400 5090 9450 5100
rect 9600 5090 9650 5100
rect 0 5080 350 5090
rect 2300 5080 2400 5090
rect 2500 5080 2650 5090
rect 3400 5080 3450 5090
rect 5200 5080 5250 5090
rect 8300 5080 8400 5090
rect 8450 5080 8500 5090
rect 9150 5080 9200 5090
rect 9250 5080 9300 5090
rect 9400 5080 9450 5090
rect 9600 5080 9650 5090
rect 0 5070 350 5080
rect 2300 5070 2400 5080
rect 2500 5070 2650 5080
rect 3400 5070 3450 5080
rect 5200 5070 5250 5080
rect 8300 5070 8400 5080
rect 8450 5070 8500 5080
rect 9150 5070 9200 5080
rect 9250 5070 9300 5080
rect 9400 5070 9450 5080
rect 9600 5070 9650 5080
rect 0 5060 350 5070
rect 2300 5060 2400 5070
rect 2500 5060 2650 5070
rect 3400 5060 3450 5070
rect 5200 5060 5250 5070
rect 8300 5060 8400 5070
rect 8450 5060 8500 5070
rect 9150 5060 9200 5070
rect 9250 5060 9300 5070
rect 9400 5060 9450 5070
rect 9600 5060 9650 5070
rect 0 5050 350 5060
rect 2300 5050 2400 5060
rect 2500 5050 2650 5060
rect 3400 5050 3450 5060
rect 5200 5050 5250 5060
rect 8300 5050 8400 5060
rect 8450 5050 8500 5060
rect 9150 5050 9200 5060
rect 9250 5050 9300 5060
rect 9400 5050 9450 5060
rect 9600 5050 9650 5060
rect 0 5040 150 5050
rect 200 5040 350 5050
rect 2300 5040 2400 5050
rect 3400 5040 3450 5050
rect 5200 5040 5250 5050
rect 5650 5040 5800 5050
rect 6300 5040 6400 5050
rect 8150 5040 8400 5050
rect 8450 5040 8500 5050
rect 9150 5040 9200 5050
rect 9400 5040 9450 5050
rect 0 5030 150 5040
rect 200 5030 350 5040
rect 2300 5030 2400 5040
rect 3400 5030 3450 5040
rect 5200 5030 5250 5040
rect 5650 5030 5800 5040
rect 6300 5030 6400 5040
rect 8150 5030 8400 5040
rect 8450 5030 8500 5040
rect 9150 5030 9200 5040
rect 9400 5030 9450 5040
rect 0 5020 150 5030
rect 200 5020 350 5030
rect 2300 5020 2400 5030
rect 3400 5020 3450 5030
rect 5200 5020 5250 5030
rect 5650 5020 5800 5030
rect 6300 5020 6400 5030
rect 8150 5020 8400 5030
rect 8450 5020 8500 5030
rect 9150 5020 9200 5030
rect 9400 5020 9450 5030
rect 0 5010 150 5020
rect 200 5010 350 5020
rect 2300 5010 2400 5020
rect 3400 5010 3450 5020
rect 5200 5010 5250 5020
rect 5650 5010 5800 5020
rect 6300 5010 6400 5020
rect 8150 5010 8400 5020
rect 8450 5010 8500 5020
rect 9150 5010 9200 5020
rect 9400 5010 9450 5020
rect 0 5000 150 5010
rect 200 5000 350 5010
rect 2300 5000 2400 5010
rect 3400 5000 3450 5010
rect 5200 5000 5250 5010
rect 5650 5000 5800 5010
rect 6300 5000 6400 5010
rect 8150 5000 8400 5010
rect 8450 5000 8500 5010
rect 9150 5000 9200 5010
rect 9400 5000 9450 5010
rect 0 4990 150 5000
rect 2350 4990 2450 5000
rect 4000 4990 4100 5000
rect 4350 4990 4400 5000
rect 4500 4990 4600 5000
rect 5150 4990 5250 5000
rect 5500 4990 5650 5000
rect 5750 4990 5900 5000
rect 6050 4990 6200 5000
rect 6300 4990 6350 5000
rect 6400 4990 6500 5000
rect 8000 4990 8200 5000
rect 8250 4990 8400 5000
rect 8750 4990 8800 5000
rect 8900 4990 9000 5000
rect 9150 4990 9200 5000
rect 0 4980 150 4990
rect 2350 4980 2450 4990
rect 4000 4980 4100 4990
rect 4350 4980 4400 4990
rect 4500 4980 4600 4990
rect 5150 4980 5250 4990
rect 5500 4980 5650 4990
rect 5750 4980 5900 4990
rect 6050 4980 6200 4990
rect 6300 4980 6350 4990
rect 6400 4980 6500 4990
rect 8000 4980 8200 4990
rect 8250 4980 8400 4990
rect 8750 4980 8800 4990
rect 8900 4980 9000 4990
rect 9150 4980 9200 4990
rect 0 4970 150 4980
rect 2350 4970 2450 4980
rect 4000 4970 4100 4980
rect 4350 4970 4400 4980
rect 4500 4970 4600 4980
rect 5150 4970 5250 4980
rect 5500 4970 5650 4980
rect 5750 4970 5900 4980
rect 6050 4970 6200 4980
rect 6300 4970 6350 4980
rect 6400 4970 6500 4980
rect 8000 4970 8200 4980
rect 8250 4970 8400 4980
rect 8750 4970 8800 4980
rect 8900 4970 9000 4980
rect 9150 4970 9200 4980
rect 0 4960 150 4970
rect 2350 4960 2450 4970
rect 4000 4960 4100 4970
rect 4350 4960 4400 4970
rect 4500 4960 4600 4970
rect 5150 4960 5250 4970
rect 5500 4960 5650 4970
rect 5750 4960 5900 4970
rect 6050 4960 6200 4970
rect 6300 4960 6350 4970
rect 6400 4960 6500 4970
rect 8000 4960 8200 4970
rect 8250 4960 8400 4970
rect 8750 4960 8800 4970
rect 8900 4960 9000 4970
rect 9150 4960 9200 4970
rect 0 4950 150 4960
rect 2350 4950 2450 4960
rect 4000 4950 4100 4960
rect 4350 4950 4400 4960
rect 4500 4950 4600 4960
rect 5150 4950 5250 4960
rect 5500 4950 5650 4960
rect 5750 4950 5900 4960
rect 6050 4950 6200 4960
rect 6300 4950 6350 4960
rect 6400 4950 6500 4960
rect 8000 4950 8200 4960
rect 8250 4950 8400 4960
rect 8750 4950 8800 4960
rect 8900 4950 9000 4960
rect 9150 4950 9200 4960
rect 0 4940 50 4950
rect 2400 4940 2450 4950
rect 3350 4940 3400 4950
rect 3900 4940 4000 4950
rect 4100 4940 4150 4950
rect 4500 4940 4800 4950
rect 5200 4940 5250 4950
rect 5450 4940 5550 4950
rect 6000 4940 6050 4950
rect 6500 4940 6700 4950
rect 7300 4940 7350 4950
rect 7850 4940 7950 4950
rect 8000 4940 8050 4950
rect 8100 4940 8150 4950
rect 8200 4940 8250 4950
rect 8600 4940 8650 4950
rect 8750 4940 8850 4950
rect 8900 4940 9000 4950
rect 9250 4940 9300 4950
rect 9550 4940 9650 4950
rect 0 4930 50 4940
rect 2400 4930 2450 4940
rect 3350 4930 3400 4940
rect 3900 4930 4000 4940
rect 4100 4930 4150 4940
rect 4500 4930 4800 4940
rect 5200 4930 5250 4940
rect 5450 4930 5550 4940
rect 6000 4930 6050 4940
rect 6500 4930 6700 4940
rect 7300 4930 7350 4940
rect 7850 4930 7950 4940
rect 8000 4930 8050 4940
rect 8100 4930 8150 4940
rect 8200 4930 8250 4940
rect 8600 4930 8650 4940
rect 8750 4930 8850 4940
rect 8900 4930 9000 4940
rect 9250 4930 9300 4940
rect 9550 4930 9650 4940
rect 0 4920 50 4930
rect 2400 4920 2450 4930
rect 3350 4920 3400 4930
rect 3900 4920 4000 4930
rect 4100 4920 4150 4930
rect 4500 4920 4800 4930
rect 5200 4920 5250 4930
rect 5450 4920 5550 4930
rect 6000 4920 6050 4930
rect 6500 4920 6700 4930
rect 7300 4920 7350 4930
rect 7850 4920 7950 4930
rect 8000 4920 8050 4930
rect 8100 4920 8150 4930
rect 8200 4920 8250 4930
rect 8600 4920 8650 4930
rect 8750 4920 8850 4930
rect 8900 4920 9000 4930
rect 9250 4920 9300 4930
rect 9550 4920 9650 4930
rect 0 4910 50 4920
rect 2400 4910 2450 4920
rect 3350 4910 3400 4920
rect 3900 4910 4000 4920
rect 4100 4910 4150 4920
rect 4500 4910 4800 4920
rect 5200 4910 5250 4920
rect 5450 4910 5550 4920
rect 6000 4910 6050 4920
rect 6500 4910 6700 4920
rect 7300 4910 7350 4920
rect 7850 4910 7950 4920
rect 8000 4910 8050 4920
rect 8100 4910 8150 4920
rect 8200 4910 8250 4920
rect 8600 4910 8650 4920
rect 8750 4910 8850 4920
rect 8900 4910 9000 4920
rect 9250 4910 9300 4920
rect 9550 4910 9650 4920
rect 0 4900 50 4910
rect 2400 4900 2450 4910
rect 3350 4900 3400 4910
rect 3900 4900 4000 4910
rect 4100 4900 4150 4910
rect 4500 4900 4800 4910
rect 5200 4900 5250 4910
rect 5450 4900 5550 4910
rect 6000 4900 6050 4910
rect 6500 4900 6700 4910
rect 7300 4900 7350 4910
rect 7850 4900 7950 4910
rect 8000 4900 8050 4910
rect 8100 4900 8150 4910
rect 8200 4900 8250 4910
rect 8600 4900 8650 4910
rect 8750 4900 8850 4910
rect 8900 4900 9000 4910
rect 9250 4900 9300 4910
rect 9550 4900 9650 4910
rect 2400 4890 2500 4900
rect 3350 4890 3400 4900
rect 3650 4890 3850 4900
rect 4850 4890 4950 4900
rect 5150 4890 5250 4900
rect 5350 4890 5500 4900
rect 6550 4890 6700 4900
rect 7300 4890 7350 4900
rect 7700 4890 7950 4900
rect 8500 4890 8550 4900
rect 8600 4890 8700 4900
rect 8750 4890 8850 4900
rect 9300 4890 9350 4900
rect 9450 4890 9600 4900
rect 9650 4890 9700 4900
rect 2400 4880 2500 4890
rect 3350 4880 3400 4890
rect 3650 4880 3850 4890
rect 4850 4880 4950 4890
rect 5150 4880 5250 4890
rect 5350 4880 5500 4890
rect 6550 4880 6700 4890
rect 7300 4880 7350 4890
rect 7700 4880 7950 4890
rect 8500 4880 8550 4890
rect 8600 4880 8700 4890
rect 8750 4880 8850 4890
rect 9300 4880 9350 4890
rect 9450 4880 9600 4890
rect 9650 4880 9700 4890
rect 2400 4870 2500 4880
rect 3350 4870 3400 4880
rect 3650 4870 3850 4880
rect 4850 4870 4950 4880
rect 5150 4870 5250 4880
rect 5350 4870 5500 4880
rect 6550 4870 6700 4880
rect 7300 4870 7350 4880
rect 7700 4870 7950 4880
rect 8500 4870 8550 4880
rect 8600 4870 8700 4880
rect 8750 4870 8850 4880
rect 9300 4870 9350 4880
rect 9450 4870 9600 4880
rect 9650 4870 9700 4880
rect 2400 4860 2500 4870
rect 3350 4860 3400 4870
rect 3650 4860 3850 4870
rect 4850 4860 4950 4870
rect 5150 4860 5250 4870
rect 5350 4860 5500 4870
rect 6550 4860 6700 4870
rect 7300 4860 7350 4870
rect 7700 4860 7950 4870
rect 8500 4860 8550 4870
rect 8600 4860 8700 4870
rect 8750 4860 8850 4870
rect 9300 4860 9350 4870
rect 9450 4860 9600 4870
rect 9650 4860 9700 4870
rect 2400 4850 2500 4860
rect 3350 4850 3400 4860
rect 3650 4850 3850 4860
rect 4850 4850 4950 4860
rect 5150 4850 5250 4860
rect 5350 4850 5500 4860
rect 6550 4850 6700 4860
rect 7300 4850 7350 4860
rect 7700 4850 7950 4860
rect 8500 4850 8550 4860
rect 8600 4850 8700 4860
rect 8750 4850 8850 4860
rect 9300 4850 9350 4860
rect 9450 4850 9600 4860
rect 9650 4850 9700 4860
rect 2450 4840 2600 4850
rect 3600 4840 3650 4850
rect 5000 4840 5050 4850
rect 5150 4840 5250 4850
rect 5350 4840 5450 4850
rect 5750 4840 5850 4850
rect 6600 4840 6700 4850
rect 7300 4840 7350 4850
rect 7700 4840 7800 4850
rect 7850 4840 7900 4850
rect 8300 4840 8350 4850
rect 8500 4840 8550 4850
rect 8650 4840 8700 4850
rect 9050 4840 9100 4850
rect 9300 4840 9350 4850
rect 9400 4840 9450 4850
rect 9500 4840 9550 4850
rect 9650 4840 9700 4850
rect 2450 4830 2600 4840
rect 3600 4830 3650 4840
rect 5000 4830 5050 4840
rect 5150 4830 5250 4840
rect 5350 4830 5450 4840
rect 5750 4830 5850 4840
rect 6600 4830 6700 4840
rect 7300 4830 7350 4840
rect 7700 4830 7800 4840
rect 7850 4830 7900 4840
rect 8300 4830 8350 4840
rect 8500 4830 8550 4840
rect 8650 4830 8700 4840
rect 9050 4830 9100 4840
rect 9300 4830 9350 4840
rect 9400 4830 9450 4840
rect 9500 4830 9550 4840
rect 9650 4830 9700 4840
rect 2450 4820 2600 4830
rect 3600 4820 3650 4830
rect 5000 4820 5050 4830
rect 5150 4820 5250 4830
rect 5350 4820 5450 4830
rect 5750 4820 5850 4830
rect 6600 4820 6700 4830
rect 7300 4820 7350 4830
rect 7700 4820 7800 4830
rect 7850 4820 7900 4830
rect 8300 4820 8350 4830
rect 8500 4820 8550 4830
rect 8650 4820 8700 4830
rect 9050 4820 9100 4830
rect 9300 4820 9350 4830
rect 9400 4820 9450 4830
rect 9500 4820 9550 4830
rect 9650 4820 9700 4830
rect 2450 4810 2600 4820
rect 3600 4810 3650 4820
rect 5000 4810 5050 4820
rect 5150 4810 5250 4820
rect 5350 4810 5450 4820
rect 5750 4810 5850 4820
rect 6600 4810 6700 4820
rect 7300 4810 7350 4820
rect 7700 4810 7800 4820
rect 7850 4810 7900 4820
rect 8300 4810 8350 4820
rect 8500 4810 8550 4820
rect 8650 4810 8700 4820
rect 9050 4810 9100 4820
rect 9300 4810 9350 4820
rect 9400 4810 9450 4820
rect 9500 4810 9550 4820
rect 9650 4810 9700 4820
rect 2450 4800 2600 4810
rect 3600 4800 3650 4810
rect 5000 4800 5050 4810
rect 5150 4800 5250 4810
rect 5350 4800 5450 4810
rect 5750 4800 5850 4810
rect 6600 4800 6700 4810
rect 7300 4800 7350 4810
rect 7700 4800 7800 4810
rect 7850 4800 7900 4810
rect 8300 4800 8350 4810
rect 8500 4800 8550 4810
rect 8650 4800 8700 4810
rect 9050 4800 9100 4810
rect 9300 4800 9350 4810
rect 9400 4800 9450 4810
rect 9500 4800 9550 4810
rect 9650 4800 9700 4810
rect 2500 4790 2650 4800
rect 3350 4790 3400 4800
rect 3500 4790 3600 4800
rect 5050 4790 5100 4800
rect 5200 4790 5250 4800
rect 5350 4790 5400 4800
rect 5700 4790 5800 4800
rect 5850 4790 5950 4800
rect 6650 4790 6750 4800
rect 8000 4790 8250 4800
rect 8300 4790 8400 4800
rect 9000 4790 9050 4800
rect 9300 4790 9350 4800
rect 2500 4780 2650 4790
rect 3350 4780 3400 4790
rect 3500 4780 3600 4790
rect 5050 4780 5100 4790
rect 5200 4780 5250 4790
rect 5350 4780 5400 4790
rect 5700 4780 5800 4790
rect 5850 4780 5950 4790
rect 6650 4780 6750 4790
rect 8000 4780 8250 4790
rect 8300 4780 8400 4790
rect 9000 4780 9050 4790
rect 9300 4780 9350 4790
rect 2500 4770 2650 4780
rect 3350 4770 3400 4780
rect 3500 4770 3600 4780
rect 5050 4770 5100 4780
rect 5200 4770 5250 4780
rect 5350 4770 5400 4780
rect 5700 4770 5800 4780
rect 5850 4770 5950 4780
rect 6650 4770 6750 4780
rect 8000 4770 8250 4780
rect 8300 4770 8400 4780
rect 9000 4770 9050 4780
rect 9300 4770 9350 4780
rect 2500 4760 2650 4770
rect 3350 4760 3400 4770
rect 3500 4760 3600 4770
rect 5050 4760 5100 4770
rect 5200 4760 5250 4770
rect 5350 4760 5400 4770
rect 5700 4760 5800 4770
rect 5850 4760 5950 4770
rect 6650 4760 6750 4770
rect 8000 4760 8250 4770
rect 8300 4760 8400 4770
rect 9000 4760 9050 4770
rect 9300 4760 9350 4770
rect 2500 4750 2650 4760
rect 3350 4750 3400 4760
rect 3500 4750 3600 4760
rect 5050 4750 5100 4760
rect 5200 4750 5250 4760
rect 5350 4750 5400 4760
rect 5700 4750 5800 4760
rect 5850 4750 5950 4760
rect 6650 4750 6750 4760
rect 8000 4750 8250 4760
rect 8300 4750 8400 4760
rect 9000 4750 9050 4760
rect 9300 4750 9350 4760
rect 3350 4740 3400 4750
rect 5100 4740 5150 4750
rect 5300 4740 5400 4750
rect 5700 4740 5800 4750
rect 5900 4740 6000 4750
rect 6650 4740 6750 4750
rect 7850 4740 7950 4750
rect 8000 4740 8250 4750
rect 8300 4740 8350 4750
rect 8800 4740 9000 4750
rect 9250 4740 9300 4750
rect 9850 4740 9900 4750
rect 3350 4730 3400 4740
rect 5100 4730 5150 4740
rect 5300 4730 5400 4740
rect 5700 4730 5800 4740
rect 5900 4730 6000 4740
rect 6650 4730 6750 4740
rect 7850 4730 7950 4740
rect 8000 4730 8250 4740
rect 8300 4730 8350 4740
rect 8800 4730 9000 4740
rect 9250 4730 9300 4740
rect 9850 4730 9900 4740
rect 3350 4720 3400 4730
rect 5100 4720 5150 4730
rect 5300 4720 5400 4730
rect 5700 4720 5800 4730
rect 5900 4720 6000 4730
rect 6650 4720 6750 4730
rect 7850 4720 7950 4730
rect 8000 4720 8250 4730
rect 8300 4720 8350 4730
rect 8800 4720 9000 4730
rect 9250 4720 9300 4730
rect 9850 4720 9900 4730
rect 3350 4710 3400 4720
rect 5100 4710 5150 4720
rect 5300 4710 5400 4720
rect 5700 4710 5800 4720
rect 5900 4710 6000 4720
rect 6650 4710 6750 4720
rect 7850 4710 7950 4720
rect 8000 4710 8250 4720
rect 8300 4710 8350 4720
rect 8800 4710 9000 4720
rect 9250 4710 9300 4720
rect 9850 4710 9900 4720
rect 3350 4700 3400 4710
rect 5100 4700 5150 4710
rect 5300 4700 5400 4710
rect 5700 4700 5800 4710
rect 5900 4700 6000 4710
rect 6650 4700 6750 4710
rect 7850 4700 7950 4710
rect 8000 4700 8250 4710
rect 8300 4700 8350 4710
rect 8800 4700 9000 4710
rect 9250 4700 9300 4710
rect 9850 4700 9900 4710
rect 3350 4690 3400 4700
rect 3450 4690 3500 4700
rect 5300 4690 5350 4700
rect 5800 4690 5950 4700
rect 6650 4690 6750 4700
rect 7350 4690 7400 4700
rect 7750 4690 7850 4700
rect 7900 4690 7950 4700
rect 8000 4690 8100 4700
rect 8600 4690 8650 4700
rect 8950 4690 9000 4700
rect 9800 4690 9850 4700
rect 3350 4680 3400 4690
rect 3450 4680 3500 4690
rect 5300 4680 5350 4690
rect 5800 4680 5950 4690
rect 6650 4680 6750 4690
rect 7350 4680 7400 4690
rect 7750 4680 7850 4690
rect 7900 4680 7950 4690
rect 8000 4680 8100 4690
rect 8600 4680 8650 4690
rect 8950 4680 9000 4690
rect 9800 4680 9850 4690
rect 3350 4670 3400 4680
rect 3450 4670 3500 4680
rect 5300 4670 5350 4680
rect 5800 4670 5950 4680
rect 6650 4670 6750 4680
rect 7350 4670 7400 4680
rect 7750 4670 7850 4680
rect 7900 4670 7950 4680
rect 8000 4670 8100 4680
rect 8600 4670 8650 4680
rect 8950 4670 9000 4680
rect 9800 4670 9850 4680
rect 3350 4660 3400 4670
rect 3450 4660 3500 4670
rect 5300 4660 5350 4670
rect 5800 4660 5950 4670
rect 6650 4660 6750 4670
rect 7350 4660 7400 4670
rect 7750 4660 7850 4670
rect 7900 4660 7950 4670
rect 8000 4660 8100 4670
rect 8600 4660 8650 4670
rect 8950 4660 9000 4670
rect 9800 4660 9850 4670
rect 3350 4650 3400 4660
rect 3450 4650 3500 4660
rect 5300 4650 5350 4660
rect 5800 4650 5950 4660
rect 6650 4650 6750 4660
rect 7350 4650 7400 4660
rect 7750 4650 7850 4660
rect 7900 4650 7950 4660
rect 8000 4650 8100 4660
rect 8600 4650 8650 4660
rect 8950 4650 9000 4660
rect 9800 4650 9850 4660
rect 3300 4640 3450 4650
rect 5200 4640 5250 4650
rect 5300 4640 5350 4650
rect 6650 4640 6750 4650
rect 7350 4640 7400 4650
rect 7500 4640 7650 4650
rect 7750 4640 7800 4650
rect 7900 4640 7950 4650
rect 8300 4640 8350 4650
rect 8500 4640 8550 4650
rect 8950 4640 9000 4650
rect 9750 4640 9800 4650
rect 3300 4630 3450 4640
rect 5200 4630 5250 4640
rect 5300 4630 5350 4640
rect 6650 4630 6750 4640
rect 7350 4630 7400 4640
rect 7500 4630 7650 4640
rect 7750 4630 7800 4640
rect 7900 4630 7950 4640
rect 8300 4630 8350 4640
rect 8500 4630 8550 4640
rect 8950 4630 9000 4640
rect 9750 4630 9800 4640
rect 3300 4620 3450 4630
rect 5200 4620 5250 4630
rect 5300 4620 5350 4630
rect 6650 4620 6750 4630
rect 7350 4620 7400 4630
rect 7500 4620 7650 4630
rect 7750 4620 7800 4630
rect 7900 4620 7950 4630
rect 8300 4620 8350 4630
rect 8500 4620 8550 4630
rect 8950 4620 9000 4630
rect 9750 4620 9800 4630
rect 3300 4610 3450 4620
rect 5200 4610 5250 4620
rect 5300 4610 5350 4620
rect 6650 4610 6750 4620
rect 7350 4610 7400 4620
rect 7500 4610 7650 4620
rect 7750 4610 7800 4620
rect 7900 4610 7950 4620
rect 8300 4610 8350 4620
rect 8500 4610 8550 4620
rect 8950 4610 9000 4620
rect 9750 4610 9800 4620
rect 3300 4600 3450 4610
rect 5200 4600 5250 4610
rect 5300 4600 5350 4610
rect 6650 4600 6750 4610
rect 7350 4600 7400 4610
rect 7500 4600 7650 4610
rect 7750 4600 7800 4610
rect 7900 4600 7950 4610
rect 8300 4600 8350 4610
rect 8500 4600 8550 4610
rect 8950 4600 9000 4610
rect 9750 4600 9800 4610
rect 3250 4590 3450 4600
rect 5250 4590 5400 4600
rect 5800 4590 6050 4600
rect 6600 4590 6750 4600
rect 7300 4590 7400 4600
rect 7500 4590 7550 4600
rect 7600 4590 7650 4600
rect 8150 4590 8200 4600
rect 8300 4590 8400 4600
rect 8500 4590 8600 4600
rect 8950 4590 9000 4600
rect 9200 4590 9250 4600
rect 9700 4590 9750 4600
rect 3250 4580 3450 4590
rect 5250 4580 5400 4590
rect 5800 4580 6050 4590
rect 6600 4580 6750 4590
rect 7300 4580 7400 4590
rect 7500 4580 7550 4590
rect 7600 4580 7650 4590
rect 8150 4580 8200 4590
rect 8300 4580 8400 4590
rect 8500 4580 8600 4590
rect 8950 4580 9000 4590
rect 9200 4580 9250 4590
rect 9700 4580 9750 4590
rect 3250 4570 3450 4580
rect 5250 4570 5400 4580
rect 5800 4570 6050 4580
rect 6600 4570 6750 4580
rect 7300 4570 7400 4580
rect 7500 4570 7550 4580
rect 7600 4570 7650 4580
rect 8150 4570 8200 4580
rect 8300 4570 8400 4580
rect 8500 4570 8600 4580
rect 8950 4570 9000 4580
rect 9200 4570 9250 4580
rect 9700 4570 9750 4580
rect 3250 4560 3450 4570
rect 5250 4560 5400 4570
rect 5800 4560 6050 4570
rect 6600 4560 6750 4570
rect 7300 4560 7400 4570
rect 7500 4560 7550 4570
rect 7600 4560 7650 4570
rect 8150 4560 8200 4570
rect 8300 4560 8400 4570
rect 8500 4560 8600 4570
rect 8950 4560 9000 4570
rect 9200 4560 9250 4570
rect 9700 4560 9750 4570
rect 3250 4550 3450 4560
rect 5250 4550 5400 4560
rect 5800 4550 6050 4560
rect 6600 4550 6750 4560
rect 7300 4550 7400 4560
rect 7500 4550 7550 4560
rect 7600 4550 7650 4560
rect 8150 4550 8200 4560
rect 8300 4550 8400 4560
rect 8500 4550 8600 4560
rect 8950 4550 9000 4560
rect 9200 4550 9250 4560
rect 9700 4550 9750 4560
rect 3250 4540 3300 4550
rect 5350 4540 5450 4550
rect 5850 4540 5900 4550
rect 6100 4540 6200 4550
rect 6550 4540 6700 4550
rect 7300 4540 7400 4550
rect 7900 4540 7950 4550
rect 8000 4540 8250 4550
rect 8300 4540 8400 4550
rect 9200 4540 9250 4550
rect 9650 4540 9700 4550
rect 3250 4530 3300 4540
rect 5350 4530 5450 4540
rect 5850 4530 5900 4540
rect 6100 4530 6200 4540
rect 6550 4530 6700 4540
rect 7300 4530 7400 4540
rect 7900 4530 7950 4540
rect 8000 4530 8250 4540
rect 8300 4530 8400 4540
rect 9200 4530 9250 4540
rect 9650 4530 9700 4540
rect 3250 4520 3300 4530
rect 5350 4520 5450 4530
rect 5850 4520 5900 4530
rect 6100 4520 6200 4530
rect 6550 4520 6700 4530
rect 7300 4520 7400 4530
rect 7900 4520 7950 4530
rect 8000 4520 8250 4530
rect 8300 4520 8400 4530
rect 9200 4520 9250 4530
rect 9650 4520 9700 4530
rect 3250 4510 3300 4520
rect 5350 4510 5450 4520
rect 5850 4510 5900 4520
rect 6100 4510 6200 4520
rect 6550 4510 6700 4520
rect 7300 4510 7400 4520
rect 7900 4510 7950 4520
rect 8000 4510 8250 4520
rect 8300 4510 8400 4520
rect 9200 4510 9250 4520
rect 9650 4510 9700 4520
rect 3250 4500 3300 4510
rect 5350 4500 5450 4510
rect 5850 4500 5900 4510
rect 6100 4500 6200 4510
rect 6550 4500 6700 4510
rect 7300 4500 7400 4510
rect 7900 4500 7950 4510
rect 8000 4500 8250 4510
rect 8300 4500 8400 4510
rect 9200 4500 9250 4510
rect 9650 4500 9700 4510
rect 5600 4490 5700 4500
rect 5850 4490 5950 4500
rect 6100 4490 6150 4500
rect 6550 4490 6700 4500
rect 7350 4490 7400 4500
rect 7800 4490 7850 4500
rect 7900 4490 8050 4500
rect 8100 4490 8250 4500
rect 8900 4490 8950 4500
rect 9600 4490 9650 4500
rect 5600 4480 5700 4490
rect 5850 4480 5950 4490
rect 6100 4480 6150 4490
rect 6550 4480 6700 4490
rect 7350 4480 7400 4490
rect 7800 4480 7850 4490
rect 7900 4480 8050 4490
rect 8100 4480 8250 4490
rect 8900 4480 8950 4490
rect 9600 4480 9650 4490
rect 5600 4470 5700 4480
rect 5850 4470 5950 4480
rect 6100 4470 6150 4480
rect 6550 4470 6700 4480
rect 7350 4470 7400 4480
rect 7800 4470 7850 4480
rect 7900 4470 8050 4480
rect 8100 4470 8250 4480
rect 8900 4470 8950 4480
rect 9600 4470 9650 4480
rect 5600 4460 5700 4470
rect 5850 4460 5950 4470
rect 6100 4460 6150 4470
rect 6550 4460 6700 4470
rect 7350 4460 7400 4470
rect 7800 4460 7850 4470
rect 7900 4460 8050 4470
rect 8100 4460 8250 4470
rect 8900 4460 8950 4470
rect 9600 4460 9650 4470
rect 5600 4450 5700 4460
rect 5850 4450 5950 4460
rect 6100 4450 6150 4460
rect 6550 4450 6700 4460
rect 7350 4450 7400 4460
rect 7800 4450 7850 4460
rect 7900 4450 8050 4460
rect 8100 4450 8250 4460
rect 8900 4450 8950 4460
rect 9600 4450 9650 4460
rect 3000 4440 3050 4450
rect 3300 4440 3400 4450
rect 5600 4440 5750 4450
rect 6550 4440 6700 4450
rect 7350 4440 7400 4450
rect 7800 4440 7850 4450
rect 7900 4440 8000 4450
rect 8850 4440 8900 4450
rect 9550 4440 9600 4450
rect 3000 4430 3050 4440
rect 3300 4430 3400 4440
rect 5600 4430 5750 4440
rect 6550 4430 6700 4440
rect 7350 4430 7400 4440
rect 7800 4430 7850 4440
rect 7900 4430 8000 4440
rect 8850 4430 8900 4440
rect 9550 4430 9600 4440
rect 3000 4420 3050 4430
rect 3300 4420 3400 4430
rect 5600 4420 5750 4430
rect 6550 4420 6700 4430
rect 7350 4420 7400 4430
rect 7800 4420 7850 4430
rect 7900 4420 8000 4430
rect 8850 4420 8900 4430
rect 9550 4420 9600 4430
rect 3000 4410 3050 4420
rect 3300 4410 3400 4420
rect 5600 4410 5750 4420
rect 6550 4410 6700 4420
rect 7350 4410 7400 4420
rect 7800 4410 7850 4420
rect 7900 4410 8000 4420
rect 8850 4410 8900 4420
rect 9550 4410 9600 4420
rect 3000 4400 3050 4410
rect 3300 4400 3400 4410
rect 5600 4400 5750 4410
rect 6550 4400 6700 4410
rect 7350 4400 7400 4410
rect 7800 4400 7850 4410
rect 7900 4400 8000 4410
rect 8850 4400 8900 4410
rect 9550 4400 9600 4410
rect 3000 4390 3050 4400
rect 5350 4390 5400 4400
rect 5600 4390 5950 4400
rect 6500 4390 6700 4400
rect 7300 4390 7400 4400
rect 8850 4390 8900 4400
rect 9150 4390 9200 4400
rect 9500 4390 9550 4400
rect 9800 4390 9850 4400
rect 3000 4380 3050 4390
rect 5350 4380 5400 4390
rect 5600 4380 5950 4390
rect 6500 4380 6700 4390
rect 7300 4380 7400 4390
rect 8850 4380 8900 4390
rect 9150 4380 9200 4390
rect 9500 4380 9550 4390
rect 9800 4380 9850 4390
rect 3000 4370 3050 4380
rect 5350 4370 5400 4380
rect 5600 4370 5950 4380
rect 6500 4370 6700 4380
rect 7300 4370 7400 4380
rect 8850 4370 8900 4380
rect 9150 4370 9200 4380
rect 9500 4370 9550 4380
rect 9800 4370 9850 4380
rect 3000 4360 3050 4370
rect 5350 4360 5400 4370
rect 5600 4360 5950 4370
rect 6500 4360 6700 4370
rect 7300 4360 7400 4370
rect 8850 4360 8900 4370
rect 9150 4360 9200 4370
rect 9500 4360 9550 4370
rect 9800 4360 9850 4370
rect 3000 4350 3050 4360
rect 5350 4350 5400 4360
rect 5600 4350 5950 4360
rect 6500 4350 6700 4360
rect 7300 4350 7400 4360
rect 8850 4350 8900 4360
rect 9150 4350 9200 4360
rect 9500 4350 9550 4360
rect 9800 4350 9850 4360
rect 4600 4340 4850 4350
rect 5350 4340 5400 4350
rect 5500 4340 5950 4350
rect 6500 4340 6650 4350
rect 7250 4340 7350 4350
rect 8850 4340 8900 4350
rect 9150 4340 9200 4350
rect 9450 4340 9500 4350
rect 9800 4340 9990 4350
rect 4600 4330 4850 4340
rect 5350 4330 5400 4340
rect 5500 4330 5950 4340
rect 6500 4330 6650 4340
rect 7250 4330 7350 4340
rect 8850 4330 8900 4340
rect 9150 4330 9200 4340
rect 9450 4330 9500 4340
rect 9800 4330 9990 4340
rect 4600 4320 4850 4330
rect 5350 4320 5400 4330
rect 5500 4320 5950 4330
rect 6500 4320 6650 4330
rect 7250 4320 7350 4330
rect 8850 4320 8900 4330
rect 9150 4320 9200 4330
rect 9450 4320 9500 4330
rect 9800 4320 9990 4330
rect 4600 4310 4850 4320
rect 5350 4310 5400 4320
rect 5500 4310 5950 4320
rect 6500 4310 6650 4320
rect 7250 4310 7350 4320
rect 8850 4310 8900 4320
rect 9150 4310 9200 4320
rect 9450 4310 9500 4320
rect 9800 4310 9990 4320
rect 4600 4300 4850 4310
rect 5350 4300 5400 4310
rect 5500 4300 5950 4310
rect 6500 4300 6650 4310
rect 7250 4300 7350 4310
rect 8850 4300 8900 4310
rect 9150 4300 9200 4310
rect 9450 4300 9500 4310
rect 9800 4300 9990 4310
rect 4600 4290 4650 4300
rect 4800 4290 4900 4300
rect 5350 4290 5450 4300
rect 5550 4290 5950 4300
rect 6450 4290 6500 4300
rect 6600 4290 6650 4300
rect 7050 4290 7150 4300
rect 8450 4290 8500 4300
rect 9150 4290 9200 4300
rect 9400 4290 9450 4300
rect 9800 4290 9990 4300
rect 4600 4280 4650 4290
rect 4800 4280 4900 4290
rect 5350 4280 5450 4290
rect 5550 4280 5950 4290
rect 6450 4280 6500 4290
rect 6600 4280 6650 4290
rect 7050 4280 7150 4290
rect 8450 4280 8500 4290
rect 9150 4280 9200 4290
rect 9400 4280 9450 4290
rect 9800 4280 9990 4290
rect 4600 4270 4650 4280
rect 4800 4270 4900 4280
rect 5350 4270 5450 4280
rect 5550 4270 5950 4280
rect 6450 4270 6500 4280
rect 6600 4270 6650 4280
rect 7050 4270 7150 4280
rect 8450 4270 8500 4280
rect 9150 4270 9200 4280
rect 9400 4270 9450 4280
rect 9800 4270 9990 4280
rect 4600 4260 4650 4270
rect 4800 4260 4900 4270
rect 5350 4260 5450 4270
rect 5550 4260 5950 4270
rect 6450 4260 6500 4270
rect 6600 4260 6650 4270
rect 7050 4260 7150 4270
rect 8450 4260 8500 4270
rect 9150 4260 9200 4270
rect 9400 4260 9450 4270
rect 9800 4260 9990 4270
rect 4600 4250 4650 4260
rect 4800 4250 4900 4260
rect 5350 4250 5450 4260
rect 5550 4250 5950 4260
rect 6450 4250 6500 4260
rect 6600 4250 6650 4260
rect 7050 4250 7150 4260
rect 8450 4250 8500 4260
rect 9150 4250 9200 4260
rect 9400 4250 9450 4260
rect 9800 4250 9990 4260
rect 4200 4240 4300 4250
rect 4550 4240 4650 4250
rect 4750 4240 4900 4250
rect 5450 4240 5500 4250
rect 5600 4240 5650 4250
rect 5700 4240 6000 4250
rect 6350 4240 6500 4250
rect 6600 4240 6650 4250
rect 7100 4240 7150 4250
rect 7400 4240 7450 4250
rect 9150 4240 9200 4250
rect 9350 4240 9400 4250
rect 9700 4240 9750 4250
rect 9850 4240 9990 4250
rect 4200 4230 4300 4240
rect 4550 4230 4650 4240
rect 4750 4230 4900 4240
rect 5450 4230 5500 4240
rect 5600 4230 5650 4240
rect 5700 4230 6000 4240
rect 6350 4230 6500 4240
rect 6600 4230 6650 4240
rect 7100 4230 7150 4240
rect 7400 4230 7450 4240
rect 9150 4230 9200 4240
rect 9350 4230 9400 4240
rect 9700 4230 9750 4240
rect 9850 4230 9990 4240
rect 4200 4220 4300 4230
rect 4550 4220 4650 4230
rect 4750 4220 4900 4230
rect 5450 4220 5500 4230
rect 5600 4220 5650 4230
rect 5700 4220 6000 4230
rect 6350 4220 6500 4230
rect 6600 4220 6650 4230
rect 7100 4220 7150 4230
rect 7400 4220 7450 4230
rect 9150 4220 9200 4230
rect 9350 4220 9400 4230
rect 9700 4220 9750 4230
rect 9850 4220 9990 4230
rect 4200 4210 4300 4220
rect 4550 4210 4650 4220
rect 4750 4210 4900 4220
rect 5450 4210 5500 4220
rect 5600 4210 5650 4220
rect 5700 4210 6000 4220
rect 6350 4210 6500 4220
rect 6600 4210 6650 4220
rect 7100 4210 7150 4220
rect 7400 4210 7450 4220
rect 9150 4210 9200 4220
rect 9350 4210 9400 4220
rect 9700 4210 9750 4220
rect 9850 4210 9990 4220
rect 4200 4200 4300 4210
rect 4550 4200 4650 4210
rect 4750 4200 4900 4210
rect 5450 4200 5500 4210
rect 5600 4200 5650 4210
rect 5700 4200 6000 4210
rect 6350 4200 6500 4210
rect 6600 4200 6650 4210
rect 7100 4200 7150 4210
rect 7400 4200 7450 4210
rect 9150 4200 9200 4210
rect 9350 4200 9400 4210
rect 9700 4200 9750 4210
rect 9850 4200 9990 4210
rect 4150 4190 4200 4200
rect 4300 4190 4350 4200
rect 4500 4190 4650 4200
rect 4700 4190 4950 4200
rect 5400 4190 5500 4200
rect 5600 4190 5700 4200
rect 5900 4190 6450 4200
rect 6600 4190 6650 4200
rect 7200 4190 7250 4200
rect 7350 4190 7450 4200
rect 8800 4190 8850 4200
rect 9200 4190 9350 4200
rect 9650 4190 9800 4200
rect 9900 4190 9990 4200
rect 4150 4180 4200 4190
rect 4300 4180 4350 4190
rect 4500 4180 4650 4190
rect 4700 4180 4950 4190
rect 5400 4180 5500 4190
rect 5600 4180 5700 4190
rect 5900 4180 6450 4190
rect 6600 4180 6650 4190
rect 7200 4180 7250 4190
rect 7350 4180 7450 4190
rect 8800 4180 8850 4190
rect 9200 4180 9350 4190
rect 9650 4180 9800 4190
rect 9900 4180 9990 4190
rect 4150 4170 4200 4180
rect 4300 4170 4350 4180
rect 4500 4170 4650 4180
rect 4700 4170 4950 4180
rect 5400 4170 5500 4180
rect 5600 4170 5700 4180
rect 5900 4170 6450 4180
rect 6600 4170 6650 4180
rect 7200 4170 7250 4180
rect 7350 4170 7450 4180
rect 8800 4170 8850 4180
rect 9200 4170 9350 4180
rect 9650 4170 9800 4180
rect 9900 4170 9990 4180
rect 4150 4160 4200 4170
rect 4300 4160 4350 4170
rect 4500 4160 4650 4170
rect 4700 4160 4950 4170
rect 5400 4160 5500 4170
rect 5600 4160 5700 4170
rect 5900 4160 6450 4170
rect 6600 4160 6650 4170
rect 7200 4160 7250 4170
rect 7350 4160 7450 4170
rect 8800 4160 8850 4170
rect 9200 4160 9350 4170
rect 9650 4160 9800 4170
rect 9900 4160 9990 4170
rect 4150 4150 4200 4160
rect 4300 4150 4350 4160
rect 4500 4150 4650 4160
rect 4700 4150 4950 4160
rect 5400 4150 5500 4160
rect 5600 4150 5700 4160
rect 5900 4150 6450 4160
rect 6600 4150 6650 4160
rect 7200 4150 7250 4160
rect 7350 4150 7450 4160
rect 8800 4150 8850 4160
rect 9200 4150 9350 4160
rect 9650 4150 9800 4160
rect 9900 4150 9990 4160
rect 4100 4140 4200 4150
rect 4350 4140 4550 4150
rect 5450 4140 5500 4150
rect 5650 4140 5700 4150
rect 5950 4140 6400 4150
rect 6550 4140 6650 4150
rect 7200 4140 7250 4150
rect 8800 4140 8850 4150
rect 9750 4140 9850 4150
rect 4100 4130 4200 4140
rect 4350 4130 4550 4140
rect 5450 4130 5500 4140
rect 5650 4130 5700 4140
rect 5950 4130 6400 4140
rect 6550 4130 6650 4140
rect 7200 4130 7250 4140
rect 8800 4130 8850 4140
rect 9750 4130 9850 4140
rect 4100 4120 4200 4130
rect 4350 4120 4550 4130
rect 5450 4120 5500 4130
rect 5650 4120 5700 4130
rect 5950 4120 6400 4130
rect 6550 4120 6650 4130
rect 7200 4120 7250 4130
rect 8800 4120 8850 4130
rect 9750 4120 9850 4130
rect 4100 4110 4200 4120
rect 4350 4110 4550 4120
rect 5450 4110 5500 4120
rect 5650 4110 5700 4120
rect 5950 4110 6400 4120
rect 6550 4110 6650 4120
rect 7200 4110 7250 4120
rect 8800 4110 8850 4120
rect 9750 4110 9850 4120
rect 4100 4100 4200 4110
rect 4350 4100 4550 4110
rect 5450 4100 5500 4110
rect 5650 4100 5700 4110
rect 5950 4100 6400 4110
rect 6550 4100 6650 4110
rect 7200 4100 7250 4110
rect 8800 4100 8850 4110
rect 9750 4100 9850 4110
rect 3200 4090 3250 4100
rect 4100 4090 4150 4100
rect 4450 4090 4550 4100
rect 4850 4090 5050 4100
rect 5450 4090 5500 4100
rect 5750 4090 6300 4100
rect 6450 4090 6650 4100
rect 9600 4090 9700 4100
rect 9800 4090 9950 4100
rect 3200 4080 3250 4090
rect 4100 4080 4150 4090
rect 4450 4080 4550 4090
rect 4850 4080 5050 4090
rect 5450 4080 5500 4090
rect 5750 4080 6300 4090
rect 6450 4080 6650 4090
rect 9600 4080 9700 4090
rect 9800 4080 9950 4090
rect 3200 4070 3250 4080
rect 4100 4070 4150 4080
rect 4450 4070 4550 4080
rect 4850 4070 5050 4080
rect 5450 4070 5500 4080
rect 5750 4070 6300 4080
rect 6450 4070 6650 4080
rect 9600 4070 9700 4080
rect 9800 4070 9950 4080
rect 3200 4060 3250 4070
rect 4100 4060 4150 4070
rect 4450 4060 4550 4070
rect 4850 4060 5050 4070
rect 5450 4060 5500 4070
rect 5750 4060 6300 4070
rect 6450 4060 6650 4070
rect 9600 4060 9700 4070
rect 9800 4060 9950 4070
rect 3200 4050 3250 4060
rect 4100 4050 4150 4060
rect 4450 4050 4550 4060
rect 4850 4050 5050 4060
rect 5450 4050 5500 4060
rect 5750 4050 6300 4060
rect 6450 4050 6650 4060
rect 9600 4050 9700 4060
rect 9800 4050 9950 4060
rect 3200 4040 3250 4050
rect 4050 4040 4100 4050
rect 4150 4040 4300 4050
rect 4500 4040 4550 4050
rect 4750 4040 4900 4050
rect 5000 4040 5100 4050
rect 5400 4040 5500 4050
rect 6050 4040 6200 4050
rect 6400 4040 6650 4050
rect 7150 4040 7200 4050
rect 3200 4030 3250 4040
rect 4050 4030 4100 4040
rect 4150 4030 4300 4040
rect 4500 4030 4550 4040
rect 4750 4030 4900 4040
rect 5000 4030 5100 4040
rect 5400 4030 5500 4040
rect 6050 4030 6200 4040
rect 6400 4030 6650 4040
rect 7150 4030 7200 4040
rect 3200 4020 3250 4030
rect 4050 4020 4100 4030
rect 4150 4020 4300 4030
rect 4500 4020 4550 4030
rect 4750 4020 4900 4030
rect 5000 4020 5100 4030
rect 5400 4020 5500 4030
rect 6050 4020 6200 4030
rect 6400 4020 6650 4030
rect 7150 4020 7200 4030
rect 3200 4010 3250 4020
rect 4050 4010 4100 4020
rect 4150 4010 4300 4020
rect 4500 4010 4550 4020
rect 4750 4010 4900 4020
rect 5000 4010 5100 4020
rect 5400 4010 5500 4020
rect 6050 4010 6200 4020
rect 6400 4010 6650 4020
rect 7150 4010 7200 4020
rect 3200 4000 3250 4010
rect 4050 4000 4100 4010
rect 4150 4000 4300 4010
rect 4500 4000 4550 4010
rect 4750 4000 4900 4010
rect 5000 4000 5100 4010
rect 5400 4000 5500 4010
rect 6050 4000 6200 4010
rect 6400 4000 6650 4010
rect 7150 4000 7200 4010
rect 3200 3990 3250 4000
rect 4000 3990 4050 4000
rect 4100 3990 4150 4000
rect 4300 3990 4350 4000
rect 4500 3990 4550 4000
rect 4700 3990 4850 4000
rect 5050 3990 5100 4000
rect 6400 3990 6600 4000
rect 7100 3990 7150 4000
rect 8350 3990 8400 4000
rect 8450 3990 8500 4000
rect 8550 3990 8650 4000
rect 3200 3980 3250 3990
rect 4000 3980 4050 3990
rect 4100 3980 4150 3990
rect 4300 3980 4350 3990
rect 4500 3980 4550 3990
rect 4700 3980 4850 3990
rect 5050 3980 5100 3990
rect 6400 3980 6600 3990
rect 7100 3980 7150 3990
rect 8350 3980 8400 3990
rect 8450 3980 8500 3990
rect 8550 3980 8650 3990
rect 3200 3970 3250 3980
rect 4000 3970 4050 3980
rect 4100 3970 4150 3980
rect 4300 3970 4350 3980
rect 4500 3970 4550 3980
rect 4700 3970 4850 3980
rect 5050 3970 5100 3980
rect 6400 3970 6600 3980
rect 7100 3970 7150 3980
rect 8350 3970 8400 3980
rect 8450 3970 8500 3980
rect 8550 3970 8650 3980
rect 3200 3960 3250 3970
rect 4000 3960 4050 3970
rect 4100 3960 4150 3970
rect 4300 3960 4350 3970
rect 4500 3960 4550 3970
rect 4700 3960 4850 3970
rect 5050 3960 5100 3970
rect 6400 3960 6600 3970
rect 7100 3960 7150 3970
rect 8350 3960 8400 3970
rect 8450 3960 8500 3970
rect 8550 3960 8650 3970
rect 3200 3950 3250 3960
rect 4000 3950 4050 3960
rect 4100 3950 4150 3960
rect 4300 3950 4350 3960
rect 4500 3950 4550 3960
rect 4700 3950 4850 3960
rect 5050 3950 5100 3960
rect 6400 3950 6600 3960
rect 7100 3950 7150 3960
rect 8350 3950 8400 3960
rect 8450 3950 8500 3960
rect 8550 3950 8650 3960
rect 3950 3940 4100 3950
rect 4550 3940 4800 3950
rect 5100 3940 5150 3950
rect 6450 3940 6600 3950
rect 7100 3940 7150 3950
rect 8200 3940 8350 3950
rect 8400 3940 8500 3950
rect 8700 3940 8750 3950
rect 9550 3940 9650 3950
rect 9750 3940 9800 3950
rect 3950 3930 4100 3940
rect 4550 3930 4800 3940
rect 5100 3930 5150 3940
rect 6450 3930 6600 3940
rect 7100 3930 7150 3940
rect 8200 3930 8350 3940
rect 8400 3930 8500 3940
rect 8700 3930 8750 3940
rect 9550 3930 9650 3940
rect 9750 3930 9800 3940
rect 3950 3920 4100 3930
rect 4550 3920 4800 3930
rect 5100 3920 5150 3930
rect 6450 3920 6600 3930
rect 7100 3920 7150 3930
rect 8200 3920 8350 3930
rect 8400 3920 8500 3930
rect 8700 3920 8750 3930
rect 9550 3920 9650 3930
rect 9750 3920 9800 3930
rect 3950 3910 4100 3920
rect 4550 3910 4800 3920
rect 5100 3910 5150 3920
rect 6450 3910 6600 3920
rect 7100 3910 7150 3920
rect 8200 3910 8350 3920
rect 8400 3910 8500 3920
rect 8700 3910 8750 3920
rect 9550 3910 9650 3920
rect 9750 3910 9800 3920
rect 3950 3900 4100 3910
rect 4550 3900 4800 3910
rect 5100 3900 5150 3910
rect 6450 3900 6600 3910
rect 7100 3900 7150 3910
rect 8200 3900 8350 3910
rect 8400 3900 8500 3910
rect 8700 3900 8750 3910
rect 9550 3900 9650 3910
rect 9750 3900 9800 3910
rect 3200 3890 3250 3900
rect 3900 3890 4050 3900
rect 4350 3890 4400 3900
rect 4550 3890 4650 3900
rect 5150 3890 5200 3900
rect 6500 3890 6600 3900
rect 7100 3890 7150 3900
rect 8200 3890 8300 3900
rect 8400 3890 8550 3900
rect 9450 3890 9550 3900
rect 9750 3890 9850 3900
rect 3200 3880 3250 3890
rect 3900 3880 4050 3890
rect 4350 3880 4400 3890
rect 4550 3880 4650 3890
rect 5150 3880 5200 3890
rect 6500 3880 6600 3890
rect 7100 3880 7150 3890
rect 8200 3880 8300 3890
rect 8400 3880 8550 3890
rect 9450 3880 9550 3890
rect 9750 3880 9850 3890
rect 3200 3870 3250 3880
rect 3900 3870 4050 3880
rect 4350 3870 4400 3880
rect 4550 3870 4650 3880
rect 5150 3870 5200 3880
rect 6500 3870 6600 3880
rect 7100 3870 7150 3880
rect 8200 3870 8300 3880
rect 8400 3870 8550 3880
rect 9450 3870 9550 3880
rect 9750 3870 9850 3880
rect 3200 3860 3250 3870
rect 3900 3860 4050 3870
rect 4350 3860 4400 3870
rect 4550 3860 4650 3870
rect 5150 3860 5200 3870
rect 6500 3860 6600 3870
rect 7100 3860 7150 3870
rect 8200 3860 8300 3870
rect 8400 3860 8550 3870
rect 9450 3860 9550 3870
rect 9750 3860 9850 3870
rect 3200 3850 3250 3860
rect 3900 3850 4050 3860
rect 4350 3850 4400 3860
rect 4550 3850 4650 3860
rect 5150 3850 5200 3860
rect 6500 3850 6600 3860
rect 7100 3850 7150 3860
rect 8200 3850 8300 3860
rect 8400 3850 8550 3860
rect 9450 3850 9550 3860
rect 9750 3850 9850 3860
rect 3200 3840 3250 3850
rect 3900 3840 4000 3850
rect 4350 3840 4400 3850
rect 5150 3840 5200 3850
rect 6550 3840 6600 3850
rect 7050 3840 7100 3850
rect 8250 3840 8700 3850
rect 9550 3840 9600 3850
rect 9800 3840 9900 3850
rect 3200 3830 3250 3840
rect 3900 3830 4000 3840
rect 4350 3830 4400 3840
rect 5150 3830 5200 3840
rect 6550 3830 6600 3840
rect 7050 3830 7100 3840
rect 8250 3830 8700 3840
rect 9550 3830 9600 3840
rect 9800 3830 9900 3840
rect 3200 3820 3250 3830
rect 3900 3820 4000 3830
rect 4350 3820 4400 3830
rect 5150 3820 5200 3830
rect 6550 3820 6600 3830
rect 7050 3820 7100 3830
rect 8250 3820 8700 3830
rect 9550 3820 9600 3830
rect 9800 3820 9900 3830
rect 3200 3810 3250 3820
rect 3900 3810 4000 3820
rect 4350 3810 4400 3820
rect 5150 3810 5200 3820
rect 6550 3810 6600 3820
rect 7050 3810 7100 3820
rect 8250 3810 8700 3820
rect 9550 3810 9600 3820
rect 9800 3810 9900 3820
rect 3200 3800 3250 3810
rect 3900 3800 4000 3810
rect 4350 3800 4400 3810
rect 5150 3800 5200 3810
rect 6550 3800 6600 3810
rect 7050 3800 7100 3810
rect 8250 3800 8700 3810
rect 9550 3800 9600 3810
rect 9800 3800 9900 3810
rect 3200 3790 3250 3800
rect 4300 3790 4450 3800
rect 4850 3790 4900 3800
rect 5150 3790 5200 3800
rect 6550 3790 6600 3800
rect 8350 3790 8550 3800
rect 9600 3790 9650 3800
rect 9850 3790 9900 3800
rect 3200 3780 3250 3790
rect 4300 3780 4450 3790
rect 4850 3780 4900 3790
rect 5150 3780 5200 3790
rect 6550 3780 6600 3790
rect 8350 3780 8550 3790
rect 9600 3780 9650 3790
rect 9850 3780 9900 3790
rect 3200 3770 3250 3780
rect 4300 3770 4450 3780
rect 4850 3770 4900 3780
rect 5150 3770 5200 3780
rect 6550 3770 6600 3780
rect 8350 3770 8550 3780
rect 9600 3770 9650 3780
rect 9850 3770 9900 3780
rect 3200 3760 3250 3770
rect 4300 3760 4450 3770
rect 4850 3760 4900 3770
rect 5150 3760 5200 3770
rect 6550 3760 6600 3770
rect 8350 3760 8550 3770
rect 9600 3760 9650 3770
rect 9850 3760 9900 3770
rect 3200 3750 3250 3760
rect 4300 3750 4450 3760
rect 4850 3750 4900 3760
rect 5150 3750 5200 3760
rect 6550 3750 6600 3760
rect 8350 3750 8550 3760
rect 9600 3750 9650 3760
rect 9850 3750 9900 3760
rect 3200 3740 3250 3750
rect 4050 3740 4150 3750
rect 4250 3740 4450 3750
rect 4800 3740 4850 3750
rect 4950 3740 5250 3750
rect 6550 3740 6600 3750
rect 7000 3740 7050 3750
rect 8450 3740 8550 3750
rect 9650 3740 9990 3750
rect 3200 3730 3250 3740
rect 4050 3730 4150 3740
rect 4250 3730 4450 3740
rect 4800 3730 4850 3740
rect 4950 3730 5250 3740
rect 6550 3730 6600 3740
rect 7000 3730 7050 3740
rect 8450 3730 8550 3740
rect 9650 3730 9990 3740
rect 3200 3720 3250 3730
rect 4050 3720 4150 3730
rect 4250 3720 4450 3730
rect 4800 3720 4850 3730
rect 4950 3720 5250 3730
rect 6550 3720 6600 3730
rect 7000 3720 7050 3730
rect 8450 3720 8550 3730
rect 9650 3720 9990 3730
rect 3200 3710 3250 3720
rect 4050 3710 4150 3720
rect 4250 3710 4450 3720
rect 4800 3710 4850 3720
rect 4950 3710 5250 3720
rect 6550 3710 6600 3720
rect 7000 3710 7050 3720
rect 8450 3710 8550 3720
rect 9650 3710 9990 3720
rect 3200 3700 3250 3710
rect 4050 3700 4150 3710
rect 4250 3700 4450 3710
rect 4800 3700 4850 3710
rect 4950 3700 5250 3710
rect 6550 3700 6600 3710
rect 7000 3700 7050 3710
rect 8450 3700 8550 3710
rect 9650 3700 9990 3710
rect 3150 3690 3200 3700
rect 4000 3690 4250 3700
rect 4300 3690 4450 3700
rect 4800 3690 4850 3700
rect 5100 3690 5250 3700
rect 6550 3690 6600 3700
rect 6950 3690 7000 3700
rect 8200 3690 8250 3700
rect 8350 3690 8400 3700
rect 8500 3690 8550 3700
rect 8600 3690 8650 3700
rect 9550 3690 9650 3700
rect 9850 3690 9950 3700
rect 3150 3680 3200 3690
rect 4000 3680 4250 3690
rect 4300 3680 4450 3690
rect 4800 3680 4850 3690
rect 5100 3680 5250 3690
rect 6550 3680 6600 3690
rect 6950 3680 7000 3690
rect 8200 3680 8250 3690
rect 8350 3680 8400 3690
rect 8500 3680 8550 3690
rect 8600 3680 8650 3690
rect 9550 3680 9650 3690
rect 9850 3680 9950 3690
rect 3150 3670 3200 3680
rect 4000 3670 4250 3680
rect 4300 3670 4450 3680
rect 4800 3670 4850 3680
rect 5100 3670 5250 3680
rect 6550 3670 6600 3680
rect 6950 3670 7000 3680
rect 8200 3670 8250 3680
rect 8350 3670 8400 3680
rect 8500 3670 8550 3680
rect 8600 3670 8650 3680
rect 9550 3670 9650 3680
rect 9850 3670 9950 3680
rect 3150 3660 3200 3670
rect 4000 3660 4250 3670
rect 4300 3660 4450 3670
rect 4800 3660 4850 3670
rect 5100 3660 5250 3670
rect 6550 3660 6600 3670
rect 6950 3660 7000 3670
rect 8200 3660 8250 3670
rect 8350 3660 8400 3670
rect 8500 3660 8550 3670
rect 8600 3660 8650 3670
rect 9550 3660 9650 3670
rect 9850 3660 9950 3670
rect 3150 3650 3200 3660
rect 4000 3650 4250 3660
rect 4300 3650 4450 3660
rect 4800 3650 4850 3660
rect 5100 3650 5250 3660
rect 6550 3650 6600 3660
rect 6950 3650 7000 3660
rect 8200 3650 8250 3660
rect 8350 3650 8400 3660
rect 8500 3650 8550 3660
rect 8600 3650 8650 3660
rect 9550 3650 9650 3660
rect 9850 3650 9950 3660
rect 4000 3640 4050 3650
rect 4350 3640 4450 3650
rect 4800 3640 4950 3650
rect 5150 3640 5250 3650
rect 6550 3640 6600 3650
rect 6900 3640 6950 3650
rect 8250 3640 8350 3650
rect 9450 3640 9550 3650
rect 9650 3640 9700 3650
rect 9850 3640 9950 3650
rect 4000 3630 4050 3640
rect 4350 3630 4450 3640
rect 4800 3630 4950 3640
rect 5150 3630 5250 3640
rect 6550 3630 6600 3640
rect 6900 3630 6950 3640
rect 8250 3630 8350 3640
rect 9450 3630 9550 3640
rect 9650 3630 9700 3640
rect 9850 3630 9950 3640
rect 4000 3620 4050 3630
rect 4350 3620 4450 3630
rect 4800 3620 4950 3630
rect 5150 3620 5250 3630
rect 6550 3620 6600 3630
rect 6900 3620 6950 3630
rect 8250 3620 8350 3630
rect 9450 3620 9550 3630
rect 9650 3620 9700 3630
rect 9850 3620 9950 3630
rect 4000 3610 4050 3620
rect 4350 3610 4450 3620
rect 4800 3610 4950 3620
rect 5150 3610 5250 3620
rect 6550 3610 6600 3620
rect 6900 3610 6950 3620
rect 8250 3610 8350 3620
rect 9450 3610 9550 3620
rect 9650 3610 9700 3620
rect 9850 3610 9950 3620
rect 4000 3600 4050 3610
rect 4350 3600 4450 3610
rect 4800 3600 4950 3610
rect 5150 3600 5250 3610
rect 6550 3600 6600 3610
rect 6900 3600 6950 3610
rect 8250 3600 8350 3610
rect 9450 3600 9550 3610
rect 9650 3600 9700 3610
rect 9850 3600 9950 3610
rect 4000 3590 4050 3600
rect 4300 3590 4500 3600
rect 4650 3590 4750 3600
rect 4800 3590 4850 3600
rect 4950 3590 5050 3600
rect 5150 3590 5300 3600
rect 6550 3590 6600 3600
rect 8300 3590 8400 3600
rect 8500 3590 8550 3600
rect 9250 3590 9400 3600
rect 9550 3590 9700 3600
rect 4000 3580 4050 3590
rect 4300 3580 4500 3590
rect 4650 3580 4750 3590
rect 4800 3580 4850 3590
rect 4950 3580 5050 3590
rect 5150 3580 5300 3590
rect 6550 3580 6600 3590
rect 8300 3580 8400 3590
rect 8500 3580 8550 3590
rect 9250 3580 9400 3590
rect 9550 3580 9700 3590
rect 4000 3570 4050 3580
rect 4300 3570 4500 3580
rect 4650 3570 4750 3580
rect 4800 3570 4850 3580
rect 4950 3570 5050 3580
rect 5150 3570 5300 3580
rect 6550 3570 6600 3580
rect 8300 3570 8400 3580
rect 8500 3570 8550 3580
rect 9250 3570 9400 3580
rect 9550 3570 9700 3580
rect 4000 3560 4050 3570
rect 4300 3560 4500 3570
rect 4650 3560 4750 3570
rect 4800 3560 4850 3570
rect 4950 3560 5050 3570
rect 5150 3560 5300 3570
rect 6550 3560 6600 3570
rect 8300 3560 8400 3570
rect 8500 3560 8550 3570
rect 9250 3560 9400 3570
rect 9550 3560 9700 3570
rect 4000 3550 4050 3560
rect 4300 3550 4500 3560
rect 4650 3550 4750 3560
rect 4800 3550 4850 3560
rect 4950 3550 5050 3560
rect 5150 3550 5300 3560
rect 6550 3550 6600 3560
rect 8300 3550 8400 3560
rect 8500 3550 8550 3560
rect 9250 3550 9400 3560
rect 9550 3550 9700 3560
rect 3350 3540 3400 3550
rect 4000 3540 4050 3550
rect 4250 3540 4300 3550
rect 4400 3540 4650 3550
rect 4800 3540 4850 3550
rect 4950 3540 5000 3550
rect 5150 3540 5300 3550
rect 6500 3540 6600 3550
rect 8350 3540 8400 3550
rect 8500 3540 8550 3550
rect 9150 3540 9250 3550
rect 9450 3540 9500 3550
rect 9550 3540 9650 3550
rect 3350 3530 3400 3540
rect 4000 3530 4050 3540
rect 4250 3530 4300 3540
rect 4400 3530 4650 3540
rect 4800 3530 4850 3540
rect 4950 3530 5000 3540
rect 5150 3530 5300 3540
rect 6500 3530 6600 3540
rect 8350 3530 8400 3540
rect 8500 3530 8550 3540
rect 9150 3530 9250 3540
rect 9450 3530 9500 3540
rect 9550 3530 9650 3540
rect 3350 3520 3400 3530
rect 4000 3520 4050 3530
rect 4250 3520 4300 3530
rect 4400 3520 4650 3530
rect 4800 3520 4850 3530
rect 4950 3520 5000 3530
rect 5150 3520 5300 3530
rect 6500 3520 6600 3530
rect 8350 3520 8400 3530
rect 8500 3520 8550 3530
rect 9150 3520 9250 3530
rect 9450 3520 9500 3530
rect 9550 3520 9650 3530
rect 3350 3510 3400 3520
rect 4000 3510 4050 3520
rect 4250 3510 4300 3520
rect 4400 3510 4650 3520
rect 4800 3510 4850 3520
rect 4950 3510 5000 3520
rect 5150 3510 5300 3520
rect 6500 3510 6600 3520
rect 8350 3510 8400 3520
rect 8500 3510 8550 3520
rect 9150 3510 9250 3520
rect 9450 3510 9500 3520
rect 9550 3510 9650 3520
rect 3350 3500 3400 3510
rect 4000 3500 4050 3510
rect 4250 3500 4300 3510
rect 4400 3500 4650 3510
rect 4800 3500 4850 3510
rect 4950 3500 5000 3510
rect 5150 3500 5300 3510
rect 6500 3500 6600 3510
rect 8350 3500 8400 3510
rect 8500 3500 8550 3510
rect 9150 3500 9250 3510
rect 9450 3500 9500 3510
rect 9550 3500 9650 3510
rect 2400 3490 2700 3500
rect 4000 3490 4100 3500
rect 4200 3490 4250 3500
rect 4750 3490 4800 3500
rect 4900 3490 4950 3500
rect 5050 3490 5300 3500
rect 6500 3490 6600 3500
rect 6800 3490 6850 3500
rect 9100 3490 9150 3500
rect 9350 3490 9550 3500
rect 9600 3490 9650 3500
rect 2400 3480 2700 3490
rect 4000 3480 4100 3490
rect 4200 3480 4250 3490
rect 4750 3480 4800 3490
rect 4900 3480 4950 3490
rect 5050 3480 5300 3490
rect 6500 3480 6600 3490
rect 6800 3480 6850 3490
rect 9100 3480 9150 3490
rect 9350 3480 9550 3490
rect 9600 3480 9650 3490
rect 2400 3470 2700 3480
rect 4000 3470 4100 3480
rect 4200 3470 4250 3480
rect 4750 3470 4800 3480
rect 4900 3470 4950 3480
rect 5050 3470 5300 3480
rect 6500 3470 6600 3480
rect 6800 3470 6850 3480
rect 9100 3470 9150 3480
rect 9350 3470 9550 3480
rect 9600 3470 9650 3480
rect 2400 3460 2700 3470
rect 4000 3460 4100 3470
rect 4200 3460 4250 3470
rect 4750 3460 4800 3470
rect 4900 3460 4950 3470
rect 5050 3460 5300 3470
rect 6500 3460 6600 3470
rect 6800 3460 6850 3470
rect 9100 3460 9150 3470
rect 9350 3460 9550 3470
rect 9600 3460 9650 3470
rect 2400 3450 2700 3460
rect 4000 3450 4100 3460
rect 4200 3450 4250 3460
rect 4750 3450 4800 3460
rect 4900 3450 4950 3460
rect 5050 3450 5300 3460
rect 6500 3450 6600 3460
rect 6800 3450 6850 3460
rect 9100 3450 9150 3460
rect 9350 3450 9550 3460
rect 9600 3450 9650 3460
rect 2300 3440 2350 3450
rect 2850 3440 2900 3450
rect 4050 3440 4250 3450
rect 4800 3440 4850 3450
rect 5100 3440 5300 3450
rect 6450 3440 6550 3450
rect 6750 3440 6800 3450
rect 9050 3440 9100 3450
rect 9250 3440 9300 3450
rect 9400 3440 9450 3450
rect 2300 3430 2350 3440
rect 2850 3430 2900 3440
rect 4050 3430 4250 3440
rect 4800 3430 4850 3440
rect 5100 3430 5300 3440
rect 6450 3430 6550 3440
rect 6750 3430 6800 3440
rect 9050 3430 9100 3440
rect 9250 3430 9300 3440
rect 9400 3430 9450 3440
rect 2300 3420 2350 3430
rect 2850 3420 2900 3430
rect 4050 3420 4250 3430
rect 4800 3420 4850 3430
rect 5100 3420 5300 3430
rect 6450 3420 6550 3430
rect 6750 3420 6800 3430
rect 9050 3420 9100 3430
rect 9250 3420 9300 3430
rect 9400 3420 9450 3430
rect 2300 3410 2350 3420
rect 2850 3410 2900 3420
rect 4050 3410 4250 3420
rect 4800 3410 4850 3420
rect 5100 3410 5300 3420
rect 6450 3410 6550 3420
rect 6750 3410 6800 3420
rect 9050 3410 9100 3420
rect 9250 3410 9300 3420
rect 9400 3410 9450 3420
rect 2300 3400 2350 3410
rect 2850 3400 2900 3410
rect 4050 3400 4250 3410
rect 4800 3400 4850 3410
rect 5100 3400 5300 3410
rect 6450 3400 6550 3410
rect 6750 3400 6800 3410
rect 9050 3400 9100 3410
rect 9250 3400 9300 3410
rect 9400 3400 9450 3410
rect 2200 3390 2250 3400
rect 2950 3390 3000 3400
rect 4100 3390 4200 3400
rect 4400 3390 4450 3400
rect 5000 3390 5050 3400
rect 5200 3390 5250 3400
rect 6400 3390 6550 3400
rect 9000 3390 9050 3400
rect 9150 3390 9200 3400
rect 9400 3390 9450 3400
rect 9650 3390 9800 3400
rect 2200 3380 2250 3390
rect 2950 3380 3000 3390
rect 4100 3380 4200 3390
rect 4400 3380 4450 3390
rect 5000 3380 5050 3390
rect 5200 3380 5250 3390
rect 6400 3380 6550 3390
rect 9000 3380 9050 3390
rect 9150 3380 9200 3390
rect 9400 3380 9450 3390
rect 9650 3380 9800 3390
rect 2200 3370 2250 3380
rect 2950 3370 3000 3380
rect 4100 3370 4200 3380
rect 4400 3370 4450 3380
rect 5000 3370 5050 3380
rect 5200 3370 5250 3380
rect 6400 3370 6550 3380
rect 9000 3370 9050 3380
rect 9150 3370 9200 3380
rect 9400 3370 9450 3380
rect 9650 3370 9800 3380
rect 2200 3360 2250 3370
rect 2950 3360 3000 3370
rect 4100 3360 4200 3370
rect 4400 3360 4450 3370
rect 5000 3360 5050 3370
rect 5200 3360 5250 3370
rect 6400 3360 6550 3370
rect 9000 3360 9050 3370
rect 9150 3360 9200 3370
rect 9400 3360 9450 3370
rect 9650 3360 9800 3370
rect 2200 3350 2250 3360
rect 2950 3350 3000 3360
rect 4100 3350 4200 3360
rect 4400 3350 4450 3360
rect 5000 3350 5050 3360
rect 5200 3350 5250 3360
rect 6400 3350 6550 3360
rect 9000 3350 9050 3360
rect 9150 3350 9200 3360
rect 9400 3350 9450 3360
rect 9650 3350 9800 3360
rect 2150 3340 2200 3350
rect 3050 3340 3100 3350
rect 4350 3340 4550 3350
rect 4900 3340 4950 3350
rect 5000 3340 5050 3350
rect 5200 3340 5250 3350
rect 6350 3340 6550 3350
rect 8500 3340 8550 3350
rect 8950 3340 9050 3350
rect 9300 3340 9400 3350
rect 9600 3340 9650 3350
rect 9750 3340 9800 3350
rect 2150 3330 2200 3340
rect 3050 3330 3100 3340
rect 4350 3330 4550 3340
rect 4900 3330 4950 3340
rect 5000 3330 5050 3340
rect 5200 3330 5250 3340
rect 6350 3330 6550 3340
rect 8500 3330 8550 3340
rect 8950 3330 9050 3340
rect 9300 3330 9400 3340
rect 9600 3330 9650 3340
rect 9750 3330 9800 3340
rect 2150 3320 2200 3330
rect 3050 3320 3100 3330
rect 4350 3320 4550 3330
rect 4900 3320 4950 3330
rect 5000 3320 5050 3330
rect 5200 3320 5250 3330
rect 6350 3320 6550 3330
rect 8500 3320 8550 3330
rect 8950 3320 9050 3330
rect 9300 3320 9400 3330
rect 9600 3320 9650 3330
rect 9750 3320 9800 3330
rect 2150 3310 2200 3320
rect 3050 3310 3100 3320
rect 4350 3310 4550 3320
rect 4900 3310 4950 3320
rect 5000 3310 5050 3320
rect 5200 3310 5250 3320
rect 6350 3310 6550 3320
rect 8500 3310 8550 3320
rect 8950 3310 9050 3320
rect 9300 3310 9400 3320
rect 9600 3310 9650 3320
rect 9750 3310 9800 3320
rect 2150 3300 2200 3310
rect 3050 3300 3100 3310
rect 4350 3300 4550 3310
rect 4900 3300 4950 3310
rect 5000 3300 5050 3310
rect 5200 3300 5250 3310
rect 6350 3300 6550 3310
rect 8500 3300 8550 3310
rect 8950 3300 9050 3310
rect 9300 3300 9400 3310
rect 9600 3300 9650 3310
rect 9750 3300 9800 3310
rect 4800 3290 4950 3300
rect 5000 3290 5050 3300
rect 5200 3290 5250 3300
rect 6300 3290 6550 3300
rect 8450 3290 8500 3300
rect 8850 3290 9050 3300
rect 9100 3290 9150 3300
rect 9300 3290 9350 3300
rect 9450 3290 9600 3300
rect 9700 3290 9750 3300
rect 9950 3290 9990 3300
rect 4800 3280 4950 3290
rect 5000 3280 5050 3290
rect 5200 3280 5250 3290
rect 6300 3280 6550 3290
rect 8450 3280 8500 3290
rect 8850 3280 9050 3290
rect 9100 3280 9150 3290
rect 9300 3280 9350 3290
rect 9450 3280 9600 3290
rect 9700 3280 9750 3290
rect 9950 3280 9990 3290
rect 4800 3270 4950 3280
rect 5000 3270 5050 3280
rect 5200 3270 5250 3280
rect 6300 3270 6550 3280
rect 8450 3270 8500 3280
rect 8850 3270 9050 3280
rect 9100 3270 9150 3280
rect 9300 3270 9350 3280
rect 9450 3270 9600 3280
rect 9700 3270 9750 3280
rect 9950 3270 9990 3280
rect 4800 3260 4950 3270
rect 5000 3260 5050 3270
rect 5200 3260 5250 3270
rect 6300 3260 6550 3270
rect 8450 3260 8500 3270
rect 8850 3260 9050 3270
rect 9100 3260 9150 3270
rect 9300 3260 9350 3270
rect 9450 3260 9600 3270
rect 9700 3260 9750 3270
rect 9950 3260 9990 3270
rect 4800 3250 4950 3260
rect 5000 3250 5050 3260
rect 5200 3250 5250 3260
rect 6300 3250 6550 3260
rect 8450 3250 8500 3260
rect 8850 3250 9050 3260
rect 9100 3250 9150 3260
rect 9300 3250 9350 3260
rect 9450 3250 9600 3260
rect 9700 3250 9750 3260
rect 9950 3250 9990 3260
rect 2100 3240 2150 3250
rect 3100 3240 3150 3250
rect 4750 3240 4900 3250
rect 5200 3240 5250 3250
rect 6300 3240 6400 3250
rect 8950 3240 9050 3250
rect 9150 3240 9300 3250
rect 9650 3240 9700 3250
rect 9900 3240 9990 3250
rect 2100 3230 2150 3240
rect 3100 3230 3150 3240
rect 4750 3230 4900 3240
rect 5200 3230 5250 3240
rect 6300 3230 6400 3240
rect 8950 3230 9050 3240
rect 9150 3230 9300 3240
rect 9650 3230 9700 3240
rect 9900 3230 9990 3240
rect 2100 3220 2150 3230
rect 3100 3220 3150 3230
rect 4750 3220 4900 3230
rect 5200 3220 5250 3230
rect 6300 3220 6400 3230
rect 8950 3220 9050 3230
rect 9150 3220 9300 3230
rect 9650 3220 9700 3230
rect 9900 3220 9990 3230
rect 2100 3210 2150 3220
rect 3100 3210 3150 3220
rect 4750 3210 4900 3220
rect 5200 3210 5250 3220
rect 6300 3210 6400 3220
rect 8950 3210 9050 3220
rect 9150 3210 9300 3220
rect 9650 3210 9700 3220
rect 9900 3210 9990 3220
rect 2100 3200 2150 3210
rect 3100 3200 3150 3210
rect 4750 3200 4900 3210
rect 5200 3200 5250 3210
rect 6300 3200 6400 3210
rect 8950 3200 9050 3210
rect 9150 3200 9300 3210
rect 9650 3200 9700 3210
rect 9900 3200 9990 3210
rect 2100 3190 2150 3200
rect 4650 3190 4850 3200
rect 4950 3190 5000 3200
rect 5200 3190 5250 3200
rect 8400 3190 8450 3200
rect 8850 3190 9000 3200
rect 9600 3190 9650 3200
rect 9850 3190 9990 3200
rect 2100 3180 2150 3190
rect 4650 3180 4850 3190
rect 4950 3180 5000 3190
rect 5200 3180 5250 3190
rect 8400 3180 8450 3190
rect 8850 3180 9000 3190
rect 9600 3180 9650 3190
rect 9850 3180 9990 3190
rect 2100 3170 2150 3180
rect 4650 3170 4850 3180
rect 4950 3170 5000 3180
rect 5200 3170 5250 3180
rect 8400 3170 8450 3180
rect 8850 3170 9000 3180
rect 9600 3170 9650 3180
rect 9850 3170 9990 3180
rect 2100 3160 2150 3170
rect 4650 3160 4850 3170
rect 4950 3160 5000 3170
rect 5200 3160 5250 3170
rect 8400 3160 8450 3170
rect 8850 3160 9000 3170
rect 9600 3160 9650 3170
rect 9850 3160 9990 3170
rect 2100 3150 2150 3160
rect 4650 3150 4850 3160
rect 4950 3150 5000 3160
rect 5200 3150 5250 3160
rect 8400 3150 8450 3160
rect 8850 3150 9000 3160
rect 9600 3150 9650 3160
rect 9850 3150 9990 3160
rect 4250 3140 4300 3150
rect 4350 3140 4450 3150
rect 4650 3140 4750 3150
rect 4950 3140 5000 3150
rect 5200 3140 5250 3150
rect 8400 3140 8450 3150
rect 8800 3140 8900 3150
rect 9550 3140 9600 3150
rect 9800 3140 9850 3150
rect 4250 3130 4300 3140
rect 4350 3130 4450 3140
rect 4650 3130 4750 3140
rect 4950 3130 5000 3140
rect 5200 3130 5250 3140
rect 8400 3130 8450 3140
rect 8800 3130 8900 3140
rect 9550 3130 9600 3140
rect 9800 3130 9850 3140
rect 4250 3120 4300 3130
rect 4350 3120 4450 3130
rect 4650 3120 4750 3130
rect 4950 3120 5000 3130
rect 5200 3120 5250 3130
rect 8400 3120 8450 3130
rect 8800 3120 8900 3130
rect 9550 3120 9600 3130
rect 9800 3120 9850 3130
rect 4250 3110 4300 3120
rect 4350 3110 4450 3120
rect 4650 3110 4750 3120
rect 4950 3110 5000 3120
rect 5200 3110 5250 3120
rect 8400 3110 8450 3120
rect 8800 3110 8900 3120
rect 9550 3110 9600 3120
rect 9800 3110 9850 3120
rect 4250 3100 4300 3110
rect 4350 3100 4450 3110
rect 4650 3100 4750 3110
rect 4950 3100 5000 3110
rect 5200 3100 5250 3110
rect 8400 3100 8450 3110
rect 8800 3100 8900 3110
rect 9550 3100 9600 3110
rect 9800 3100 9850 3110
rect 2050 3090 2100 3100
rect 3900 3090 4000 3100
rect 4300 3090 4500 3100
rect 4950 3090 5000 3100
rect 5150 3090 5200 3100
rect 8400 3090 8450 3100
rect 8800 3090 9000 3100
rect 9500 3090 9550 3100
rect 9750 3090 9800 3100
rect 9900 3090 9990 3100
rect 2050 3080 2100 3090
rect 3900 3080 4000 3090
rect 4300 3080 4500 3090
rect 4950 3080 5000 3090
rect 5150 3080 5200 3090
rect 8400 3080 8450 3090
rect 8800 3080 9000 3090
rect 9500 3080 9550 3090
rect 9750 3080 9800 3090
rect 9900 3080 9990 3090
rect 2050 3070 2100 3080
rect 3900 3070 4000 3080
rect 4300 3070 4500 3080
rect 4950 3070 5000 3080
rect 5150 3070 5200 3080
rect 8400 3070 8450 3080
rect 8800 3070 9000 3080
rect 9500 3070 9550 3080
rect 9750 3070 9800 3080
rect 9900 3070 9990 3080
rect 2050 3060 2100 3070
rect 3900 3060 4000 3070
rect 4300 3060 4500 3070
rect 4950 3060 5000 3070
rect 5150 3060 5200 3070
rect 8400 3060 8450 3070
rect 8800 3060 9000 3070
rect 9500 3060 9550 3070
rect 9750 3060 9800 3070
rect 9900 3060 9990 3070
rect 2050 3050 2100 3060
rect 3900 3050 4000 3060
rect 4300 3050 4500 3060
rect 4950 3050 5000 3060
rect 5150 3050 5200 3060
rect 8400 3050 8450 3060
rect 8800 3050 9000 3060
rect 9500 3050 9550 3060
rect 9750 3050 9800 3060
rect 9900 3050 9990 3060
rect 2050 3040 2100 3050
rect 3100 3040 3150 3050
rect 3900 3040 3950 3050
rect 4000 3040 4050 3050
rect 4350 3040 4450 3050
rect 4900 3040 5200 3050
rect 8350 3040 8450 3050
rect 8600 3040 8900 3050
rect 9750 3040 9800 3050
rect 9900 3040 9950 3050
rect 2050 3030 2100 3040
rect 3100 3030 3150 3040
rect 3900 3030 3950 3040
rect 4000 3030 4050 3040
rect 4350 3030 4450 3040
rect 4900 3030 5200 3040
rect 8350 3030 8450 3040
rect 8600 3030 8900 3040
rect 9750 3030 9800 3040
rect 9900 3030 9950 3040
rect 2050 3020 2100 3030
rect 3100 3020 3150 3030
rect 3900 3020 3950 3030
rect 4000 3020 4050 3030
rect 4350 3020 4450 3030
rect 4900 3020 5200 3030
rect 8350 3020 8450 3030
rect 8600 3020 8900 3030
rect 9750 3020 9800 3030
rect 9900 3020 9950 3030
rect 2050 3010 2100 3020
rect 3100 3010 3150 3020
rect 3900 3010 3950 3020
rect 4000 3010 4050 3020
rect 4350 3010 4450 3020
rect 4900 3010 5200 3020
rect 8350 3010 8450 3020
rect 8600 3010 8900 3020
rect 9750 3010 9800 3020
rect 9900 3010 9950 3020
rect 2050 3000 2100 3010
rect 3100 3000 3150 3010
rect 3900 3000 3950 3010
rect 4000 3000 4050 3010
rect 4350 3000 4450 3010
rect 4900 3000 5200 3010
rect 8350 3000 8450 3010
rect 8600 3000 8900 3010
rect 9750 3000 9800 3010
rect 9900 3000 9950 3010
rect 2050 2990 2100 3000
rect 3100 2990 3150 3000
rect 4400 2990 4450 3000
rect 4950 2990 5150 3000
rect 8300 2990 8350 3000
rect 8550 2990 8700 3000
rect 9450 2990 9500 3000
rect 9750 2990 9950 3000
rect 2050 2980 2100 2990
rect 3100 2980 3150 2990
rect 4400 2980 4450 2990
rect 4950 2980 5150 2990
rect 8300 2980 8350 2990
rect 8550 2980 8700 2990
rect 9450 2980 9500 2990
rect 9750 2980 9950 2990
rect 2050 2970 2100 2980
rect 3100 2970 3150 2980
rect 4400 2970 4450 2980
rect 4950 2970 5150 2980
rect 8300 2970 8350 2980
rect 8550 2970 8700 2980
rect 9450 2970 9500 2980
rect 9750 2970 9950 2980
rect 2050 2960 2100 2970
rect 3100 2960 3150 2970
rect 4400 2960 4450 2970
rect 4950 2960 5150 2970
rect 8300 2960 8350 2970
rect 8550 2960 8700 2970
rect 9450 2960 9500 2970
rect 9750 2960 9950 2970
rect 2050 2950 2100 2960
rect 3100 2950 3150 2960
rect 4400 2950 4450 2960
rect 4950 2950 5150 2960
rect 8300 2950 8350 2960
rect 8550 2950 8700 2960
rect 9450 2950 9500 2960
rect 9750 2950 9950 2960
rect 2050 2940 2100 2950
rect 3100 2940 3150 2950
rect 4150 2940 4200 2950
rect 5000 2940 5100 2950
rect 8500 2940 8650 2950
rect 9400 2940 9450 2950
rect 9650 2940 9750 2950
rect 9900 2940 9990 2950
rect 2050 2930 2100 2940
rect 3100 2930 3150 2940
rect 4150 2930 4200 2940
rect 5000 2930 5100 2940
rect 8500 2930 8650 2940
rect 9400 2930 9450 2940
rect 9650 2930 9750 2940
rect 9900 2930 9990 2940
rect 2050 2920 2100 2930
rect 3100 2920 3150 2930
rect 4150 2920 4200 2930
rect 5000 2920 5100 2930
rect 8500 2920 8650 2930
rect 9400 2920 9450 2930
rect 9650 2920 9750 2930
rect 9900 2920 9990 2930
rect 2050 2910 2100 2920
rect 3100 2910 3150 2920
rect 4150 2910 4200 2920
rect 5000 2910 5100 2920
rect 8500 2910 8650 2920
rect 9400 2910 9450 2920
rect 9650 2910 9750 2920
rect 9900 2910 9990 2920
rect 2050 2900 2100 2910
rect 3100 2900 3150 2910
rect 4150 2900 4200 2910
rect 5000 2900 5100 2910
rect 8500 2900 8650 2910
rect 9400 2900 9450 2910
rect 9650 2900 9750 2910
rect 9900 2900 9990 2910
rect 3100 2890 3150 2900
rect 4200 2890 4250 2900
rect 8250 2890 8300 2900
rect 8500 2890 8600 2900
rect 9650 2890 9750 2900
rect 9900 2890 9990 2900
rect 3100 2880 3150 2890
rect 4200 2880 4250 2890
rect 8250 2880 8300 2890
rect 8500 2880 8600 2890
rect 9650 2880 9750 2890
rect 9900 2880 9990 2890
rect 3100 2870 3150 2880
rect 4200 2870 4250 2880
rect 8250 2870 8300 2880
rect 8500 2870 8600 2880
rect 9650 2870 9750 2880
rect 9900 2870 9990 2880
rect 3100 2860 3150 2870
rect 4200 2860 4250 2870
rect 8250 2860 8300 2870
rect 8500 2860 8600 2870
rect 9650 2860 9750 2870
rect 9900 2860 9990 2870
rect 3100 2850 3150 2860
rect 4200 2850 4250 2860
rect 8250 2850 8300 2860
rect 8500 2850 8600 2860
rect 9650 2850 9750 2860
rect 9900 2850 9990 2860
rect 3050 2840 3100 2850
rect 7200 2840 7250 2850
rect 7500 2840 7550 2850
rect 8200 2840 8250 2850
rect 8500 2840 8600 2850
rect 9100 2840 9150 2850
rect 9400 2840 9450 2850
rect 9600 2840 9700 2850
rect 9900 2840 9990 2850
rect 3050 2830 3100 2840
rect 7200 2830 7250 2840
rect 7500 2830 7550 2840
rect 8200 2830 8250 2840
rect 8500 2830 8600 2840
rect 9100 2830 9150 2840
rect 9400 2830 9450 2840
rect 9600 2830 9700 2840
rect 9900 2830 9990 2840
rect 3050 2820 3100 2830
rect 7200 2820 7250 2830
rect 7500 2820 7550 2830
rect 8200 2820 8250 2830
rect 8500 2820 8600 2830
rect 9100 2820 9150 2830
rect 9400 2820 9450 2830
rect 9600 2820 9700 2830
rect 9900 2820 9990 2830
rect 3050 2810 3100 2820
rect 7200 2810 7250 2820
rect 7500 2810 7550 2820
rect 8200 2810 8250 2820
rect 8500 2810 8600 2820
rect 9100 2810 9150 2820
rect 9400 2810 9450 2820
rect 9600 2810 9700 2820
rect 9900 2810 9990 2820
rect 3050 2800 3100 2810
rect 7200 2800 7250 2810
rect 7500 2800 7550 2810
rect 8200 2800 8250 2810
rect 8500 2800 8600 2810
rect 9100 2800 9150 2810
rect 9400 2800 9450 2810
rect 9600 2800 9700 2810
rect 9900 2800 9990 2810
rect 2050 2790 2100 2800
rect 2200 2790 2450 2800
rect 2800 2790 3100 2800
rect 3950 2790 4000 2800
rect 7550 2790 7600 2800
rect 8500 2790 8600 2800
rect 9300 2790 9400 2800
rect 9450 2790 9650 2800
rect 9700 2790 9750 2800
rect 9900 2790 9950 2800
rect 2050 2780 2100 2790
rect 2200 2780 2450 2790
rect 2800 2780 3100 2790
rect 3950 2780 4000 2790
rect 7550 2780 7600 2790
rect 8500 2780 8600 2790
rect 9300 2780 9400 2790
rect 9450 2780 9650 2790
rect 9700 2780 9750 2790
rect 9900 2780 9950 2790
rect 2050 2770 2100 2780
rect 2200 2770 2450 2780
rect 2800 2770 3100 2780
rect 3950 2770 4000 2780
rect 7550 2770 7600 2780
rect 8500 2770 8600 2780
rect 9300 2770 9400 2780
rect 9450 2770 9650 2780
rect 9700 2770 9750 2780
rect 9900 2770 9950 2780
rect 2050 2760 2100 2770
rect 2200 2760 2450 2770
rect 2800 2760 3100 2770
rect 3950 2760 4000 2770
rect 7550 2760 7600 2770
rect 8500 2760 8600 2770
rect 9300 2760 9400 2770
rect 9450 2760 9650 2770
rect 9700 2760 9750 2770
rect 9900 2760 9950 2770
rect 2050 2750 2100 2760
rect 2200 2750 2450 2760
rect 2800 2750 3100 2760
rect 3950 2750 4000 2760
rect 7550 2750 7600 2760
rect 8500 2750 8600 2760
rect 9300 2750 9400 2760
rect 9450 2750 9650 2760
rect 9700 2750 9750 2760
rect 9900 2750 9950 2760
rect 2050 2740 2100 2750
rect 2250 2740 2450 2750
rect 2750 2740 3000 2750
rect 3100 2740 3150 2750
rect 7050 2740 7100 2750
rect 7600 2740 7650 2750
rect 8550 2740 8650 2750
rect 9300 2740 9450 2750
rect 9500 2740 9600 2750
rect 9700 2740 9750 2750
rect 2050 2730 2100 2740
rect 2250 2730 2450 2740
rect 2750 2730 3000 2740
rect 3100 2730 3150 2740
rect 7050 2730 7100 2740
rect 7600 2730 7650 2740
rect 8550 2730 8650 2740
rect 9300 2730 9450 2740
rect 9500 2730 9600 2740
rect 9700 2730 9750 2740
rect 2050 2720 2100 2730
rect 2250 2720 2450 2730
rect 2750 2720 3000 2730
rect 3100 2720 3150 2730
rect 7050 2720 7100 2730
rect 7600 2720 7650 2730
rect 8550 2720 8650 2730
rect 9300 2720 9450 2730
rect 9500 2720 9600 2730
rect 9700 2720 9750 2730
rect 2050 2710 2100 2720
rect 2250 2710 2450 2720
rect 2750 2710 3000 2720
rect 3100 2710 3150 2720
rect 7050 2710 7100 2720
rect 7600 2710 7650 2720
rect 8550 2710 8650 2720
rect 9300 2710 9450 2720
rect 9500 2710 9600 2720
rect 9700 2710 9750 2720
rect 2050 2700 2100 2710
rect 2250 2700 2450 2710
rect 2750 2700 3000 2710
rect 3100 2700 3150 2710
rect 7050 2700 7100 2710
rect 7600 2700 7650 2710
rect 8550 2700 8650 2710
rect 9300 2700 9450 2710
rect 9500 2700 9600 2710
rect 9700 2700 9750 2710
rect 2000 2690 2050 2700
rect 2100 2690 2200 2700
rect 2450 2690 2500 2700
rect 2750 2690 2800 2700
rect 3000 2690 3100 2700
rect 3900 2690 3950 2700
rect 4200 2690 4250 2700
rect 6950 2690 7000 2700
rect 7650 2690 7700 2700
rect 8550 2690 8650 2700
rect 9250 2690 9300 2700
rect 9600 2690 9750 2700
rect 9900 2690 9950 2700
rect 2000 2680 2050 2690
rect 2100 2680 2200 2690
rect 2450 2680 2500 2690
rect 2750 2680 2800 2690
rect 3000 2680 3100 2690
rect 3900 2680 3950 2690
rect 4200 2680 4250 2690
rect 6950 2680 7000 2690
rect 7650 2680 7700 2690
rect 8550 2680 8650 2690
rect 9250 2680 9300 2690
rect 9600 2680 9750 2690
rect 9900 2680 9950 2690
rect 2000 2670 2050 2680
rect 2100 2670 2200 2680
rect 2450 2670 2500 2680
rect 2750 2670 2800 2680
rect 3000 2670 3100 2680
rect 3900 2670 3950 2680
rect 4200 2670 4250 2680
rect 6950 2670 7000 2680
rect 7650 2670 7700 2680
rect 8550 2670 8650 2680
rect 9250 2670 9300 2680
rect 9600 2670 9750 2680
rect 9900 2670 9950 2680
rect 2000 2660 2050 2670
rect 2100 2660 2200 2670
rect 2450 2660 2500 2670
rect 2750 2660 2800 2670
rect 3000 2660 3100 2670
rect 3900 2660 3950 2670
rect 4200 2660 4250 2670
rect 6950 2660 7000 2670
rect 7650 2660 7700 2670
rect 8550 2660 8650 2670
rect 9250 2660 9300 2670
rect 9600 2660 9750 2670
rect 9900 2660 9950 2670
rect 2000 2650 2050 2660
rect 2100 2650 2200 2660
rect 2450 2650 2500 2660
rect 2750 2650 2800 2660
rect 3000 2650 3100 2660
rect 3900 2650 3950 2660
rect 4200 2650 4250 2660
rect 6950 2650 7000 2660
rect 7650 2650 7700 2660
rect 8550 2650 8650 2660
rect 9250 2650 9300 2660
rect 9600 2650 9750 2660
rect 9900 2650 9950 2660
rect 2000 2640 2050 2650
rect 2450 2640 2500 2650
rect 2700 2640 2750 2650
rect 6900 2640 6950 2650
rect 7150 2640 7250 2650
rect 8050 2640 8100 2650
rect 8400 2640 8700 2650
rect 8750 2640 8850 2650
rect 9200 2640 9250 2650
rect 9700 2640 9850 2650
rect 2000 2630 2050 2640
rect 2450 2630 2500 2640
rect 2700 2630 2750 2640
rect 6900 2630 6950 2640
rect 7150 2630 7250 2640
rect 8050 2630 8100 2640
rect 8400 2630 8700 2640
rect 8750 2630 8850 2640
rect 9200 2630 9250 2640
rect 9700 2630 9850 2640
rect 2000 2620 2050 2630
rect 2450 2620 2500 2630
rect 2700 2620 2750 2630
rect 6900 2620 6950 2630
rect 7150 2620 7250 2630
rect 8050 2620 8100 2630
rect 8400 2620 8700 2630
rect 8750 2620 8850 2630
rect 9200 2620 9250 2630
rect 9700 2620 9850 2630
rect 2000 2610 2050 2620
rect 2450 2610 2500 2620
rect 2700 2610 2750 2620
rect 6900 2610 6950 2620
rect 7150 2610 7250 2620
rect 8050 2610 8100 2620
rect 8400 2610 8700 2620
rect 8750 2610 8850 2620
rect 9200 2610 9250 2620
rect 9700 2610 9850 2620
rect 2000 2600 2050 2610
rect 2450 2600 2500 2610
rect 2700 2600 2750 2610
rect 6900 2600 6950 2610
rect 7150 2600 7250 2610
rect 8050 2600 8100 2610
rect 8400 2600 8700 2610
rect 8750 2600 8850 2610
rect 9200 2600 9250 2610
rect 9700 2600 9850 2610
rect 2750 2590 2800 2600
rect 3950 2590 4000 2600
rect 4050 2590 4200 2600
rect 6850 2590 6900 2600
rect 7100 2590 7200 2600
rect 8000 2590 8050 2600
rect 8400 2590 8850 2600
rect 9400 2590 9600 2600
rect 9800 2590 9850 2600
rect 2750 2580 2800 2590
rect 3950 2580 4000 2590
rect 4050 2580 4200 2590
rect 6850 2580 6900 2590
rect 7100 2580 7200 2590
rect 8000 2580 8050 2590
rect 8400 2580 8850 2590
rect 9400 2580 9600 2590
rect 9800 2580 9850 2590
rect 2750 2570 2800 2580
rect 3950 2570 4000 2580
rect 4050 2570 4200 2580
rect 6850 2570 6900 2580
rect 7100 2570 7200 2580
rect 8000 2570 8050 2580
rect 8400 2570 8850 2580
rect 9400 2570 9600 2580
rect 9800 2570 9850 2580
rect 2750 2560 2800 2570
rect 3950 2560 4000 2570
rect 4050 2560 4200 2570
rect 6850 2560 6900 2570
rect 7100 2560 7200 2570
rect 8000 2560 8050 2570
rect 8400 2560 8850 2570
rect 9400 2560 9600 2570
rect 9800 2560 9850 2570
rect 2750 2550 2800 2560
rect 3950 2550 4000 2560
rect 4050 2550 4200 2560
rect 6850 2550 6900 2560
rect 7100 2550 7200 2560
rect 8000 2550 8050 2560
rect 8400 2550 8850 2560
rect 9400 2550 9600 2560
rect 9800 2550 9850 2560
rect 2400 2540 2450 2550
rect 2800 2540 3100 2550
rect 6800 2540 6850 2550
rect 7150 2540 7250 2550
rect 7300 2540 7350 2550
rect 7750 2540 7800 2550
rect 8400 2540 8850 2550
rect 9150 2540 9200 2550
rect 9300 2540 9350 2550
rect 9600 2540 9700 2550
rect 9900 2540 9950 2550
rect 2400 2530 2450 2540
rect 2800 2530 3100 2540
rect 6800 2530 6850 2540
rect 7150 2530 7250 2540
rect 7300 2530 7350 2540
rect 7750 2530 7800 2540
rect 8400 2530 8850 2540
rect 9150 2530 9200 2540
rect 9300 2530 9350 2540
rect 9600 2530 9700 2540
rect 9900 2530 9950 2540
rect 2400 2520 2450 2530
rect 2800 2520 3100 2530
rect 6800 2520 6850 2530
rect 7150 2520 7250 2530
rect 7300 2520 7350 2530
rect 7750 2520 7800 2530
rect 8400 2520 8850 2530
rect 9150 2520 9200 2530
rect 9300 2520 9350 2530
rect 9600 2520 9700 2530
rect 9900 2520 9950 2530
rect 2400 2510 2450 2520
rect 2800 2510 3100 2520
rect 6800 2510 6850 2520
rect 7150 2510 7250 2520
rect 7300 2510 7350 2520
rect 7750 2510 7800 2520
rect 8400 2510 8850 2520
rect 9150 2510 9200 2520
rect 9300 2510 9350 2520
rect 9600 2510 9700 2520
rect 9900 2510 9950 2520
rect 2400 2500 2450 2510
rect 2800 2500 3100 2510
rect 6800 2500 6850 2510
rect 7150 2500 7250 2510
rect 7300 2500 7350 2510
rect 7750 2500 7800 2510
rect 8400 2500 8850 2510
rect 9150 2500 9200 2510
rect 9300 2500 9350 2510
rect 9600 2500 9700 2510
rect 9900 2500 9950 2510
rect 1950 2490 2000 2500
rect 2050 2490 2350 2500
rect 3000 2490 3200 2500
rect 6800 2490 6900 2500
rect 7200 2490 7250 2500
rect 7350 2490 7400 2500
rect 7800 2490 7900 2500
rect 8400 2490 8950 2500
rect 9700 2490 9750 2500
rect 1950 2480 2000 2490
rect 2050 2480 2350 2490
rect 3000 2480 3200 2490
rect 6800 2480 6900 2490
rect 7200 2480 7250 2490
rect 7350 2480 7400 2490
rect 7800 2480 7900 2490
rect 8400 2480 8950 2490
rect 9700 2480 9750 2490
rect 1950 2470 2000 2480
rect 2050 2470 2350 2480
rect 3000 2470 3200 2480
rect 6800 2470 6900 2480
rect 7200 2470 7250 2480
rect 7350 2470 7400 2480
rect 7800 2470 7900 2480
rect 8400 2470 8950 2480
rect 9700 2470 9750 2480
rect 1950 2460 2000 2470
rect 2050 2460 2350 2470
rect 3000 2460 3200 2470
rect 6800 2460 6900 2470
rect 7200 2460 7250 2470
rect 7350 2460 7400 2470
rect 7800 2460 7900 2470
rect 8400 2460 8950 2470
rect 9700 2460 9750 2470
rect 1950 2450 2000 2460
rect 2050 2450 2350 2460
rect 3000 2450 3200 2460
rect 6800 2450 6900 2460
rect 7200 2450 7250 2460
rect 7350 2450 7400 2460
rect 7800 2450 7900 2460
rect 8400 2450 8950 2460
rect 9700 2450 9750 2460
rect 2100 2440 2250 2450
rect 3200 2440 3250 2450
rect 6850 2440 6950 2450
rect 8400 2440 9250 2450
rect 9800 2440 9850 2450
rect 2100 2430 2250 2440
rect 3200 2430 3250 2440
rect 6850 2430 6950 2440
rect 8400 2430 9250 2440
rect 9800 2430 9850 2440
rect 2100 2420 2250 2430
rect 3200 2420 3250 2430
rect 6850 2420 6950 2430
rect 8400 2420 9250 2430
rect 9800 2420 9850 2430
rect 2100 2410 2250 2420
rect 3200 2410 3250 2420
rect 6850 2410 6950 2420
rect 8400 2410 9250 2420
rect 9800 2410 9850 2420
rect 2100 2400 2250 2410
rect 3200 2400 3250 2410
rect 6850 2400 6950 2410
rect 8400 2400 9250 2410
rect 9800 2400 9850 2410
rect 3200 2390 3250 2400
rect 6950 2390 7100 2400
rect 7350 2390 7400 2400
rect 7450 2390 7500 2400
rect 8350 2390 8400 2400
rect 8500 2390 9150 2400
rect 9200 2390 9250 2400
rect 9500 2390 9550 2400
rect 9800 2390 9850 2400
rect 3200 2380 3250 2390
rect 6950 2380 7100 2390
rect 7350 2380 7400 2390
rect 7450 2380 7500 2390
rect 8350 2380 8400 2390
rect 8500 2380 9150 2390
rect 9200 2380 9250 2390
rect 9500 2380 9550 2390
rect 9800 2380 9850 2390
rect 3200 2370 3250 2380
rect 6950 2370 7100 2380
rect 7350 2370 7400 2380
rect 7450 2370 7500 2380
rect 8350 2370 8400 2380
rect 8500 2370 9150 2380
rect 9200 2370 9250 2380
rect 9500 2370 9550 2380
rect 9800 2370 9850 2380
rect 3200 2360 3250 2370
rect 6950 2360 7100 2370
rect 7350 2360 7400 2370
rect 7450 2360 7500 2370
rect 8350 2360 8400 2370
rect 8500 2360 9150 2370
rect 9200 2360 9250 2370
rect 9500 2360 9550 2370
rect 9800 2360 9850 2370
rect 3200 2350 3250 2360
rect 6950 2350 7100 2360
rect 7350 2350 7400 2360
rect 7450 2350 7500 2360
rect 8350 2350 8400 2360
rect 8500 2350 9150 2360
rect 9200 2350 9250 2360
rect 9500 2350 9550 2360
rect 9800 2350 9850 2360
rect 1900 2340 1950 2350
rect 3200 2340 3250 2350
rect 7100 2340 7250 2350
rect 7450 2340 7500 2350
rect 7550 2340 7600 2350
rect 8350 2340 8400 2350
rect 8600 2340 8650 2350
rect 8750 2340 9150 2350
rect 9800 2340 9850 2350
rect 1900 2330 1950 2340
rect 3200 2330 3250 2340
rect 7100 2330 7250 2340
rect 7450 2330 7500 2340
rect 7550 2330 7600 2340
rect 8350 2330 8400 2340
rect 8600 2330 8650 2340
rect 8750 2330 9150 2340
rect 9800 2330 9850 2340
rect 1900 2320 1950 2330
rect 3200 2320 3250 2330
rect 7100 2320 7250 2330
rect 7450 2320 7500 2330
rect 7550 2320 7600 2330
rect 8350 2320 8400 2330
rect 8600 2320 8650 2330
rect 8750 2320 9150 2330
rect 9800 2320 9850 2330
rect 1900 2310 1950 2320
rect 3200 2310 3250 2320
rect 7100 2310 7250 2320
rect 7450 2310 7500 2320
rect 7550 2310 7600 2320
rect 8350 2310 8400 2320
rect 8600 2310 8650 2320
rect 8750 2310 9150 2320
rect 9800 2310 9850 2320
rect 1900 2300 1950 2310
rect 3200 2300 3250 2310
rect 7100 2300 7250 2310
rect 7450 2300 7500 2310
rect 7550 2300 7600 2310
rect 8350 2300 8400 2310
rect 8600 2300 8650 2310
rect 8750 2300 9150 2310
rect 9800 2300 9850 2310
rect 1900 2290 1950 2300
rect 7250 2290 7400 2300
rect 7450 2290 7500 2300
rect 7600 2290 7650 2300
rect 8650 2290 9100 2300
rect 9800 2290 9850 2300
rect 1900 2280 1950 2290
rect 7250 2280 7400 2290
rect 7450 2280 7500 2290
rect 7600 2280 7650 2290
rect 8650 2280 9100 2290
rect 9800 2280 9850 2290
rect 1900 2270 1950 2280
rect 7250 2270 7400 2280
rect 7450 2270 7500 2280
rect 7600 2270 7650 2280
rect 8650 2270 9100 2280
rect 9800 2270 9850 2280
rect 1900 2260 1950 2270
rect 7250 2260 7400 2270
rect 7450 2260 7500 2270
rect 7600 2260 7650 2270
rect 8650 2260 9100 2270
rect 9800 2260 9850 2270
rect 1900 2250 1950 2260
rect 7250 2250 7400 2260
rect 7450 2250 7500 2260
rect 7600 2250 7650 2260
rect 8650 2250 9100 2260
rect 9800 2250 9850 2260
rect 2500 2240 2750 2250
rect 7400 2240 7500 2250
rect 7650 2240 7700 2250
rect 8850 2240 9000 2250
rect 9250 2240 9300 2250
rect 9800 2240 9850 2250
rect 2500 2230 2750 2240
rect 7400 2230 7500 2240
rect 7650 2230 7700 2240
rect 8850 2230 9000 2240
rect 9250 2230 9300 2240
rect 9800 2230 9850 2240
rect 2500 2220 2750 2230
rect 7400 2220 7500 2230
rect 7650 2220 7700 2230
rect 8850 2220 9000 2230
rect 9250 2220 9300 2230
rect 9800 2220 9850 2230
rect 2500 2210 2750 2220
rect 7400 2210 7500 2220
rect 7650 2210 7700 2220
rect 8850 2210 9000 2220
rect 9250 2210 9300 2220
rect 9800 2210 9850 2220
rect 2500 2200 2750 2210
rect 7400 2200 7500 2210
rect 7650 2200 7700 2210
rect 8850 2200 9000 2210
rect 9250 2200 9300 2210
rect 9800 2200 9850 2210
rect 2250 2190 2300 2200
rect 2350 2190 2450 2200
rect 2800 2190 2850 2200
rect 6400 2190 6450 2200
rect 7750 2190 7800 2200
rect 9250 2190 9300 2200
rect 9350 2190 9450 2200
rect 9800 2190 9850 2200
rect 9950 2190 9990 2200
rect 2250 2180 2300 2190
rect 2350 2180 2450 2190
rect 2800 2180 2850 2190
rect 6400 2180 6450 2190
rect 7750 2180 7800 2190
rect 9250 2180 9300 2190
rect 9350 2180 9450 2190
rect 9800 2180 9850 2190
rect 9950 2180 9990 2190
rect 2250 2170 2300 2180
rect 2350 2170 2450 2180
rect 2800 2170 2850 2180
rect 6400 2170 6450 2180
rect 7750 2170 7800 2180
rect 9250 2170 9300 2180
rect 9350 2170 9450 2180
rect 9800 2170 9850 2180
rect 9950 2170 9990 2180
rect 2250 2160 2300 2170
rect 2350 2160 2450 2170
rect 2800 2160 2850 2170
rect 6400 2160 6450 2170
rect 7750 2160 7800 2170
rect 9250 2160 9300 2170
rect 9350 2160 9450 2170
rect 9800 2160 9850 2170
rect 9950 2160 9990 2170
rect 2250 2150 2300 2160
rect 2350 2150 2450 2160
rect 2800 2150 2850 2160
rect 6400 2150 6450 2160
rect 7750 2150 7800 2160
rect 9250 2150 9300 2160
rect 9350 2150 9450 2160
rect 9800 2150 9850 2160
rect 9950 2150 9990 2160
rect 1900 2140 1950 2150
rect 2200 2140 2300 2150
rect 2350 2140 2400 2150
rect 2700 2140 2850 2150
rect 3200 2140 3250 2150
rect 6400 2140 6450 2150
rect 7850 2140 7900 2150
rect 8350 2140 8400 2150
rect 9300 2140 9350 2150
rect 9450 2140 9500 2150
rect 9700 2140 9800 2150
rect 1900 2130 1950 2140
rect 2200 2130 2300 2140
rect 2350 2130 2400 2140
rect 2700 2130 2850 2140
rect 3200 2130 3250 2140
rect 6400 2130 6450 2140
rect 7850 2130 7900 2140
rect 8350 2130 8400 2140
rect 9300 2130 9350 2140
rect 9450 2130 9500 2140
rect 9700 2130 9800 2140
rect 1900 2120 1950 2130
rect 2200 2120 2300 2130
rect 2350 2120 2400 2130
rect 2700 2120 2850 2130
rect 3200 2120 3250 2130
rect 6400 2120 6450 2130
rect 7850 2120 7900 2130
rect 8350 2120 8400 2130
rect 9300 2120 9350 2130
rect 9450 2120 9500 2130
rect 9700 2120 9800 2130
rect 1900 2110 1950 2120
rect 2200 2110 2300 2120
rect 2350 2110 2400 2120
rect 2700 2110 2850 2120
rect 3200 2110 3250 2120
rect 6400 2110 6450 2120
rect 7850 2110 7900 2120
rect 8350 2110 8400 2120
rect 9300 2110 9350 2120
rect 9450 2110 9500 2120
rect 9700 2110 9800 2120
rect 1900 2100 1950 2110
rect 2200 2100 2300 2110
rect 2350 2100 2400 2110
rect 2700 2100 2850 2110
rect 3200 2100 3250 2110
rect 6400 2100 6450 2110
rect 7850 2100 7900 2110
rect 8350 2100 8400 2110
rect 9300 2100 9350 2110
rect 9450 2100 9500 2110
rect 9700 2100 9800 2110
rect 1900 2090 1950 2100
rect 2150 2090 2250 2100
rect 3200 2090 3250 2100
rect 6400 2090 6450 2100
rect 6800 2090 6900 2100
rect 7900 2090 8000 2100
rect 8350 2090 8400 2100
rect 1900 2080 1950 2090
rect 2150 2080 2250 2090
rect 3200 2080 3250 2090
rect 6400 2080 6450 2090
rect 6800 2080 6900 2090
rect 7900 2080 8000 2090
rect 8350 2080 8400 2090
rect 1900 2070 1950 2080
rect 2150 2070 2250 2080
rect 3200 2070 3250 2080
rect 6400 2070 6450 2080
rect 6800 2070 6900 2080
rect 7900 2070 8000 2080
rect 8350 2070 8400 2080
rect 1900 2060 1950 2070
rect 2150 2060 2250 2070
rect 3200 2060 3250 2070
rect 6400 2060 6450 2070
rect 6800 2060 6900 2070
rect 7900 2060 8000 2070
rect 8350 2060 8400 2070
rect 1900 2050 1950 2060
rect 2150 2050 2250 2060
rect 3200 2050 3250 2060
rect 6400 2050 6450 2060
rect 6800 2050 6900 2060
rect 7900 2050 8000 2060
rect 8350 2050 8400 2060
rect 1900 2040 2000 2050
rect 2050 2040 2200 2050
rect 3150 2040 3200 2050
rect 6400 2040 6450 2050
rect 6850 2040 6950 2050
rect 8350 2040 8400 2050
rect 9450 2040 9500 2050
rect 9600 2040 9650 2050
rect 1900 2030 2000 2040
rect 2050 2030 2200 2040
rect 3150 2030 3200 2040
rect 6400 2030 6450 2040
rect 6850 2030 6950 2040
rect 8350 2030 8400 2040
rect 9450 2030 9500 2040
rect 9600 2030 9650 2040
rect 1900 2020 2000 2030
rect 2050 2020 2200 2030
rect 3150 2020 3200 2030
rect 6400 2020 6450 2030
rect 6850 2020 6950 2030
rect 8350 2020 8400 2030
rect 9450 2020 9500 2030
rect 9600 2020 9650 2030
rect 1900 2010 2000 2020
rect 2050 2010 2200 2020
rect 3150 2010 3200 2020
rect 6400 2010 6450 2020
rect 6850 2010 6950 2020
rect 8350 2010 8400 2020
rect 9450 2010 9500 2020
rect 9600 2010 9650 2020
rect 1900 2000 2000 2010
rect 2050 2000 2200 2010
rect 3150 2000 3200 2010
rect 6400 2000 6450 2010
rect 6850 2000 6950 2010
rect 8350 2000 8400 2010
rect 9450 2000 9500 2010
rect 9600 2000 9650 2010
rect 1900 1990 2200 2000
rect 3100 1990 3200 2000
rect 6400 1990 6450 2000
rect 6850 1990 7050 2000
rect 7950 1990 8000 2000
rect 8350 1990 8400 2000
rect 8450 1990 8550 2000
rect 9050 1990 9150 2000
rect 1900 1980 2200 1990
rect 3100 1980 3200 1990
rect 6400 1980 6450 1990
rect 6850 1980 7050 1990
rect 7950 1980 8000 1990
rect 8350 1980 8400 1990
rect 8450 1980 8550 1990
rect 9050 1980 9150 1990
rect 1900 1970 2200 1980
rect 3100 1970 3200 1980
rect 6400 1970 6450 1980
rect 6850 1970 7050 1980
rect 7950 1970 8000 1980
rect 8350 1970 8400 1980
rect 8450 1970 8550 1980
rect 9050 1970 9150 1980
rect 1900 1960 2200 1970
rect 3100 1960 3200 1970
rect 6400 1960 6450 1970
rect 6850 1960 7050 1970
rect 7950 1960 8000 1970
rect 8350 1960 8400 1970
rect 8450 1960 8550 1970
rect 9050 1960 9150 1970
rect 1900 1950 2200 1960
rect 3100 1950 3200 1960
rect 6400 1950 6450 1960
rect 6850 1950 7050 1960
rect 7950 1950 8000 1960
rect 8350 1950 8400 1960
rect 8450 1950 8550 1960
rect 9050 1950 9150 1960
rect 1900 1940 2150 1950
rect 2500 1940 2750 1950
rect 3100 1940 3200 1950
rect 6850 1940 7300 1950
rect 7850 1940 7950 1950
rect 8350 1940 8400 1950
rect 8450 1940 9150 1950
rect 9600 1940 9750 1950
rect 9850 1940 9990 1950
rect 1900 1930 2150 1940
rect 2500 1930 2750 1940
rect 3100 1930 3200 1940
rect 6850 1930 7300 1940
rect 7850 1930 7950 1940
rect 8350 1930 8400 1940
rect 8450 1930 9150 1940
rect 9600 1930 9750 1940
rect 9850 1930 9990 1940
rect 1900 1920 2150 1930
rect 2500 1920 2750 1930
rect 3100 1920 3200 1930
rect 6850 1920 7300 1930
rect 7850 1920 7950 1930
rect 8350 1920 8400 1930
rect 8450 1920 9150 1930
rect 9600 1920 9750 1930
rect 9850 1920 9990 1930
rect 1900 1910 2150 1920
rect 2500 1910 2750 1920
rect 3100 1910 3200 1920
rect 6850 1910 7300 1920
rect 7850 1910 7950 1920
rect 8350 1910 8400 1920
rect 8450 1910 9150 1920
rect 9600 1910 9750 1920
rect 9850 1910 9990 1920
rect 1900 1900 2150 1910
rect 2500 1900 2750 1910
rect 3100 1900 3200 1910
rect 6850 1900 7300 1910
rect 7850 1900 7950 1910
rect 8350 1900 8400 1910
rect 8450 1900 9150 1910
rect 9600 1900 9750 1910
rect 9850 1900 9990 1910
rect 1900 1890 2150 1900
rect 2350 1890 2400 1900
rect 2850 1890 2950 1900
rect 3100 1890 3250 1900
rect 6850 1890 7300 1900
rect 7850 1890 7950 1900
rect 8350 1890 8400 1900
rect 8450 1890 8650 1900
rect 8950 1890 9250 1900
rect 9650 1890 9700 1900
rect 9750 1890 9800 1900
rect 9950 1890 9990 1900
rect 1900 1880 2150 1890
rect 2350 1880 2400 1890
rect 2850 1880 2950 1890
rect 3100 1880 3250 1890
rect 6850 1880 7300 1890
rect 7850 1880 7950 1890
rect 8350 1880 8400 1890
rect 8450 1880 8650 1890
rect 8950 1880 9250 1890
rect 9650 1880 9700 1890
rect 9750 1880 9800 1890
rect 9950 1880 9990 1890
rect 1900 1870 2150 1880
rect 2350 1870 2400 1880
rect 2850 1870 2950 1880
rect 3100 1870 3250 1880
rect 6850 1870 7300 1880
rect 7850 1870 7950 1880
rect 8350 1870 8400 1880
rect 8450 1870 8650 1880
rect 8950 1870 9250 1880
rect 9650 1870 9700 1880
rect 9750 1870 9800 1880
rect 9950 1870 9990 1880
rect 1900 1860 2150 1870
rect 2350 1860 2400 1870
rect 2850 1860 2950 1870
rect 3100 1860 3250 1870
rect 6850 1860 7300 1870
rect 7850 1860 7950 1870
rect 8350 1860 8400 1870
rect 8450 1860 8650 1870
rect 8950 1860 9250 1870
rect 9650 1860 9700 1870
rect 9750 1860 9800 1870
rect 9950 1860 9990 1870
rect 1900 1850 2150 1860
rect 2350 1850 2400 1860
rect 2850 1850 2950 1860
rect 3100 1850 3250 1860
rect 6850 1850 7300 1860
rect 7850 1850 7950 1860
rect 8350 1850 8400 1860
rect 8450 1850 8650 1860
rect 8950 1850 9250 1860
rect 9650 1850 9700 1860
rect 9750 1850 9800 1860
rect 9950 1850 9990 1860
rect 1900 1840 2300 1850
rect 2900 1840 2950 1850
rect 3150 1840 3250 1850
rect 6850 1840 7300 1850
rect 7850 1840 7950 1850
rect 8500 1840 8650 1850
rect 8950 1840 9100 1850
rect 9200 1840 9450 1850
rect 9650 1840 9700 1850
rect 9750 1840 9800 1850
rect 1900 1830 2300 1840
rect 2900 1830 2950 1840
rect 3150 1830 3250 1840
rect 6850 1830 7300 1840
rect 7850 1830 7950 1840
rect 8500 1830 8650 1840
rect 8950 1830 9100 1840
rect 9200 1830 9450 1840
rect 9650 1830 9700 1840
rect 9750 1830 9800 1840
rect 1900 1820 2300 1830
rect 2900 1820 2950 1830
rect 3150 1820 3250 1830
rect 6850 1820 7300 1830
rect 7850 1820 7950 1830
rect 8500 1820 8650 1830
rect 8950 1820 9100 1830
rect 9200 1820 9450 1830
rect 9650 1820 9700 1830
rect 9750 1820 9800 1830
rect 1900 1810 2300 1820
rect 2900 1810 2950 1820
rect 3150 1810 3250 1820
rect 6850 1810 7300 1820
rect 7850 1810 7950 1820
rect 8500 1810 8650 1820
rect 8950 1810 9100 1820
rect 9200 1810 9450 1820
rect 9650 1810 9700 1820
rect 9750 1810 9800 1820
rect 1900 1800 2300 1810
rect 2900 1800 2950 1810
rect 3150 1800 3250 1810
rect 6850 1800 7300 1810
rect 7850 1800 7950 1810
rect 8500 1800 8650 1810
rect 8950 1800 9100 1810
rect 9200 1800 9450 1810
rect 9650 1800 9700 1810
rect 9750 1800 9800 1810
rect 1900 1790 2050 1800
rect 2200 1790 2350 1800
rect 2750 1790 2800 1800
rect 3150 1790 3250 1800
rect 4100 1790 4200 1800
rect 6850 1790 7300 1800
rect 7900 1790 7950 1800
rect 8500 1790 8600 1800
rect 8900 1790 9100 1800
rect 9200 1790 9250 1800
rect 9750 1790 9800 1800
rect 9900 1790 9990 1800
rect 1900 1780 2050 1790
rect 2200 1780 2350 1790
rect 2750 1780 2800 1790
rect 3150 1780 3250 1790
rect 4100 1780 4200 1790
rect 6850 1780 7300 1790
rect 7900 1780 7950 1790
rect 8500 1780 8600 1790
rect 8900 1780 9100 1790
rect 9200 1780 9250 1790
rect 9750 1780 9800 1790
rect 9900 1780 9990 1790
rect 1900 1770 2050 1780
rect 2200 1770 2350 1780
rect 2750 1770 2800 1780
rect 3150 1770 3250 1780
rect 4100 1770 4200 1780
rect 6850 1770 7300 1780
rect 7900 1770 7950 1780
rect 8500 1770 8600 1780
rect 8900 1770 9100 1780
rect 9200 1770 9250 1780
rect 9750 1770 9800 1780
rect 9900 1770 9990 1780
rect 1900 1760 2050 1770
rect 2200 1760 2350 1770
rect 2750 1760 2800 1770
rect 3150 1760 3250 1770
rect 4100 1760 4200 1770
rect 6850 1760 7300 1770
rect 7900 1760 7950 1770
rect 8500 1760 8600 1770
rect 8900 1760 9100 1770
rect 9200 1760 9250 1770
rect 9750 1760 9800 1770
rect 9900 1760 9990 1770
rect 1900 1750 2050 1760
rect 2200 1750 2350 1760
rect 2750 1750 2800 1760
rect 3150 1750 3250 1760
rect 4100 1750 4200 1760
rect 6850 1750 7300 1760
rect 7900 1750 7950 1760
rect 8500 1750 8600 1760
rect 8900 1750 9100 1760
rect 9200 1750 9250 1760
rect 9750 1750 9800 1760
rect 9900 1750 9990 1760
rect 1950 1740 2050 1750
rect 2400 1740 2700 1750
rect 3150 1740 3200 1750
rect 4150 1740 4200 1750
rect 5250 1740 5300 1750
rect 6850 1740 7050 1750
rect 7100 1740 7300 1750
rect 7900 1740 7950 1750
rect 8300 1740 8350 1750
rect 8500 1740 8600 1750
rect 8900 1740 9100 1750
rect 9200 1740 9250 1750
rect 9800 1740 9850 1750
rect 9900 1740 9950 1750
rect 1950 1730 2050 1740
rect 2400 1730 2700 1740
rect 3150 1730 3200 1740
rect 4150 1730 4200 1740
rect 5250 1730 5300 1740
rect 6850 1730 7050 1740
rect 7100 1730 7300 1740
rect 7900 1730 7950 1740
rect 8300 1730 8350 1740
rect 8500 1730 8600 1740
rect 8900 1730 9100 1740
rect 9200 1730 9250 1740
rect 9800 1730 9850 1740
rect 9900 1730 9950 1740
rect 1950 1720 2050 1730
rect 2400 1720 2700 1730
rect 3150 1720 3200 1730
rect 4150 1720 4200 1730
rect 5250 1720 5300 1730
rect 6850 1720 7050 1730
rect 7100 1720 7300 1730
rect 7900 1720 7950 1730
rect 8300 1720 8350 1730
rect 8500 1720 8600 1730
rect 8900 1720 9100 1730
rect 9200 1720 9250 1730
rect 9800 1720 9850 1730
rect 9900 1720 9950 1730
rect 1950 1710 2050 1720
rect 2400 1710 2700 1720
rect 3150 1710 3200 1720
rect 4150 1710 4200 1720
rect 5250 1710 5300 1720
rect 6850 1710 7050 1720
rect 7100 1710 7300 1720
rect 7900 1710 7950 1720
rect 8300 1710 8350 1720
rect 8500 1710 8600 1720
rect 8900 1710 9100 1720
rect 9200 1710 9250 1720
rect 9800 1710 9850 1720
rect 9900 1710 9950 1720
rect 1950 1700 2050 1710
rect 2400 1700 2700 1710
rect 3150 1700 3200 1710
rect 4150 1700 4200 1710
rect 5250 1700 5300 1710
rect 6850 1700 7050 1710
rect 7100 1700 7300 1710
rect 7900 1700 7950 1710
rect 8300 1700 8350 1710
rect 8500 1700 8600 1710
rect 8900 1700 9100 1710
rect 9200 1700 9250 1710
rect 9800 1700 9850 1710
rect 9900 1700 9950 1710
rect 1950 1690 2050 1700
rect 2450 1690 2700 1700
rect 3100 1690 3200 1700
rect 4100 1690 4150 1700
rect 6850 1690 7000 1700
rect 7150 1690 7300 1700
rect 7900 1690 7950 1700
rect 8300 1690 8350 1700
rect 8550 1690 8650 1700
rect 8850 1690 9100 1700
rect 9200 1690 9250 1700
rect 9700 1690 9800 1700
rect 9850 1690 9950 1700
rect 1950 1680 2050 1690
rect 2450 1680 2700 1690
rect 3100 1680 3200 1690
rect 4100 1680 4150 1690
rect 6850 1680 7000 1690
rect 7150 1680 7300 1690
rect 7900 1680 7950 1690
rect 8300 1680 8350 1690
rect 8550 1680 8650 1690
rect 8850 1680 9100 1690
rect 9200 1680 9250 1690
rect 9700 1680 9800 1690
rect 9850 1680 9950 1690
rect 1950 1670 2050 1680
rect 2450 1670 2700 1680
rect 3100 1670 3200 1680
rect 4100 1670 4150 1680
rect 6850 1670 7000 1680
rect 7150 1670 7300 1680
rect 7900 1670 7950 1680
rect 8300 1670 8350 1680
rect 8550 1670 8650 1680
rect 8850 1670 9100 1680
rect 9200 1670 9250 1680
rect 9700 1670 9800 1680
rect 9850 1670 9950 1680
rect 1950 1660 2050 1670
rect 2450 1660 2700 1670
rect 3100 1660 3200 1670
rect 4100 1660 4150 1670
rect 6850 1660 7000 1670
rect 7150 1660 7300 1670
rect 7900 1660 7950 1670
rect 8300 1660 8350 1670
rect 8550 1660 8650 1670
rect 8850 1660 9100 1670
rect 9200 1660 9250 1670
rect 9700 1660 9800 1670
rect 9850 1660 9950 1670
rect 1950 1650 2050 1660
rect 2450 1650 2700 1660
rect 3100 1650 3200 1660
rect 4100 1650 4150 1660
rect 6850 1650 7000 1660
rect 7150 1650 7300 1660
rect 7900 1650 7950 1660
rect 8300 1650 8350 1660
rect 8550 1650 8650 1660
rect 8850 1650 9100 1660
rect 9200 1650 9250 1660
rect 9700 1650 9800 1660
rect 9850 1650 9950 1660
rect 2000 1640 2100 1650
rect 2400 1640 2750 1650
rect 3050 1640 3150 1650
rect 5450 1640 5500 1650
rect 6850 1640 7000 1650
rect 7150 1640 7350 1650
rect 7900 1640 7950 1650
rect 8300 1640 8350 1650
rect 8500 1640 8650 1650
rect 8800 1640 9150 1650
rect 9200 1640 9250 1650
rect 9800 1640 9900 1650
rect 2000 1630 2100 1640
rect 2400 1630 2750 1640
rect 3050 1630 3150 1640
rect 5450 1630 5500 1640
rect 6850 1630 7000 1640
rect 7150 1630 7350 1640
rect 7900 1630 7950 1640
rect 8300 1630 8350 1640
rect 8500 1630 8650 1640
rect 8800 1630 9150 1640
rect 9200 1630 9250 1640
rect 9800 1630 9900 1640
rect 2000 1620 2100 1630
rect 2400 1620 2750 1630
rect 3050 1620 3150 1630
rect 5450 1620 5500 1630
rect 6850 1620 7000 1630
rect 7150 1620 7350 1630
rect 7900 1620 7950 1630
rect 8300 1620 8350 1630
rect 8500 1620 8650 1630
rect 8800 1620 9150 1630
rect 9200 1620 9250 1630
rect 9800 1620 9900 1630
rect 2000 1610 2100 1620
rect 2400 1610 2750 1620
rect 3050 1610 3150 1620
rect 5450 1610 5500 1620
rect 6850 1610 7000 1620
rect 7150 1610 7350 1620
rect 7900 1610 7950 1620
rect 8300 1610 8350 1620
rect 8500 1610 8650 1620
rect 8800 1610 9150 1620
rect 9200 1610 9250 1620
rect 9800 1610 9900 1620
rect 2000 1600 2100 1610
rect 2400 1600 2750 1610
rect 3050 1600 3150 1610
rect 5450 1600 5500 1610
rect 6850 1600 7000 1610
rect 7150 1600 7350 1610
rect 7900 1600 7950 1610
rect 8300 1600 8350 1610
rect 8500 1600 8650 1610
rect 8800 1600 9150 1610
rect 9200 1600 9250 1610
rect 9800 1600 9900 1610
rect 2000 1590 2150 1600
rect 2400 1590 2700 1600
rect 3000 1590 3100 1600
rect 4250 1590 4300 1600
rect 5650 1590 5700 1600
rect 6850 1590 7000 1600
rect 7150 1590 7350 1600
rect 7900 1590 8000 1600
rect 8450 1590 9050 1600
rect 9700 1590 9800 1600
rect 9850 1590 9990 1600
rect 2000 1580 2150 1590
rect 2400 1580 2700 1590
rect 3000 1580 3100 1590
rect 4250 1580 4300 1590
rect 5650 1580 5700 1590
rect 6850 1580 7000 1590
rect 7150 1580 7350 1590
rect 7900 1580 8000 1590
rect 8450 1580 9050 1590
rect 9700 1580 9800 1590
rect 9850 1580 9990 1590
rect 2000 1570 2150 1580
rect 2400 1570 2700 1580
rect 3000 1570 3100 1580
rect 4250 1570 4300 1580
rect 5650 1570 5700 1580
rect 6850 1570 7000 1580
rect 7150 1570 7350 1580
rect 7900 1570 8000 1580
rect 8450 1570 9050 1580
rect 9700 1570 9800 1580
rect 9850 1570 9990 1580
rect 2000 1560 2150 1570
rect 2400 1560 2700 1570
rect 3000 1560 3100 1570
rect 4250 1560 4300 1570
rect 5650 1560 5700 1570
rect 6850 1560 7000 1570
rect 7150 1560 7350 1570
rect 7900 1560 8000 1570
rect 8450 1560 9050 1570
rect 9700 1560 9800 1570
rect 9850 1560 9990 1570
rect 2000 1550 2150 1560
rect 2400 1550 2700 1560
rect 3000 1550 3100 1560
rect 4250 1550 4300 1560
rect 5650 1550 5700 1560
rect 6850 1550 7000 1560
rect 7150 1550 7350 1560
rect 7900 1550 8000 1560
rect 8450 1550 9050 1560
rect 9700 1550 9800 1560
rect 9850 1550 9990 1560
rect 2050 1540 2200 1550
rect 2900 1540 3050 1550
rect 4250 1540 4350 1550
rect 6850 1540 7000 1550
rect 7200 1540 7350 1550
rect 7900 1540 8000 1550
rect 8450 1540 9050 1550
rect 9850 1540 9950 1550
rect 2050 1530 2200 1540
rect 2900 1530 3050 1540
rect 4250 1530 4350 1540
rect 6850 1530 7000 1540
rect 7200 1530 7350 1540
rect 7900 1530 8000 1540
rect 8450 1530 9050 1540
rect 9850 1530 9950 1540
rect 2050 1520 2200 1530
rect 2900 1520 3050 1530
rect 4250 1520 4350 1530
rect 6850 1520 7000 1530
rect 7200 1520 7350 1530
rect 7900 1520 8000 1530
rect 8450 1520 9050 1530
rect 9850 1520 9950 1530
rect 2050 1510 2200 1520
rect 2900 1510 3050 1520
rect 4250 1510 4350 1520
rect 6850 1510 7000 1520
rect 7200 1510 7350 1520
rect 7900 1510 8000 1520
rect 8450 1510 9050 1520
rect 9850 1510 9950 1520
rect 2050 1500 2200 1510
rect 2900 1500 3050 1510
rect 4250 1500 4350 1510
rect 6850 1500 7000 1510
rect 7200 1500 7350 1510
rect 7900 1500 8000 1510
rect 8450 1500 9050 1510
rect 9850 1500 9950 1510
rect 2100 1490 2250 1500
rect 2900 1490 2950 1500
rect 4150 1490 4250 1500
rect 6850 1490 6950 1500
rect 7250 1490 7350 1500
rect 7900 1490 8000 1500
rect 8250 1490 8300 1500
rect 8450 1490 8600 1500
rect 8700 1490 9200 1500
rect 9600 1490 9700 1500
rect 9800 1490 9850 1500
rect 9900 1490 9950 1500
rect 2100 1480 2250 1490
rect 2900 1480 2950 1490
rect 4150 1480 4250 1490
rect 6850 1480 6950 1490
rect 7250 1480 7350 1490
rect 7900 1480 8000 1490
rect 8250 1480 8300 1490
rect 8450 1480 8600 1490
rect 8700 1480 9200 1490
rect 9600 1480 9700 1490
rect 9800 1480 9850 1490
rect 9900 1480 9950 1490
rect 2100 1470 2250 1480
rect 2900 1470 2950 1480
rect 4150 1470 4250 1480
rect 6850 1470 6950 1480
rect 7250 1470 7350 1480
rect 7900 1470 8000 1480
rect 8250 1470 8300 1480
rect 8450 1470 8600 1480
rect 8700 1470 9200 1480
rect 9600 1470 9700 1480
rect 9800 1470 9850 1480
rect 9900 1470 9950 1480
rect 2100 1460 2250 1470
rect 2900 1460 2950 1470
rect 4150 1460 4250 1470
rect 6850 1460 6950 1470
rect 7250 1460 7350 1470
rect 7900 1460 8000 1470
rect 8250 1460 8300 1470
rect 8450 1460 8600 1470
rect 8700 1460 9200 1470
rect 9600 1460 9700 1470
rect 9800 1460 9850 1470
rect 9900 1460 9950 1470
rect 2100 1450 2250 1460
rect 2900 1450 2950 1460
rect 4150 1450 4250 1460
rect 6850 1450 6950 1460
rect 7250 1450 7350 1460
rect 7900 1450 8000 1460
rect 8250 1450 8300 1460
rect 8450 1450 8600 1460
rect 8700 1450 9200 1460
rect 9600 1450 9700 1460
rect 9800 1450 9850 1460
rect 9900 1450 9950 1460
rect 2150 1440 2250 1450
rect 2850 1440 2900 1450
rect 4200 1440 4300 1450
rect 4350 1440 4400 1450
rect 6850 1440 6900 1450
rect 7250 1440 7350 1450
rect 7950 1440 8000 1450
rect 8200 1440 8250 1450
rect 8450 1440 9100 1450
rect 9550 1440 9700 1450
rect 9750 1440 9800 1450
rect 9950 1440 9990 1450
rect 2150 1430 2250 1440
rect 2850 1430 2900 1440
rect 4200 1430 4300 1440
rect 4350 1430 4400 1440
rect 6850 1430 6900 1440
rect 7250 1430 7350 1440
rect 7950 1430 8000 1440
rect 8200 1430 8250 1440
rect 8450 1430 9100 1440
rect 9550 1430 9700 1440
rect 9750 1430 9800 1440
rect 9950 1430 9990 1440
rect 2150 1420 2250 1430
rect 2850 1420 2900 1430
rect 4200 1420 4300 1430
rect 4350 1420 4400 1430
rect 6850 1420 6900 1430
rect 7250 1420 7350 1430
rect 7950 1420 8000 1430
rect 8200 1420 8250 1430
rect 8450 1420 9100 1430
rect 9550 1420 9700 1430
rect 9750 1420 9800 1430
rect 9950 1420 9990 1430
rect 2150 1410 2250 1420
rect 2850 1410 2900 1420
rect 4200 1410 4300 1420
rect 4350 1410 4400 1420
rect 6850 1410 6900 1420
rect 7250 1410 7350 1420
rect 7950 1410 8000 1420
rect 8200 1410 8250 1420
rect 8450 1410 9100 1420
rect 9550 1410 9700 1420
rect 9750 1410 9800 1420
rect 9950 1410 9990 1420
rect 2150 1400 2250 1410
rect 2850 1400 2900 1410
rect 4200 1400 4300 1410
rect 4350 1400 4400 1410
rect 6850 1400 6900 1410
rect 7250 1400 7350 1410
rect 7950 1400 8000 1410
rect 8200 1400 8250 1410
rect 8450 1400 9100 1410
rect 9550 1400 9700 1410
rect 9750 1400 9800 1410
rect 9950 1400 9990 1410
rect 2200 1390 2350 1400
rect 2750 1390 2800 1400
rect 4250 1390 4400 1400
rect 7250 1390 7350 1400
rect 7950 1390 8000 1400
rect 8150 1390 8200 1400
rect 8450 1390 9100 1400
rect 9200 1390 9300 1400
rect 9600 1390 9650 1400
rect 9750 1390 9850 1400
rect 9900 1390 9990 1400
rect 2200 1380 2350 1390
rect 2750 1380 2800 1390
rect 4250 1380 4400 1390
rect 7250 1380 7350 1390
rect 7950 1380 8000 1390
rect 8150 1380 8200 1390
rect 8450 1380 9100 1390
rect 9200 1380 9300 1390
rect 9600 1380 9650 1390
rect 9750 1380 9850 1390
rect 9900 1380 9990 1390
rect 2200 1370 2350 1380
rect 2750 1370 2800 1380
rect 4250 1370 4400 1380
rect 7250 1370 7350 1380
rect 7950 1370 8000 1380
rect 8150 1370 8200 1380
rect 8450 1370 9100 1380
rect 9200 1370 9300 1380
rect 9600 1370 9650 1380
rect 9750 1370 9850 1380
rect 9900 1370 9990 1380
rect 2200 1360 2350 1370
rect 2750 1360 2800 1370
rect 4250 1360 4400 1370
rect 7250 1360 7350 1370
rect 7950 1360 8000 1370
rect 8150 1360 8200 1370
rect 8450 1360 9100 1370
rect 9200 1360 9300 1370
rect 9600 1360 9650 1370
rect 9750 1360 9850 1370
rect 9900 1360 9990 1370
rect 2200 1350 2350 1360
rect 2750 1350 2800 1360
rect 4250 1350 4400 1360
rect 7250 1350 7350 1360
rect 7950 1350 8000 1360
rect 8150 1350 8200 1360
rect 8450 1350 9100 1360
rect 9200 1350 9300 1360
rect 9600 1350 9650 1360
rect 9750 1350 9850 1360
rect 9900 1350 9990 1360
rect 2350 1340 2500 1350
rect 2650 1340 2750 1350
rect 3600 1340 3650 1350
rect 4250 1340 4300 1350
rect 7300 1340 7350 1350
rect 7950 1340 8150 1350
rect 8450 1340 9150 1350
rect 9250 1340 9300 1350
rect 9600 1340 9650 1350
rect 9700 1340 9850 1350
rect 9950 1340 9990 1350
rect 2350 1330 2500 1340
rect 2650 1330 2750 1340
rect 3600 1330 3650 1340
rect 4250 1330 4300 1340
rect 7300 1330 7350 1340
rect 7950 1330 8150 1340
rect 8450 1330 9150 1340
rect 9250 1330 9300 1340
rect 9600 1330 9650 1340
rect 9700 1330 9850 1340
rect 9950 1330 9990 1340
rect 2350 1320 2500 1330
rect 2650 1320 2750 1330
rect 3600 1320 3650 1330
rect 4250 1320 4300 1330
rect 7300 1320 7350 1330
rect 7950 1320 8150 1330
rect 8450 1320 9150 1330
rect 9250 1320 9300 1330
rect 9600 1320 9650 1330
rect 9700 1320 9850 1330
rect 9950 1320 9990 1330
rect 2350 1310 2500 1320
rect 2650 1310 2750 1320
rect 3600 1310 3650 1320
rect 4250 1310 4300 1320
rect 7300 1310 7350 1320
rect 7950 1310 8150 1320
rect 8450 1310 9150 1320
rect 9250 1310 9300 1320
rect 9600 1310 9650 1320
rect 9700 1310 9850 1320
rect 9950 1310 9990 1320
rect 2350 1300 2500 1310
rect 2650 1300 2750 1310
rect 3600 1300 3650 1310
rect 4250 1300 4300 1310
rect 7300 1300 7350 1310
rect 7950 1300 8150 1310
rect 8450 1300 9150 1310
rect 9250 1300 9300 1310
rect 9600 1300 9650 1310
rect 9700 1300 9850 1310
rect 9950 1300 9990 1310
rect 3500 1290 3550 1300
rect 4200 1290 4250 1300
rect 4400 1290 4450 1300
rect 7300 1290 7350 1300
rect 7950 1290 8150 1300
rect 8450 1290 9050 1300
rect 9600 1290 9650 1300
rect 9700 1290 9750 1300
rect 3500 1280 3550 1290
rect 4200 1280 4250 1290
rect 4400 1280 4450 1290
rect 7300 1280 7350 1290
rect 7950 1280 8150 1290
rect 8450 1280 9050 1290
rect 9600 1280 9650 1290
rect 9700 1280 9750 1290
rect 3500 1270 3550 1280
rect 4200 1270 4250 1280
rect 4400 1270 4450 1280
rect 7300 1270 7350 1280
rect 7950 1270 8150 1280
rect 8450 1270 9050 1280
rect 9600 1270 9650 1280
rect 9700 1270 9750 1280
rect 3500 1260 3550 1270
rect 4200 1260 4250 1270
rect 4400 1260 4450 1270
rect 7300 1260 7350 1270
rect 7950 1260 8150 1270
rect 8450 1260 9050 1270
rect 9600 1260 9650 1270
rect 9700 1260 9750 1270
rect 3500 1250 3550 1260
rect 4200 1250 4250 1260
rect 4400 1250 4450 1260
rect 7300 1250 7350 1260
rect 7950 1250 8150 1260
rect 8450 1250 9050 1260
rect 9600 1250 9650 1260
rect 9700 1250 9750 1260
rect 3650 1240 3700 1250
rect 3750 1240 3800 1250
rect 4200 1240 4250 1250
rect 4400 1240 4450 1250
rect 5250 1240 5350 1250
rect 7300 1240 7350 1250
rect 7950 1240 8150 1250
rect 8450 1240 8850 1250
rect 9300 1240 9350 1250
rect 9650 1240 9750 1250
rect 9800 1240 9850 1250
rect 9900 1240 9950 1250
rect 3650 1230 3700 1240
rect 3750 1230 3800 1240
rect 4200 1230 4250 1240
rect 4400 1230 4450 1240
rect 5250 1230 5350 1240
rect 7300 1230 7350 1240
rect 7950 1230 8150 1240
rect 8450 1230 8850 1240
rect 9300 1230 9350 1240
rect 9650 1230 9750 1240
rect 9800 1230 9850 1240
rect 9900 1230 9950 1240
rect 3650 1220 3700 1230
rect 3750 1220 3800 1230
rect 4200 1220 4250 1230
rect 4400 1220 4450 1230
rect 5250 1220 5350 1230
rect 7300 1220 7350 1230
rect 7950 1220 8150 1230
rect 8450 1220 8850 1230
rect 9300 1220 9350 1230
rect 9650 1220 9750 1230
rect 9800 1220 9850 1230
rect 9900 1220 9950 1230
rect 3650 1210 3700 1220
rect 3750 1210 3800 1220
rect 4200 1210 4250 1220
rect 4400 1210 4450 1220
rect 5250 1210 5350 1220
rect 7300 1210 7350 1220
rect 7950 1210 8150 1220
rect 8450 1210 8850 1220
rect 9300 1210 9350 1220
rect 9650 1210 9750 1220
rect 9800 1210 9850 1220
rect 9900 1210 9950 1220
rect 3650 1200 3700 1210
rect 3750 1200 3800 1210
rect 4200 1200 4250 1210
rect 4400 1200 4450 1210
rect 5250 1200 5350 1210
rect 7300 1200 7350 1210
rect 7950 1200 8150 1210
rect 8450 1200 8850 1210
rect 9300 1200 9350 1210
rect 9650 1200 9750 1210
rect 9800 1200 9850 1210
rect 9900 1200 9950 1210
rect 3700 1190 3750 1200
rect 3800 1190 3850 1200
rect 4200 1190 4250 1200
rect 6700 1190 6800 1200
rect 7300 1190 7350 1200
rect 7950 1190 8150 1200
rect 8450 1190 8700 1200
rect 9100 1190 9150 1200
rect 9300 1190 9400 1200
rect 9500 1190 9600 1200
rect 9650 1190 9700 1200
rect 9800 1190 9850 1200
rect 9950 1190 9990 1200
rect 3700 1180 3750 1190
rect 3800 1180 3850 1190
rect 4200 1180 4250 1190
rect 6700 1180 6800 1190
rect 7300 1180 7350 1190
rect 7950 1180 8150 1190
rect 8450 1180 8700 1190
rect 9100 1180 9150 1190
rect 9300 1180 9400 1190
rect 9500 1180 9600 1190
rect 9650 1180 9700 1190
rect 9800 1180 9850 1190
rect 9950 1180 9990 1190
rect 3700 1170 3750 1180
rect 3800 1170 3850 1180
rect 4200 1170 4250 1180
rect 6700 1170 6800 1180
rect 7300 1170 7350 1180
rect 7950 1170 8150 1180
rect 8450 1170 8700 1180
rect 9100 1170 9150 1180
rect 9300 1170 9400 1180
rect 9500 1170 9600 1180
rect 9650 1170 9700 1180
rect 9800 1170 9850 1180
rect 9950 1170 9990 1180
rect 3700 1160 3750 1170
rect 3800 1160 3850 1170
rect 4200 1160 4250 1170
rect 6700 1160 6800 1170
rect 7300 1160 7350 1170
rect 7950 1160 8150 1170
rect 8450 1160 8700 1170
rect 9100 1160 9150 1170
rect 9300 1160 9400 1170
rect 9500 1160 9600 1170
rect 9650 1160 9700 1170
rect 9800 1160 9850 1170
rect 9950 1160 9990 1170
rect 3700 1150 3750 1160
rect 3800 1150 3850 1160
rect 4200 1150 4250 1160
rect 6700 1150 6800 1160
rect 7300 1150 7350 1160
rect 7950 1150 8150 1160
rect 8450 1150 8700 1160
rect 9100 1150 9150 1160
rect 9300 1150 9400 1160
rect 9500 1150 9600 1160
rect 9650 1150 9700 1160
rect 9800 1150 9850 1160
rect 9950 1150 9990 1160
rect 3750 1140 3800 1150
rect 3900 1140 3950 1150
rect 6600 1140 6650 1150
rect 6750 1140 6800 1150
rect 7300 1140 7350 1150
rect 8000 1140 8150 1150
rect 8450 1140 8650 1150
rect 9100 1140 9150 1150
rect 9300 1140 9400 1150
rect 9500 1140 9550 1150
rect 9600 1140 9650 1150
rect 9850 1140 9990 1150
rect 3750 1130 3800 1140
rect 3900 1130 3950 1140
rect 6600 1130 6650 1140
rect 6750 1130 6800 1140
rect 7300 1130 7350 1140
rect 8000 1130 8150 1140
rect 8450 1130 8650 1140
rect 9100 1130 9150 1140
rect 9300 1130 9400 1140
rect 9500 1130 9550 1140
rect 9600 1130 9650 1140
rect 9850 1130 9990 1140
rect 3750 1120 3800 1130
rect 3900 1120 3950 1130
rect 6600 1120 6650 1130
rect 6750 1120 6800 1130
rect 7300 1120 7350 1130
rect 8000 1120 8150 1130
rect 8450 1120 8650 1130
rect 9100 1120 9150 1130
rect 9300 1120 9400 1130
rect 9500 1120 9550 1130
rect 9600 1120 9650 1130
rect 9850 1120 9990 1130
rect 3750 1110 3800 1120
rect 3900 1110 3950 1120
rect 6600 1110 6650 1120
rect 6750 1110 6800 1120
rect 7300 1110 7350 1120
rect 8000 1110 8150 1120
rect 8450 1110 8650 1120
rect 9100 1110 9150 1120
rect 9300 1110 9400 1120
rect 9500 1110 9550 1120
rect 9600 1110 9650 1120
rect 9850 1110 9990 1120
rect 3750 1100 3800 1110
rect 3900 1100 3950 1110
rect 6600 1100 6650 1110
rect 6750 1100 6800 1110
rect 7300 1100 7350 1110
rect 8000 1100 8150 1110
rect 8450 1100 8650 1110
rect 9100 1100 9150 1110
rect 9300 1100 9400 1110
rect 9500 1100 9550 1110
rect 9600 1100 9650 1110
rect 9850 1100 9990 1110
rect 3750 1090 3850 1100
rect 3950 1090 4000 1100
rect 4450 1090 4500 1100
rect 6550 1090 6600 1100
rect 6750 1090 6800 1100
rect 7300 1090 7350 1100
rect 8000 1090 8150 1100
rect 8500 1090 8550 1100
rect 9100 1090 9450 1100
rect 9500 1090 9600 1100
rect 9700 1090 9750 1100
rect 9850 1090 9950 1100
rect 3750 1080 3850 1090
rect 3950 1080 4000 1090
rect 4450 1080 4500 1090
rect 6550 1080 6600 1090
rect 6750 1080 6800 1090
rect 7300 1080 7350 1090
rect 8000 1080 8150 1090
rect 8500 1080 8550 1090
rect 9100 1080 9450 1090
rect 9500 1080 9600 1090
rect 9700 1080 9750 1090
rect 9850 1080 9950 1090
rect 3750 1070 3850 1080
rect 3950 1070 4000 1080
rect 4450 1070 4500 1080
rect 6550 1070 6600 1080
rect 6750 1070 6800 1080
rect 7300 1070 7350 1080
rect 8000 1070 8150 1080
rect 8500 1070 8550 1080
rect 9100 1070 9450 1080
rect 9500 1070 9600 1080
rect 9700 1070 9750 1080
rect 9850 1070 9950 1080
rect 3750 1060 3850 1070
rect 3950 1060 4000 1070
rect 4450 1060 4500 1070
rect 6550 1060 6600 1070
rect 6750 1060 6800 1070
rect 7300 1060 7350 1070
rect 8000 1060 8150 1070
rect 8500 1060 8550 1070
rect 9100 1060 9450 1070
rect 9500 1060 9600 1070
rect 9700 1060 9750 1070
rect 9850 1060 9950 1070
rect 3750 1050 3850 1060
rect 3950 1050 4000 1060
rect 4450 1050 4500 1060
rect 6550 1050 6600 1060
rect 6750 1050 6800 1060
rect 7300 1050 7350 1060
rect 8000 1050 8150 1060
rect 8500 1050 8550 1060
rect 9100 1050 9450 1060
rect 9500 1050 9600 1060
rect 9700 1050 9750 1060
rect 9850 1050 9950 1060
rect 2100 1040 2200 1050
rect 3850 1040 3900 1050
rect 4050 1040 4100 1050
rect 4200 1040 4250 1050
rect 4550 1040 4650 1050
rect 6500 1040 6550 1050
rect 6750 1040 6800 1050
rect 7300 1040 7350 1050
rect 8000 1040 8100 1050
rect 8400 1040 8500 1050
rect 9250 1040 9300 1050
rect 9350 1040 9450 1050
rect 9500 1040 9600 1050
rect 9700 1040 9750 1050
rect 9850 1040 9990 1050
rect 2100 1030 2200 1040
rect 3850 1030 3900 1040
rect 4050 1030 4100 1040
rect 4200 1030 4250 1040
rect 4550 1030 4650 1040
rect 6500 1030 6550 1040
rect 6750 1030 6800 1040
rect 7300 1030 7350 1040
rect 8000 1030 8100 1040
rect 8400 1030 8500 1040
rect 9250 1030 9300 1040
rect 9350 1030 9450 1040
rect 9500 1030 9600 1040
rect 9700 1030 9750 1040
rect 9850 1030 9990 1040
rect 2100 1020 2200 1030
rect 3850 1020 3900 1030
rect 4050 1020 4100 1030
rect 4200 1020 4250 1030
rect 4550 1020 4650 1030
rect 6500 1020 6550 1030
rect 6750 1020 6800 1030
rect 7300 1020 7350 1030
rect 8000 1020 8100 1030
rect 8400 1020 8500 1030
rect 9250 1020 9300 1030
rect 9350 1020 9450 1030
rect 9500 1020 9600 1030
rect 9700 1020 9750 1030
rect 9850 1020 9990 1030
rect 2100 1010 2200 1020
rect 3850 1010 3900 1020
rect 4050 1010 4100 1020
rect 4200 1010 4250 1020
rect 4550 1010 4650 1020
rect 6500 1010 6550 1020
rect 6750 1010 6800 1020
rect 7300 1010 7350 1020
rect 8000 1010 8100 1020
rect 8400 1010 8500 1020
rect 9250 1010 9300 1020
rect 9350 1010 9450 1020
rect 9500 1010 9600 1020
rect 9700 1010 9750 1020
rect 9850 1010 9990 1020
rect 2100 1000 2200 1010
rect 3850 1000 3900 1010
rect 4050 1000 4100 1010
rect 4200 1000 4250 1010
rect 4550 1000 4650 1010
rect 6500 1000 6550 1010
rect 6750 1000 6800 1010
rect 7300 1000 7350 1010
rect 8000 1000 8100 1010
rect 8400 1000 8500 1010
rect 9250 1000 9300 1010
rect 9350 1000 9450 1010
rect 9500 1000 9600 1010
rect 9700 1000 9750 1010
rect 9850 1000 9990 1010
rect 2050 990 2300 1000
rect 3850 990 3900 1000
rect 4100 990 4200 1000
rect 4700 990 4750 1000
rect 6500 990 6550 1000
rect 6850 990 6900 1000
rect 7300 990 7350 1000
rect 8000 990 8100 1000
rect 8400 990 8550 1000
rect 9150 990 9250 1000
rect 9450 990 9550 1000
rect 9750 990 9850 1000
rect 2050 980 2300 990
rect 3850 980 3900 990
rect 4100 980 4200 990
rect 4700 980 4750 990
rect 6500 980 6550 990
rect 6850 980 6900 990
rect 7300 980 7350 990
rect 8000 980 8100 990
rect 8400 980 8550 990
rect 9150 980 9250 990
rect 9450 980 9550 990
rect 9750 980 9850 990
rect 2050 970 2300 980
rect 3850 970 3900 980
rect 4100 970 4200 980
rect 4700 970 4750 980
rect 6500 970 6550 980
rect 6850 970 6900 980
rect 7300 970 7350 980
rect 8000 970 8100 980
rect 8400 970 8550 980
rect 9150 970 9250 980
rect 9450 970 9550 980
rect 9750 970 9850 980
rect 2050 960 2300 970
rect 3850 960 3900 970
rect 4100 960 4200 970
rect 4700 960 4750 970
rect 6500 960 6550 970
rect 6850 960 6900 970
rect 7300 960 7350 970
rect 8000 960 8100 970
rect 8400 960 8550 970
rect 9150 960 9250 970
rect 9450 960 9550 970
rect 9750 960 9850 970
rect 2050 950 2300 960
rect 3850 950 3900 960
rect 4100 950 4200 960
rect 4700 950 4750 960
rect 6500 950 6550 960
rect 6850 950 6900 960
rect 7300 950 7350 960
rect 8000 950 8100 960
rect 8400 950 8550 960
rect 9150 950 9250 960
rect 9450 950 9550 960
rect 9750 950 9850 960
rect 2050 940 2700 950
rect 3850 940 3900 950
rect 4800 940 4850 950
rect 6500 940 6550 950
rect 6800 940 6900 950
rect 7300 940 7350 950
rect 8000 940 8100 950
rect 8450 940 8550 950
rect 9150 940 9200 950
rect 9500 940 9550 950
rect 2050 930 2700 940
rect 3850 930 3900 940
rect 4800 930 4850 940
rect 6500 930 6550 940
rect 6800 930 6900 940
rect 7300 930 7350 940
rect 8000 930 8100 940
rect 8450 930 8550 940
rect 9150 930 9200 940
rect 9500 930 9550 940
rect 2050 920 2700 930
rect 3850 920 3900 930
rect 4800 920 4850 930
rect 6500 920 6550 930
rect 6800 920 6900 930
rect 7300 920 7350 930
rect 8000 920 8100 930
rect 8450 920 8550 930
rect 9150 920 9200 930
rect 9500 920 9550 930
rect 2050 910 2700 920
rect 3850 910 3900 920
rect 4800 910 4850 920
rect 6500 910 6550 920
rect 6800 910 6900 920
rect 7300 910 7350 920
rect 8000 910 8100 920
rect 8450 910 8550 920
rect 9150 910 9200 920
rect 9500 910 9550 920
rect 2050 900 2700 910
rect 3850 900 3900 910
rect 4800 900 4850 910
rect 6500 900 6550 910
rect 6800 900 6900 910
rect 7300 900 7350 910
rect 8000 900 8100 910
rect 8450 900 8550 910
rect 9150 900 9200 910
rect 9500 900 9550 910
rect 700 890 750 900
rect 2050 890 2650 900
rect 3900 890 4050 900
rect 6500 890 6600 900
rect 6800 890 6900 900
rect 7300 890 7350 900
rect 8000 890 8100 900
rect 8450 890 8600 900
rect 9150 890 9200 900
rect 9400 890 9500 900
rect 700 880 750 890
rect 2050 880 2650 890
rect 3900 880 4050 890
rect 6500 880 6600 890
rect 6800 880 6900 890
rect 7300 880 7350 890
rect 8000 880 8100 890
rect 8450 880 8600 890
rect 9150 880 9200 890
rect 9400 880 9500 890
rect 700 870 750 880
rect 2050 870 2650 880
rect 3900 870 4050 880
rect 6500 870 6600 880
rect 6800 870 6900 880
rect 7300 870 7350 880
rect 8000 870 8100 880
rect 8450 870 8600 880
rect 9150 870 9200 880
rect 9400 870 9500 880
rect 700 860 750 870
rect 2050 860 2650 870
rect 3900 860 4050 870
rect 6500 860 6600 870
rect 6800 860 6900 870
rect 7300 860 7350 870
rect 8000 860 8100 870
rect 8450 860 8600 870
rect 9150 860 9200 870
rect 9400 860 9500 870
rect 700 850 750 860
rect 2050 850 2650 860
rect 3900 850 4050 860
rect 6500 850 6600 860
rect 6800 850 6900 860
rect 7300 850 7350 860
rect 8000 850 8100 860
rect 8450 850 8600 860
rect 9150 850 9200 860
rect 9400 850 9500 860
rect 700 840 750 850
rect 2100 840 2600 850
rect 4000 840 4050 850
rect 4250 840 4350 850
rect 4850 840 4900 850
rect 6500 840 6600 850
rect 6800 840 6900 850
rect 7300 840 7350 850
rect 8000 840 8100 850
rect 700 830 750 840
rect 2100 830 2600 840
rect 4000 830 4050 840
rect 4250 830 4350 840
rect 4850 830 4900 840
rect 6500 830 6600 840
rect 6800 830 6900 840
rect 7300 830 7350 840
rect 8000 830 8100 840
rect 700 820 750 830
rect 2100 820 2600 830
rect 4000 820 4050 830
rect 4250 820 4350 830
rect 4850 820 4900 830
rect 6500 820 6600 830
rect 6800 820 6900 830
rect 7300 820 7350 830
rect 8000 820 8100 830
rect 700 810 750 820
rect 2100 810 2600 820
rect 4000 810 4050 820
rect 4250 810 4350 820
rect 4850 810 4900 820
rect 6500 810 6600 820
rect 6800 810 6900 820
rect 7300 810 7350 820
rect 8000 810 8100 820
rect 700 800 750 810
rect 2100 800 2600 810
rect 4000 800 4050 810
rect 4250 800 4350 810
rect 4850 800 4900 810
rect 6500 800 6600 810
rect 6800 800 6900 810
rect 7300 800 7350 810
rect 8000 800 8100 810
rect 650 790 700 800
rect 2100 790 2350 800
rect 2450 790 2550 800
rect 4000 790 4050 800
rect 4300 790 4350 800
rect 6550 790 6600 800
rect 6800 790 6900 800
rect 7250 790 7350 800
rect 8050 790 8100 800
rect 9200 790 9250 800
rect 9350 790 9450 800
rect 650 780 700 790
rect 2100 780 2350 790
rect 2450 780 2550 790
rect 4000 780 4050 790
rect 4300 780 4350 790
rect 6550 780 6600 790
rect 6800 780 6900 790
rect 7250 780 7350 790
rect 8050 780 8100 790
rect 9200 780 9250 790
rect 9350 780 9450 790
rect 650 770 700 780
rect 2100 770 2350 780
rect 2450 770 2550 780
rect 4000 770 4050 780
rect 4300 770 4350 780
rect 6550 770 6600 780
rect 6800 770 6900 780
rect 7250 770 7350 780
rect 8050 770 8100 780
rect 9200 770 9250 780
rect 9350 770 9450 780
rect 650 760 700 770
rect 2100 760 2350 770
rect 2450 760 2550 770
rect 4000 760 4050 770
rect 4300 760 4350 770
rect 6550 760 6600 770
rect 6800 760 6900 770
rect 7250 760 7350 770
rect 8050 760 8100 770
rect 9200 760 9250 770
rect 9350 760 9450 770
rect 650 750 700 760
rect 2100 750 2350 760
rect 2450 750 2550 760
rect 4000 750 4050 760
rect 4300 750 4350 760
rect 6550 750 6600 760
rect 6800 750 6900 760
rect 7250 750 7350 760
rect 8050 750 8100 760
rect 9200 750 9250 760
rect 9350 750 9450 760
rect 650 740 700 750
rect 1150 740 1200 750
rect 2100 740 2250 750
rect 2400 740 2450 750
rect 3450 740 3550 750
rect 4000 740 4200 750
rect 4750 740 4850 750
rect 6550 740 6600 750
rect 7250 740 7350 750
rect 8050 740 8100 750
rect 9200 740 9250 750
rect 9300 740 9350 750
rect 650 730 700 740
rect 1150 730 1200 740
rect 2100 730 2250 740
rect 2400 730 2450 740
rect 3450 730 3550 740
rect 4000 730 4200 740
rect 4750 730 4850 740
rect 6550 730 6600 740
rect 7250 730 7350 740
rect 8050 730 8100 740
rect 9200 730 9250 740
rect 9300 730 9350 740
rect 650 720 700 730
rect 1150 720 1200 730
rect 2100 720 2250 730
rect 2400 720 2450 730
rect 3450 720 3550 730
rect 4000 720 4200 730
rect 4750 720 4850 730
rect 6550 720 6600 730
rect 7250 720 7350 730
rect 8050 720 8100 730
rect 9200 720 9250 730
rect 9300 720 9350 730
rect 650 710 700 720
rect 1150 710 1200 720
rect 2100 710 2250 720
rect 2400 710 2450 720
rect 3450 710 3550 720
rect 4000 710 4200 720
rect 4750 710 4850 720
rect 6550 710 6600 720
rect 7250 710 7350 720
rect 8050 710 8100 720
rect 9200 710 9250 720
rect 9300 710 9350 720
rect 650 700 700 710
rect 1150 700 1200 710
rect 2100 700 2250 710
rect 2400 700 2450 710
rect 3450 700 3550 710
rect 4000 700 4200 710
rect 4750 700 4850 710
rect 6550 700 6600 710
rect 7250 700 7350 710
rect 8050 700 8100 710
rect 9200 700 9250 710
rect 9300 700 9350 710
rect 1100 690 1150 700
rect 2150 690 2350 700
rect 3300 690 3350 700
rect 4050 690 4100 700
rect 4150 690 4200 700
rect 4800 690 4900 700
rect 6600 690 6650 700
rect 6900 690 6950 700
rect 7250 690 7300 700
rect 8050 690 8100 700
rect 9200 690 9250 700
rect 9300 690 9400 700
rect 9600 690 9700 700
rect 1100 680 1150 690
rect 2150 680 2350 690
rect 3300 680 3350 690
rect 4050 680 4100 690
rect 4150 680 4200 690
rect 4800 680 4900 690
rect 6600 680 6650 690
rect 6900 680 6950 690
rect 7250 680 7300 690
rect 8050 680 8100 690
rect 9200 680 9250 690
rect 9300 680 9400 690
rect 9600 680 9700 690
rect 1100 670 1150 680
rect 2150 670 2350 680
rect 3300 670 3350 680
rect 4050 670 4100 680
rect 4150 670 4200 680
rect 4800 670 4900 680
rect 6600 670 6650 680
rect 6900 670 6950 680
rect 7250 670 7300 680
rect 8050 670 8100 680
rect 9200 670 9250 680
rect 9300 670 9400 680
rect 9600 670 9700 680
rect 1100 660 1150 670
rect 2150 660 2350 670
rect 3300 660 3350 670
rect 4050 660 4100 670
rect 4150 660 4200 670
rect 4800 660 4900 670
rect 6600 660 6650 670
rect 6900 660 6950 670
rect 7250 660 7300 670
rect 8050 660 8100 670
rect 9200 660 9250 670
rect 9300 660 9400 670
rect 9600 660 9700 670
rect 1100 650 1150 660
rect 2150 650 2350 660
rect 3300 650 3350 660
rect 4050 650 4100 660
rect 4150 650 4200 660
rect 4800 650 4900 660
rect 6600 650 6650 660
rect 6900 650 6950 660
rect 7250 650 7300 660
rect 8050 650 8100 660
rect 9200 650 9250 660
rect 9300 650 9400 660
rect 9600 650 9700 660
rect 2150 640 2200 650
rect 3250 640 3300 650
rect 4050 640 4150 650
rect 4650 640 4700 650
rect 4800 640 4850 650
rect 4900 640 4950 650
rect 6600 640 6700 650
rect 6850 640 6950 650
rect 7200 640 7300 650
rect 9200 640 9350 650
rect 9600 640 9700 650
rect 2150 630 2200 640
rect 3250 630 3300 640
rect 4050 630 4150 640
rect 4650 630 4700 640
rect 4800 630 4850 640
rect 4900 630 4950 640
rect 6600 630 6700 640
rect 6850 630 6950 640
rect 7200 630 7300 640
rect 9200 630 9350 640
rect 9600 630 9700 640
rect 2150 620 2200 630
rect 3250 620 3300 630
rect 4050 620 4150 630
rect 4650 620 4700 630
rect 4800 620 4850 630
rect 4900 620 4950 630
rect 6600 620 6700 630
rect 6850 620 6950 630
rect 7200 620 7300 630
rect 9200 620 9350 630
rect 9600 620 9700 630
rect 2150 610 2200 620
rect 3250 610 3300 620
rect 4050 610 4150 620
rect 4650 610 4700 620
rect 4800 610 4850 620
rect 4900 610 4950 620
rect 6600 610 6700 620
rect 6850 610 6950 620
rect 7200 610 7300 620
rect 9200 610 9350 620
rect 9600 610 9700 620
rect 2150 600 2200 610
rect 3250 600 3300 610
rect 4050 600 4150 610
rect 4650 600 4700 610
rect 4800 600 4850 610
rect 4900 600 4950 610
rect 6600 600 6700 610
rect 6850 600 6950 610
rect 7200 600 7300 610
rect 9200 600 9350 610
rect 9600 600 9700 610
rect 350 590 450 600
rect 550 590 650 600
rect 950 590 1050 600
rect 3100 590 3150 600
rect 4350 590 4500 600
rect 4550 590 4600 600
rect 4900 590 4950 600
rect 6650 590 6700 600
rect 6850 590 6900 600
rect 6950 590 7000 600
rect 7150 590 7300 600
rect 9200 590 9250 600
rect 350 580 450 590
rect 550 580 650 590
rect 950 580 1050 590
rect 3100 580 3150 590
rect 4350 580 4500 590
rect 4550 580 4600 590
rect 4900 580 4950 590
rect 6650 580 6700 590
rect 6850 580 6900 590
rect 6950 580 7000 590
rect 7150 580 7300 590
rect 9200 580 9250 590
rect 350 570 450 580
rect 550 570 650 580
rect 950 570 1050 580
rect 3100 570 3150 580
rect 4350 570 4500 580
rect 4550 570 4600 580
rect 4900 570 4950 580
rect 6650 570 6700 580
rect 6850 570 6900 580
rect 6950 570 7000 580
rect 7150 570 7300 580
rect 9200 570 9250 580
rect 350 560 450 570
rect 550 560 650 570
rect 950 560 1050 570
rect 3100 560 3150 570
rect 4350 560 4500 570
rect 4550 560 4600 570
rect 4900 560 4950 570
rect 6650 560 6700 570
rect 6850 560 6900 570
rect 6950 560 7000 570
rect 7150 560 7300 570
rect 9200 560 9250 570
rect 350 550 450 560
rect 550 550 650 560
rect 950 550 1050 560
rect 3100 550 3150 560
rect 4350 550 4500 560
rect 4550 550 4600 560
rect 4900 550 4950 560
rect 6650 550 6700 560
rect 6850 550 6900 560
rect 6950 550 7000 560
rect 7150 550 7300 560
rect 9200 550 9250 560
rect 350 540 400 550
rect 500 540 600 550
rect 1250 540 1300 550
rect 1450 540 1500 550
rect 2950 540 3000 550
rect 4200 540 4300 550
rect 4750 540 4800 550
rect 4850 540 4900 550
rect 6700 540 6750 550
rect 6850 540 6900 550
rect 6950 540 7250 550
rect 9250 540 9300 550
rect 9900 540 9990 550
rect 350 530 400 540
rect 500 530 600 540
rect 1250 530 1300 540
rect 1450 530 1500 540
rect 2950 530 3000 540
rect 4200 530 4300 540
rect 4750 530 4800 540
rect 4850 530 4900 540
rect 6700 530 6750 540
rect 6850 530 6900 540
rect 6950 530 7250 540
rect 9250 530 9300 540
rect 9900 530 9990 540
rect 350 520 400 530
rect 500 520 600 530
rect 1250 520 1300 530
rect 1450 520 1500 530
rect 2950 520 3000 530
rect 4200 520 4300 530
rect 4750 520 4800 530
rect 4850 520 4900 530
rect 6700 520 6750 530
rect 6850 520 6900 530
rect 6950 520 7250 530
rect 9250 520 9300 530
rect 9900 520 9990 530
rect 350 510 400 520
rect 500 510 600 520
rect 1250 510 1300 520
rect 1450 510 1500 520
rect 2950 510 3000 520
rect 4200 510 4300 520
rect 4750 510 4800 520
rect 4850 510 4900 520
rect 6700 510 6750 520
rect 6850 510 6900 520
rect 6950 510 7250 520
rect 9250 510 9300 520
rect 9900 510 9990 520
rect 350 500 400 510
rect 500 500 600 510
rect 1250 500 1300 510
rect 1450 500 1500 510
rect 2950 500 3000 510
rect 4200 500 4300 510
rect 4750 500 4800 510
rect 4850 500 4900 510
rect 6700 500 6750 510
rect 6850 500 6900 510
rect 6950 500 7250 510
rect 9250 500 9300 510
rect 9900 500 9990 510
rect 150 490 300 500
rect 400 490 500 500
rect 1150 490 1200 500
rect 1500 490 1550 500
rect 2800 490 2900 500
rect 4200 490 4250 500
rect 4750 490 4800 500
rect 4850 490 4900 500
rect 6700 490 7250 500
rect 9850 490 9990 500
rect 150 480 300 490
rect 400 480 500 490
rect 1150 480 1200 490
rect 1500 480 1550 490
rect 2800 480 2900 490
rect 4200 480 4250 490
rect 4750 480 4800 490
rect 4850 480 4900 490
rect 6700 480 7250 490
rect 9850 480 9990 490
rect 150 470 300 480
rect 400 470 500 480
rect 1150 470 1200 480
rect 1500 470 1550 480
rect 2800 470 2900 480
rect 4200 470 4250 480
rect 4750 470 4800 480
rect 4850 470 4900 480
rect 6700 470 7250 480
rect 9850 470 9990 480
rect 150 460 300 470
rect 400 460 500 470
rect 1150 460 1200 470
rect 1500 460 1550 470
rect 2800 460 2900 470
rect 4200 460 4250 470
rect 4750 460 4800 470
rect 4850 460 4900 470
rect 6700 460 7250 470
rect 9850 460 9990 470
rect 150 450 300 460
rect 400 450 500 460
rect 1150 450 1200 460
rect 1500 450 1550 460
rect 2800 450 2900 460
rect 4200 450 4250 460
rect 4750 450 4800 460
rect 4850 450 4900 460
rect 6700 450 7250 460
rect 9850 450 9990 460
rect 100 440 150 450
rect 250 440 350 450
rect 1100 440 1150 450
rect 1550 440 1700 450
rect 1800 440 2000 450
rect 2250 440 2300 450
rect 2550 440 2700 450
rect 4150 440 4200 450
rect 4750 440 4800 450
rect 6750 440 7200 450
rect 9200 440 9400 450
rect 100 430 150 440
rect 250 430 350 440
rect 1100 430 1150 440
rect 1550 430 1700 440
rect 1800 430 2000 440
rect 2250 430 2300 440
rect 2550 430 2700 440
rect 4150 430 4200 440
rect 4750 430 4800 440
rect 6750 430 7200 440
rect 9200 430 9400 440
rect 100 420 150 430
rect 250 420 350 430
rect 1100 420 1150 430
rect 1550 420 1700 430
rect 1800 420 2000 430
rect 2250 420 2300 430
rect 2550 420 2700 430
rect 4150 420 4200 430
rect 4750 420 4800 430
rect 6750 420 7200 430
rect 9200 420 9400 430
rect 100 410 150 420
rect 250 410 350 420
rect 1100 410 1150 420
rect 1550 410 1700 420
rect 1800 410 2000 420
rect 2250 410 2300 420
rect 2550 410 2700 420
rect 4150 410 4200 420
rect 4750 410 4800 420
rect 6750 410 7200 420
rect 9200 410 9400 420
rect 100 400 150 410
rect 250 400 350 410
rect 1100 400 1150 410
rect 1550 400 1700 410
rect 1800 400 2000 410
rect 2250 400 2300 410
rect 2550 400 2700 410
rect 4150 400 4200 410
rect 4750 400 4800 410
rect 6750 400 7200 410
rect 9200 400 9400 410
rect 50 390 100 400
rect 300 390 350 400
rect 4150 390 4200 400
rect 6800 390 7200 400
rect 9200 390 9250 400
rect 9400 390 9450 400
rect 50 380 100 390
rect 300 380 350 390
rect 4150 380 4200 390
rect 6800 380 7200 390
rect 9200 380 9250 390
rect 9400 380 9450 390
rect 50 370 100 380
rect 300 370 350 380
rect 4150 370 4200 380
rect 6800 370 7200 380
rect 9200 370 9250 380
rect 9400 370 9450 380
rect 50 360 100 370
rect 300 360 350 370
rect 4150 360 4200 370
rect 6800 360 7200 370
rect 9200 360 9250 370
rect 9400 360 9450 370
rect 50 350 100 360
rect 300 350 350 360
rect 4150 350 4200 360
rect 6800 350 7200 360
rect 9200 350 9250 360
rect 9400 350 9450 360
rect 50 340 100 350
rect 250 340 350 350
rect 1050 340 1100 350
rect 4100 340 4150 350
rect 4300 340 4350 350
rect 4750 340 4950 350
rect 6850 340 7100 350
rect 9150 340 9250 350
rect 9400 340 9450 350
rect 50 330 100 340
rect 250 330 350 340
rect 1050 330 1100 340
rect 4100 330 4150 340
rect 4300 330 4350 340
rect 4750 330 4950 340
rect 6850 330 7100 340
rect 9150 330 9250 340
rect 9400 330 9450 340
rect 50 320 100 330
rect 250 320 350 330
rect 1050 320 1100 330
rect 4100 320 4150 330
rect 4300 320 4350 330
rect 4750 320 4950 330
rect 6850 320 7100 330
rect 9150 320 9250 330
rect 9400 320 9450 330
rect 50 310 100 320
rect 250 310 350 320
rect 1050 310 1100 320
rect 4100 310 4150 320
rect 4300 310 4350 320
rect 4750 310 4950 320
rect 6850 310 7100 320
rect 9150 310 9250 320
rect 9400 310 9450 320
rect 50 300 100 310
rect 250 300 350 310
rect 1050 300 1100 310
rect 4100 300 4150 310
rect 4300 300 4350 310
rect 4750 300 4950 310
rect 6850 300 7100 310
rect 9150 300 9250 310
rect 9400 300 9450 310
rect 50 290 350 300
rect 500 290 600 300
rect 700 290 800 300
rect 4050 290 4100 300
rect 4250 290 4500 300
rect 4700 290 5000 300
rect 9100 290 9200 300
rect 9450 290 9500 300
rect 50 280 350 290
rect 500 280 600 290
rect 700 280 800 290
rect 4050 280 4100 290
rect 4250 280 4500 290
rect 4700 280 5000 290
rect 9100 280 9200 290
rect 9450 280 9500 290
rect 50 270 350 280
rect 500 270 600 280
rect 700 270 800 280
rect 4050 270 4100 280
rect 4250 270 4500 280
rect 4700 270 5000 280
rect 9100 270 9200 280
rect 9450 270 9500 280
rect 50 260 350 270
rect 500 260 600 270
rect 700 260 800 270
rect 4050 260 4100 270
rect 4250 260 4500 270
rect 4700 260 5000 270
rect 9100 260 9200 270
rect 9450 260 9500 270
rect 50 250 350 260
rect 500 250 600 260
rect 700 250 800 260
rect 4050 250 4100 260
rect 4250 250 4500 260
rect 4700 250 5000 260
rect 9100 250 9200 260
rect 9450 250 9500 260
rect 250 240 350 250
rect 450 240 600 250
rect 700 240 850 250
rect 1000 240 1050 250
rect 4100 240 4150 250
rect 4250 240 4300 250
rect 4400 240 4500 250
rect 4650 240 4850 250
rect 4900 240 5000 250
rect 9100 240 9200 250
rect 9350 240 9450 250
rect 9750 240 9900 250
rect 9950 240 9990 250
rect 250 230 350 240
rect 450 230 600 240
rect 700 230 850 240
rect 1000 230 1050 240
rect 4100 230 4150 240
rect 4250 230 4300 240
rect 4400 230 4500 240
rect 4650 230 4850 240
rect 4900 230 5000 240
rect 9100 230 9200 240
rect 9350 230 9450 240
rect 9750 230 9900 240
rect 9950 230 9990 240
rect 250 220 350 230
rect 450 220 600 230
rect 700 220 850 230
rect 1000 220 1050 230
rect 4100 220 4150 230
rect 4250 220 4300 230
rect 4400 220 4500 230
rect 4650 220 4850 230
rect 4900 220 5000 230
rect 9100 220 9200 230
rect 9350 220 9450 230
rect 9750 220 9900 230
rect 9950 220 9990 230
rect 250 210 350 220
rect 450 210 600 220
rect 700 210 850 220
rect 1000 210 1050 220
rect 4100 210 4150 220
rect 4250 210 4300 220
rect 4400 210 4500 220
rect 4650 210 4850 220
rect 4900 210 5000 220
rect 9100 210 9200 220
rect 9350 210 9450 220
rect 9750 210 9900 220
rect 9950 210 9990 220
rect 250 200 350 210
rect 450 200 600 210
rect 700 200 850 210
rect 1000 200 1050 210
rect 4100 200 4150 210
rect 4250 200 4300 210
rect 4400 200 4500 210
rect 4650 200 4850 210
rect 4900 200 5000 210
rect 9100 200 9200 210
rect 9350 200 9450 210
rect 9750 200 9900 210
rect 9950 200 9990 210
rect 1000 190 1050 200
rect 4600 190 4800 200
rect 4900 190 5000 200
rect 9100 190 9150 200
rect 9700 190 9750 200
rect 1000 180 1050 190
rect 4600 180 4800 190
rect 4900 180 5000 190
rect 9100 180 9150 190
rect 9700 180 9750 190
rect 1000 170 1050 180
rect 4600 170 4800 180
rect 4900 170 5000 180
rect 9100 170 9150 180
rect 9700 170 9750 180
rect 1000 160 1050 170
rect 4600 160 4800 170
rect 4900 160 5000 170
rect 9100 160 9150 170
rect 9700 160 9750 170
rect 1000 150 1050 160
rect 4600 150 4800 160
rect 4900 150 5000 160
rect 9100 150 9150 160
rect 9700 150 9750 160
rect 0 140 100 150
rect 1000 140 1050 150
rect 4200 140 4250 150
rect 4950 140 5000 150
rect 9100 140 9150 150
rect 9350 140 9450 150
rect 9700 140 9750 150
rect 0 130 100 140
rect 1000 130 1050 140
rect 4200 130 4250 140
rect 4950 130 5000 140
rect 9100 130 9150 140
rect 9350 130 9450 140
rect 9700 130 9750 140
rect 0 120 100 130
rect 1000 120 1050 130
rect 4200 120 4250 130
rect 4950 120 5000 130
rect 9100 120 9150 130
rect 9350 120 9450 130
rect 9700 120 9750 130
rect 0 110 100 120
rect 1000 110 1050 120
rect 4200 110 4250 120
rect 4950 110 5000 120
rect 9100 110 9150 120
rect 9350 110 9450 120
rect 9700 110 9750 120
rect 0 100 100 110
rect 1000 100 1050 110
rect 4200 100 4250 110
rect 4950 100 5000 110
rect 9100 100 9150 110
rect 9350 100 9450 110
rect 9700 100 9750 110
rect 0 90 100 100
rect 1000 90 1050 100
rect 4250 90 4300 100
rect 4950 90 5050 100
rect 8900 90 8950 100
rect 9050 90 9150 100
rect 9450 90 9750 100
rect 0 80 100 90
rect 1000 80 1050 90
rect 4250 80 4300 90
rect 4950 80 5050 90
rect 8900 80 8950 90
rect 9050 80 9150 90
rect 9450 80 9750 90
rect 0 70 100 80
rect 1000 70 1050 80
rect 4250 70 4300 80
rect 4950 70 5050 80
rect 8900 70 8950 80
rect 9050 70 9150 80
rect 9450 70 9750 80
rect 0 60 100 70
rect 1000 60 1050 70
rect 4250 60 4300 70
rect 4950 60 5050 70
rect 8900 60 8950 70
rect 9050 60 9150 70
rect 9450 60 9750 70
rect 0 50 100 60
rect 1000 50 1050 60
rect 4250 50 4300 60
rect 4950 50 5050 60
rect 8900 50 8950 60
rect 9050 50 9150 60
rect 9450 50 9750 60
rect 0 40 100 50
rect 1000 40 1050 50
rect 4300 40 4350 50
rect 4950 40 5000 50
rect 9050 40 9150 50
rect 9500 40 9750 50
rect 9950 40 9990 50
rect 0 30 100 40
rect 1000 30 1050 40
rect 4300 30 4350 40
rect 4950 30 5000 40
rect 9050 30 9150 40
rect 9500 30 9750 40
rect 9950 30 9990 40
rect 0 20 100 30
rect 1000 20 1050 30
rect 4300 20 4350 30
rect 4950 20 5000 30
rect 9050 20 9150 30
rect 9500 20 9750 30
rect 9950 20 9990 30
rect 0 10 100 20
rect 1000 10 1050 20
rect 4300 10 4350 20
rect 4950 10 5000 20
rect 9050 10 9150 20
rect 9500 10 9750 20
rect 9950 10 9990 20
rect 0 0 100 10
rect 1000 0 1050 10
rect 4300 0 4350 10
rect 4950 0 5000 10
rect 9050 0 9150 10
rect 9500 0 9750 10
rect 9950 0 9990 10
<< end >>
