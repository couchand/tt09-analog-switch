VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_couchand_analog_switch
  CLASS BLOCK ;
  FOREIGN tt_um_couchand_analog_switch ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.088000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
        RECT 151.500 -0.500 153.000 0.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.176000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
        RECT 132.500 -0.500 134.000 0.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.776000 ;
    PORT
      LAYER met4 ;
        RECT 138.000 225.760 139.000 226.000 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 60.000 116.200 62.970 121.900 ;
      LAYER nwell ;
        RECT 63.500 117.500 66.470 121.990 ;
        RECT 63.500 116.150 66.700 117.500 ;
        RECT 63.500 116.140 66.950 116.150 ;
      LAYER pwell ;
        RECT 60.000 110.350 62.970 116.050 ;
      LAYER nwell ;
        RECT 63.500 116.000 66.970 116.140 ;
        RECT 64.000 110.350 66.970 116.000 ;
      LAYER li1 ;
        RECT 54.000 123.000 55.500 123.500 ;
        RECT 54.000 122.500 66.000 123.000 ;
        RECT 54.000 122.000 55.500 122.500 ;
        RECT 64.000 121.810 66.000 122.500 ;
        RECT 60.180 121.550 62.790 121.720 ;
        RECT 60.180 119.200 60.350 121.550 ;
        RECT 60.980 121.040 61.340 121.210 ;
        RECT 61.630 121.040 61.990 121.210 ;
        RECT 60.750 119.200 60.920 120.870 ;
        RECT 60.180 119.025 60.920 119.200 ;
        RECT 60.180 116.550 60.350 119.025 ;
        RECT 60.750 117.230 60.920 119.025 ;
        RECT 61.400 117.230 61.570 120.870 ;
        RECT 62.050 119.200 62.220 120.870 ;
        RECT 62.620 119.200 62.790 121.550 ;
        RECT 62.050 119.025 62.790 119.200 ;
        RECT 62.050 117.230 62.220 119.025 ;
        RECT 60.980 116.890 61.340 117.060 ;
        RECT 61.630 116.890 61.990 117.060 ;
        RECT 62.620 116.550 62.790 119.025 ;
        RECT 60.180 116.380 62.790 116.550 ;
        RECT 63.680 121.640 66.290 121.810 ;
        RECT 63.680 119.200 63.850 121.640 ;
        RECT 64.480 121.130 64.840 121.300 ;
        RECT 65.130 121.130 65.490 121.300 ;
        RECT 64.250 119.200 64.420 120.915 ;
        RECT 63.680 119.025 64.420 119.200 ;
        RECT 63.680 116.550 63.850 119.025 ;
        RECT 64.250 117.275 64.420 119.025 ;
        RECT 64.900 117.275 65.070 120.915 ;
        RECT 65.550 119.200 65.720 120.915 ;
        RECT 66.120 119.200 66.290 121.640 ;
        RECT 65.550 119.025 66.290 119.200 ;
        RECT 65.550 117.275 65.720 119.025 ;
        RECT 64.480 116.890 64.840 117.060 ;
        RECT 65.130 116.890 65.490 117.060 ;
        RECT 66.120 116.550 66.290 119.025 ;
        RECT 63.680 116.450 66.290 116.550 ;
        RECT 60.500 115.870 62.500 116.380 ;
        RECT 63.400 116.200 66.750 116.450 ;
        RECT 64.550 115.960 66.450 116.200 ;
        RECT 60.180 115.700 62.790 115.870 ;
        RECT 60.180 110.700 60.350 115.700 ;
        RECT 60.980 115.190 61.340 115.360 ;
        RECT 61.630 115.190 61.990 115.360 ;
        RECT 60.750 111.380 60.920 115.020 ;
        RECT 61.400 111.380 61.570 115.020 ;
        RECT 62.050 111.380 62.220 115.020 ;
        RECT 60.980 111.040 61.340 111.210 ;
        RECT 61.630 111.040 61.990 111.210 ;
        RECT 62.620 110.700 62.790 115.700 ;
        RECT 60.180 110.530 62.790 110.700 ;
        RECT 64.180 115.790 66.790 115.960 ;
        RECT 64.180 110.700 64.350 115.790 ;
        RECT 64.980 115.280 65.340 115.450 ;
        RECT 65.630 115.280 65.990 115.450 ;
        RECT 64.750 111.425 64.920 115.065 ;
        RECT 65.400 111.425 65.570 115.065 ;
        RECT 66.050 111.425 66.220 115.065 ;
        RECT 64.980 111.040 65.340 111.210 ;
        RECT 65.630 111.040 65.990 111.210 ;
        RECT 66.620 110.700 66.790 115.790 ;
        RECT 64.180 110.530 66.790 110.700 ;
        RECT 54.000 110.000 55.500 110.500 ;
        RECT 60.600 110.300 62.400 110.530 ;
        RECT 60.350 110.000 63.700 110.300 ;
        RECT 54.000 109.500 63.500 110.000 ;
        RECT 54.000 109.000 55.500 109.500 ;
      LAYER mcon ;
        RECT 54.500 122.500 55.000 123.000 ;
        RECT 61.060 121.040 61.260 121.210 ;
        RECT 61.710 121.040 61.910 121.210 ;
        RECT 60.750 117.310 60.920 120.790 ;
        RECT 61.400 117.310 61.570 120.790 ;
        RECT 62.050 117.310 62.220 120.790 ;
        RECT 61.060 116.890 61.260 117.060 ;
        RECT 61.710 116.890 61.910 117.060 ;
        RECT 64.560 121.130 64.760 121.300 ;
        RECT 65.210 121.130 65.410 121.300 ;
        RECT 64.250 117.355 64.420 120.835 ;
        RECT 64.900 117.355 65.070 120.835 ;
        RECT 65.550 117.355 65.720 120.835 ;
        RECT 64.560 116.890 64.760 117.060 ;
        RECT 65.210 116.890 65.410 117.060 ;
        RECT 61.060 115.190 61.260 115.360 ;
        RECT 61.710 115.190 61.910 115.360 ;
        RECT 60.750 111.460 60.920 114.940 ;
        RECT 61.400 111.460 61.570 114.940 ;
        RECT 62.050 111.460 62.220 114.940 ;
        RECT 61.060 111.040 61.260 111.210 ;
        RECT 61.710 111.040 61.910 111.210 ;
        RECT 65.060 115.280 65.260 115.450 ;
        RECT 65.710 115.280 65.910 115.450 ;
        RECT 64.750 111.505 64.920 114.985 ;
        RECT 65.400 111.505 65.570 114.985 ;
        RECT 66.050 111.505 66.220 114.985 ;
        RECT 65.060 111.040 65.260 111.210 ;
        RECT 65.710 111.040 65.910 111.210 ;
        RECT 54.500 109.500 55.000 110.000 ;
      LAYER met1 ;
        RECT 62.500 125.000 64.000 126.500 ;
        RECT 1.000 122.000 55.500 123.500 ;
        RECT 63.000 121.350 63.500 125.000 ;
        RECT 63.000 121.250 65.500 121.350 ;
        RECT 60.975 121.100 65.500 121.250 ;
        RECT 60.975 121.000 63.500 121.100 ;
        RECT 60.720 117.250 60.950 120.850 ;
        RECT 61.370 120.200 61.600 120.850 ;
        RECT 61.300 119.825 61.675 120.200 ;
        RECT 61.370 117.250 61.600 119.825 ;
        RECT 62.020 117.250 62.250 120.850 ;
        RECT 64.220 117.295 64.450 120.895 ;
        RECT 64.870 120.200 65.100 120.895 ;
        RECT 64.800 119.825 65.175 120.200 ;
        RECT 64.870 117.295 65.100 119.825 ;
        RECT 65.520 117.295 65.750 120.895 ;
        RECT 60.975 116.850 65.500 117.100 ;
        RECT 63.600 115.500 63.850 116.850 ;
        RECT 62.950 115.400 63.350 115.500 ;
        RECT 60.950 115.150 63.350 115.400 ;
        RECT 62.950 115.100 63.350 115.150 ;
        RECT 60.720 113.750 60.950 115.000 ;
        RECT 60.650 113.350 61.050 113.750 ;
        RECT 60.720 111.400 60.950 113.350 ;
        RECT 61.370 112.500 61.600 115.000 ;
        RECT 62.020 113.750 62.250 115.000 ;
        RECT 61.950 113.350 62.350 113.750 ;
        RECT 61.300 112.100 61.700 112.500 ;
        RECT 61.370 111.400 61.600 112.100 ;
        RECT 62.020 111.400 62.250 113.350 ;
        RECT 63.100 111.250 63.350 115.100 ;
        RECT 60.950 111.000 63.350 111.250 ;
        RECT 63.600 115.250 66.050 115.500 ;
        RECT 63.600 111.250 63.850 115.250 ;
        RECT 64.720 113.750 64.950 115.045 ;
        RECT 64.650 113.350 65.050 113.750 ;
        RECT 64.720 111.445 64.950 113.350 ;
        RECT 65.370 112.500 65.600 115.045 ;
        RECT 66.020 113.750 66.250 115.045 ;
        RECT 65.950 113.350 66.350 113.750 ;
        RECT 65.300 112.100 65.700 112.500 ;
        RECT 65.370 111.445 65.600 112.100 ;
        RECT 66.020 111.445 66.250 113.350 ;
        RECT 63.600 111.000 66.050 111.250 ;
        RECT 4.000 109.000 55.500 110.500 ;
      LAYER via ;
        RECT 63.000 125.500 63.500 126.000 ;
        RECT 1.500 122.500 2.500 123.000 ;
        RECT 61.350 119.875 61.625 120.150 ;
        RECT 64.850 119.875 65.125 120.150 ;
        RECT 63.000 115.150 63.300 115.450 ;
        RECT 60.700 113.400 61.000 113.700 ;
        RECT 62.000 113.400 62.300 113.700 ;
        RECT 61.350 112.150 61.650 112.450 ;
        RECT 64.700 113.400 65.000 113.700 ;
        RECT 66.000 113.400 66.300 113.700 ;
        RECT 65.350 112.150 65.650 112.450 ;
        RECT 4.500 109.500 5.500 110.000 ;
      LAYER met2 ;
        RECT 62.500 125.000 64.000 126.500 ;
        RECT 1.000 121.500 3.000 124.000 ;
        RECT 61.300 120.150 61.675 120.200 ;
        RECT 64.800 120.150 65.175 120.200 ;
        RECT 61.300 119.875 65.175 120.150 ;
        RECT 61.300 119.825 61.675 119.875 ;
        RECT 63.000 115.500 63.250 119.875 ;
        RECT 64.800 119.825 65.175 119.875 ;
        RECT 62.950 115.100 63.350 115.500 ;
        RECT 71.500 113.800 73.000 114.500 ;
        RECT 60.600 113.300 73.000 113.800 ;
        RECT 71.500 113.000 73.000 113.300 ;
        RECT 61.200 112.000 73.000 112.500 ;
        RECT 71.500 111.000 73.000 112.000 ;
        RECT 4.000 108.500 6.000 111.000 ;
      LAYER via2 ;
        RECT 63.000 125.500 63.500 126.000 ;
        RECT 1.500 122.500 2.500 123.000 ;
        RECT 72.000 113.500 72.500 114.000 ;
        RECT 72.000 111.500 72.500 112.000 ;
        RECT 4.500 109.500 5.500 110.000 ;
      LAYER met3 ;
        RECT 62.500 125.000 64.000 126.500 ;
        RECT 1.000 121.500 3.000 124.000 ;
        RECT 71.500 113.000 73.000 114.500 ;
        RECT 71.500 111.000 153.000 112.500 ;
        RECT 4.000 108.500 6.000 111.000 ;
      LAYER via3 ;
        RECT 63.000 125.500 63.500 126.000 ;
        RECT 1.500 122.500 2.500 123.000 ;
        RECT 72.000 113.500 72.500 114.000 ;
        RECT 152.000 111.500 152.500 112.000 ;
        RECT 4.500 109.500 5.500 110.000 ;
      LAYER met4 ;
        RECT 138.000 224.760 138.310 225.760 ;
        RECT 138.610 224.760 139.000 225.760 ;
        RECT 138.000 126.500 139.000 224.760 ;
        RECT 62.500 125.000 139.000 126.500 ;
        RECT 71.500 113.000 134.000 114.500 ;
        RECT 132.500 1.000 134.000 113.000 ;
        RECT 133.390 0.000 134.000 1.000 ;
        RECT 151.500 1.000 153.000 112.500 ;
        RECT 151.500 0.000 151.810 1.000 ;
        RECT 152.710 0.000 153.000 1.000 ;
  END
END tt_um_couchand_analog_switch
END LIBRARY

