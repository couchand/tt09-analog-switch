magic
tech sky130A
timestamp 1730993132
<< locali >>
rect 5400 12300 5550 12350
rect 5400 12250 5450 12300
rect 5500 12250 6600 12300
rect 5400 12200 5550 12250
rect 6400 12200 6600 12250
rect 5400 11000 5550 11050
rect 5400 10950 5450 11000
rect 5500 10950 6350 11000
rect 5400 10900 5550 10950
<< viali >>
rect 5450 12250 5500 12300
rect 5450 10950 5500 11000
<< metal1 >>
rect 6250 12600 6400 12650
rect 6250 12550 6300 12600
rect 6350 12550 6400 12600
rect 6250 12500 6400 12550
rect 100 12300 5550 12350
rect 100 12250 150 12300
rect 250 12250 5450 12300
rect 5500 12250 5550 12300
rect 100 12200 5550 12250
rect 6300 12100 6350 12500
rect 6950 11650 7100 11700
rect 6950 11640 7000 11650
rect 6380 11600 7000 11640
rect 7050 11600 7100 11650
rect 6380 11590 7100 11600
rect 6950 11550 7100 11590
rect 400 11000 5550 11050
rect 400 10950 450 11000
rect 550 10950 5450 11000
rect 5500 10950 5550 11000
rect 400 10900 5550 10950
<< via1 >>
rect 6300 12550 6350 12600
rect 150 12250 250 12300
rect 7000 11600 7050 11650
rect 450 10950 550 11000
<< metal2 >>
rect 6950 12900 9500 12950
rect 6950 12850 9400 12900
rect 9450 12850 9500 12900
rect 6950 12800 9500 12850
rect 6250 12600 6400 12650
rect 6250 12550 6300 12600
rect 6350 12550 6400 12600
rect 6250 12500 6400 12550
rect 100 12300 300 12400
rect 100 12250 150 12300
rect 250 12250 300 12300
rect 100 12150 300 12250
rect 6950 11650 7100 12800
rect 6950 11600 7000 11650
rect 7050 11600 7100 11650
rect 6950 11550 7100 11600
rect 7150 11400 7300 11450
rect 7150 11380 7200 11400
rect 6060 11350 7200 11380
rect 7250 11350 7300 11400
rect 6060 11330 7300 11350
rect 7150 11300 7300 11330
rect 6120 11200 7300 11250
rect 7150 11150 7200 11200
rect 7250 11150 7300 11200
rect 7150 11100 7300 11150
rect 400 11000 600 11100
rect 400 10950 450 11000
rect 550 10950 600 11000
rect 400 10850 600 10950
<< via2 >>
rect 9400 12850 9450 12900
rect 6300 12550 6350 12600
rect 150 12250 250 12300
rect 7200 11350 7250 11400
rect 7200 11150 7250 11200
rect 450 10950 550 11000
<< metal3 >>
rect 9350 12900 9500 12950
rect 9350 12850 9400 12900
rect 9450 12850 9500 12900
rect 9350 12800 9500 12850
rect 6250 12600 6400 12650
rect 6250 12550 6300 12600
rect 6350 12550 6400 12600
rect 6250 12500 6400 12550
rect 100 12300 300 12400
rect 100 12250 150 12300
rect 250 12250 300 12300
rect 100 12150 300 12250
rect 7150 11400 7300 11450
rect 7150 11350 7200 11400
rect 7250 11350 7300 11400
rect 7150 11300 7300 11350
rect 7150 11200 15300 11250
rect 7150 11150 7200 11200
rect 7250 11150 15200 11200
rect 15250 11150 15300 11200
rect 7150 11100 15300 11150
rect 400 11000 600 11100
rect 400 10950 450 11000
rect 550 10950 600 11000
rect 400 10850 600 10950
<< via3 >>
rect 9400 12850 9450 12900
rect 6300 12550 6350 12600
rect 150 12250 250 12300
rect 7200 11350 7250 11400
rect 15200 11150 15250 11200
rect 450 10950 550 11000
<< metal4 >>
rect 3067 22476 3097 22576
rect 3343 22476 3373 22576
rect 3619 22476 3649 22576
rect 3895 22476 3925 22576
rect 4171 22476 4201 22576
rect 4447 22476 4477 22576
rect 4723 22476 4753 22576
rect 4999 22476 5029 22576
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22476 6961 22576
rect 7207 22476 7237 22576
rect 7483 22476 7513 22576
rect 7759 22476 7789 22576
rect 8035 22476 8065 22576
rect 8311 22476 8341 22576
rect 8587 22476 8617 22576
rect 8863 22476 8893 22576
rect 9139 22476 9169 22576
rect 9415 22500 9445 22576
rect 100 12300 300 22076
rect 100 12250 150 12300
rect 250 12250 300 12300
rect 100 500 300 12250
rect 400 11000 600 22076
rect 9350 12900 9500 22500
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22480 13861 22576
rect 13825 22450 13870 22480
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 9350 12850 9400 12900
rect 9450 12850 9500 12900
rect 9350 12800 9500 12850
rect 13750 12650 13900 22450
rect 6250 12600 13900 12650
rect 6250 12550 6300 12600
rect 6350 12550 13900 12600
rect 6250 12500 13900 12550
rect 7150 11400 13350 11450
rect 7150 11350 7200 11400
rect 7250 11350 13350 11400
rect 7150 11300 13350 11350
rect 400 10950 450 11000
rect 550 10950 600 11000
rect 400 500 600 10950
rect 13200 100 13350 11300
rect 15150 11200 15300 11250
rect 15150 11150 15200 11200
rect 15250 11150 15300 11200
rect 15150 100 15300 11150
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13249 0 13339 100
rect 15181 0 15271 100
use FAMILY  FAMILY_0 ~/dev/personal/chacha-silicon/tt09-analog-switch
timestamp 1730992266
transform 1 0 2000 0 1 1000
box 0 0 9990 7500
use SWTCH_UNIT  SWTCH_UNIT_0 ~/dev/personal/chacha-silicon/tt09-analog-switch/swtch_unit_sky130nm/design/SWTCH_UNIT_SKY130NM
timestamp 1730751262
transform 1 0 6000 0 1 11600
box 0 -600 697 610
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 100 500 300 22076 1 FreeSans 1 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 1 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
