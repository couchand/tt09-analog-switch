magic
tech sky130A
timestamp 1730992266
<< locali >>
rect 2270 7490 3340 7500
rect 3560 7490 3680 7500
rect 2250 7480 2260 7490
rect 2270 7480 3330 7490
rect 3570 7480 3680 7490
rect 9920 7480 9960 7490
rect 2220 7470 3330 7480
rect 3570 7470 3670 7480
rect 9840 7470 9940 7480
rect 2220 7460 3330 7470
rect 3570 7460 3660 7470
rect 9820 7460 9850 7470
rect 9860 7460 9930 7470
rect 2210 7450 3330 7460
rect 3580 7450 3660 7460
rect 9820 7450 9850 7460
rect 9870 7450 9920 7460
rect 2190 7440 3330 7450
rect 3580 7440 3660 7450
rect 9810 7440 9920 7450
rect 2190 7430 3330 7440
rect 3600 7430 3660 7440
rect 9790 7430 9910 7440
rect 2170 7420 3330 7430
rect 3580 7420 3640 7430
rect 9770 7420 9910 7430
rect 2150 7410 3330 7420
rect 3590 7410 3640 7420
rect 9750 7410 9890 7420
rect 2140 7400 3330 7410
rect 3600 7400 3620 7410
rect 3630 7400 3640 7410
rect 9710 7400 9890 7410
rect 2140 7390 3330 7400
rect 9690 7390 9860 7400
rect 2130 7380 2140 7390
rect 2150 7380 3330 7390
rect 9670 7380 9710 7390
rect 9750 7380 9800 7390
rect 2130 7370 3340 7380
rect 9650 7370 9690 7380
rect 2110 7360 3350 7370
rect 9650 7360 9680 7370
rect 2110 7350 3340 7360
rect 9650 7350 9670 7360
rect 2090 7340 3350 7350
rect 9650 7340 9670 7350
rect 2080 7330 3340 7340
rect 9650 7330 9670 7340
rect 9790 7330 9800 7340
rect 9880 7330 9890 7340
rect 2080 7320 3340 7330
rect 9770 7320 9780 7330
rect 9790 7320 9800 7330
rect 2080 7310 3340 7320
rect 9770 7310 9800 7320
rect 2070 7300 2080 7310
rect 2090 7300 3330 7310
rect 2070 7290 2530 7300
rect 2540 7290 3350 7300
rect 2060 7280 2530 7290
rect 2550 7280 3330 7290
rect 2050 7270 2380 7280
rect 2390 7270 2520 7280
rect 2590 7270 3340 7280
rect 2050 7260 2520 7270
rect 2570 7260 3320 7270
rect 3360 7260 3370 7270
rect 2050 7250 2510 7260
rect 2560 7250 3320 7260
rect 3330 7250 3340 7260
rect 2030 7240 2340 7250
rect 2350 7240 2440 7250
rect 2460 7240 2500 7250
rect 2570 7240 3330 7250
rect 2020 7230 2320 7240
rect 2330 7230 2430 7240
rect 2460 7230 2500 7240
rect 2540 7230 3350 7240
rect 2030 7220 2320 7230
rect 2330 7220 2410 7230
rect 2460 7220 2490 7230
rect 2500 7220 2510 7230
rect 2530 7220 3350 7230
rect 3370 7220 3380 7230
rect 2020 7210 2410 7220
rect 2450 7210 2490 7220
rect 2500 7210 3350 7220
rect 3360 7210 3390 7220
rect 2020 7200 2190 7210
rect 2200 7200 2210 7210
rect 2220 7200 2260 7210
rect 2270 7200 2400 7210
rect 2440 7200 3340 7210
rect 3360 7200 3370 7210
rect 3430 7200 3440 7210
rect 9860 7200 9880 7210
rect 2010 7190 2140 7200
rect 2170 7190 2190 7200
rect 2200 7190 2220 7200
rect 2230 7190 2240 7200
rect 2250 7190 2260 7200
rect 2270 7190 2290 7200
rect 2300 7190 2330 7200
rect 2420 7190 3310 7200
rect 3440 7190 3450 7200
rect 9850 7190 9890 7200
rect 2000 7180 2130 7190
rect 2210 7180 2220 7190
rect 2300 7180 2310 7190
rect 2340 7180 2370 7190
rect 2390 7180 3340 7190
rect 3440 7180 3450 7190
rect 9850 7180 9890 7190
rect 2000 7170 2110 7180
rect 2120 7170 2130 7180
rect 2330 7170 3350 7180
rect 9850 7170 9900 7180
rect 2000 7160 2110 7170
rect 2280 7160 2290 7170
rect 2320 7160 3350 7170
rect 1990 7150 2100 7160
rect 2260 7150 2270 7160
rect 2280 7150 3350 7160
rect 1980 7140 2090 7150
rect 2260 7140 3360 7150
rect 9880 7140 9900 7150
rect 1990 7130 2080 7140
rect 2230 7130 3370 7140
rect 9860 7130 9920 7140
rect 1980 7120 2060 7130
rect 2210 7120 3410 7130
rect 9860 7120 9920 7130
rect 1980 7110 2040 7120
rect 2200 7110 3460 7120
rect 9850 7110 9930 7120
rect 1990 7100 2030 7110
rect 2160 7100 3420 7110
rect 9850 7100 9940 7110
rect 2000 7090 2020 7100
rect 2040 7090 2060 7100
rect 2140 7090 2260 7100
rect 2280 7090 3420 7100
rect 9840 7090 9950 7100
rect 9990 7090 9990 7100
rect 2140 7080 3410 7090
rect 9840 7080 9960 7090
rect 9980 7080 9990 7090
rect 2130 7070 2170 7080
rect 2180 7070 3440 7080
rect 9830 7070 9990 7080
rect 2100 7060 2170 7070
rect 2190 7060 3390 7070
rect 3400 7060 3430 7070
rect 9830 7060 9990 7070
rect 2100 7050 2290 7060
rect 2360 7050 3440 7060
rect 9810 7050 9980 7060
rect 2090 7040 2240 7050
rect 2380 7040 2520 7050
rect 2540 7040 2560 7050
rect 2810 7040 2840 7050
rect 2850 7040 3440 7050
rect 3470 7040 3480 7050
rect 3510 7040 3520 7050
rect 9800 7040 9950 7050
rect 2070 7030 2220 7040
rect 2410 7030 2450 7040
rect 2480 7030 2490 7040
rect 3030 7030 3170 7040
rect 3180 7030 3470 7040
rect 3490 7030 3500 7040
rect 9790 7030 9930 7040
rect 2070 7020 2200 7030
rect 2420 7020 2450 7030
rect 3090 7020 3480 7030
rect 9780 7020 9920 7030
rect 2050 7010 2200 7020
rect 3130 7010 3470 7020
rect 9770 7010 9910 7020
rect 2050 7000 2180 7010
rect 3180 7000 3470 7010
rect 9720 7000 9840 7010
rect 9860 7000 9890 7010
rect 9980 7000 9990 7010
rect 2020 6990 2030 7000
rect 2040 6990 2170 7000
rect 3210 6990 3480 7000
rect 9690 6990 9810 7000
rect 9920 6990 9960 7000
rect 9970 6990 9990 7000
rect 2010 6980 2180 6990
rect 3240 6980 3490 6990
rect 9670 6980 9780 6990
rect 9880 6980 9990 6990
rect 1990 6970 2180 6980
rect 3280 6970 3500 6980
rect 9670 6970 9760 6980
rect 9870 6970 9990 6980
rect 1990 6960 2180 6970
rect 3300 6960 3510 6970
rect 9670 6960 9740 6970
rect 9860 6960 9990 6970
rect 1990 6950 2190 6960
rect 3330 6950 3520 6960
rect 9660 6950 9720 6960
rect 9850 6950 9990 6960
rect 1950 6940 2190 6950
rect 3360 6940 3530 6950
rect 9660 6940 9710 6950
rect 9840 6940 9990 6950
rect 1950 6930 2200 6940
rect 3380 6930 3550 6940
rect 9660 6930 9680 6940
rect 9840 6930 9990 6940
rect 1940 6920 2210 6930
rect 3410 6920 3560 6930
rect 9660 6920 9680 6930
rect 9840 6920 9990 6930
rect 1930 6910 2220 6920
rect 3430 6910 3590 6920
rect 9840 6910 9990 6920
rect 1910 6900 2230 6910
rect 3450 6900 3520 6910
rect 3530 6900 3600 6910
rect 9850 6900 9990 6910
rect 1900 6890 2250 6900
rect 3480 6890 3530 6900
rect 3540 6890 3620 6900
rect 9850 6890 9990 6900
rect 1900 6880 2260 6890
rect 3500 6880 3630 6890
rect 9850 6880 9990 6890
rect 1900 6870 2260 6880
rect 3520 6870 3570 6880
rect 3580 6870 3650 6880
rect 9860 6870 9990 6880
rect 1940 6860 2280 6870
rect 3540 6860 3580 6870
rect 3600 6860 3670 6870
rect 9860 6860 9950 6870
rect 9980 6860 9990 6870
rect 1910 6850 2290 6860
rect 3560 6850 3680 6860
rect 9860 6850 9940 6860
rect 9990 6850 9990 6860
rect 1900 6840 2300 6850
rect 3570 6840 3610 6850
rect 3630 6840 3690 6850
rect 9870 6840 9920 6850
rect 9990 6840 9990 6850
rect 1900 6830 2330 6840
rect 3590 6830 3700 6840
rect 9870 6830 9930 6840
rect 9990 6830 9990 6840
rect 1900 6820 2350 6830
rect 3610 6820 3650 6830
rect 3660 6820 3710 6830
rect 9860 6820 9910 6830
rect 9990 6820 9990 6830
rect 1900 6810 2370 6820
rect 3630 6810 3670 6820
rect 3680 6810 3730 6820
rect 9860 6810 9920 6820
rect 9990 6810 9990 6820
rect 1890 6800 1950 6810
rect 1970 6800 2390 6810
rect 3640 6800 3740 6810
rect 9870 6800 9920 6810
rect 1900 6790 1940 6800
rect 1960 6790 1980 6800
rect 2020 6790 2290 6800
rect 2360 6790 2410 6800
rect 3660 6790 3680 6800
rect 3710 6790 3760 6800
rect 9860 6790 9920 6800
rect 1900 6780 1920 6790
rect 1940 6780 1960 6790
rect 2030 6780 2270 6790
rect 2370 6780 2460 6790
rect 3670 6780 3770 6790
rect 9860 6780 9930 6790
rect 1910 6770 1960 6780
rect 2040 6770 2260 6780
rect 2390 6770 2500 6780
rect 3690 6770 3710 6780
rect 3730 6770 3780 6780
rect 9860 6770 9940 6780
rect 1910 6760 1960 6770
rect 2040 6760 2250 6770
rect 2410 6760 2530 6770
rect 2570 6760 2650 6770
rect 3700 6760 3720 6770
rect 3740 6760 3790 6770
rect 9850 6760 9950 6770
rect 1900 6750 1950 6760
rect 1990 6750 2030 6760
rect 2060 6750 2260 6760
rect 2430 6750 2730 6760
rect 3720 6750 3740 6760
rect 3750 6750 3800 6760
rect 9840 6750 9960 6760
rect 1910 6740 1940 6750
rect 1990 6740 2250 6750
rect 2450 6740 2820 6750
rect 3730 6740 3750 6750
rect 3770 6740 3810 6750
rect 9840 6740 9990 6750
rect 1980 6730 2240 6740
rect 2470 6730 2900 6740
rect 3740 6730 3770 6740
rect 3780 6730 3830 6740
rect 9840 6730 9990 6740
rect 1980 6720 2230 6730
rect 2490 6720 3030 6730
rect 3760 6720 3780 6730
rect 3790 6720 3840 6730
rect 9550 6720 9560 6730
rect 9850 6720 9990 6730
rect 1980 6710 2230 6720
rect 2520 6710 3100 6720
rect 3770 6710 3780 6720
rect 3800 6710 3850 6720
rect 9540 6710 9560 6720
rect 9850 6710 9990 6720
rect 1950 6700 1960 6710
rect 1980 6700 2220 6710
rect 2550 6700 3200 6710
rect 3780 6700 3800 6710
rect 3810 6700 3860 6710
rect 9550 6700 9560 6710
rect 9840 6700 9990 6710
rect 1960 6690 2220 6700
rect 2580 6690 3230 6700
rect 3790 6690 3810 6700
rect 3830 6690 3870 6700
rect 9840 6690 9980 6700
rect 1970 6680 2220 6690
rect 2630 6680 3320 6690
rect 3810 6680 3820 6690
rect 3830 6680 3880 6690
rect 9710 6680 9720 6690
rect 9830 6680 9950 6690
rect 1930 6670 1950 6680
rect 1960 6670 2230 6680
rect 2670 6670 3370 6680
rect 3850 6670 3890 6680
rect 9820 6670 9920 6680
rect 1930 6660 2220 6670
rect 2660 6660 3420 6670
rect 3850 6660 3900 6670
rect 9810 6660 9890 6670
rect 1900 6650 1930 6660
rect 1940 6650 2210 6660
rect 2650 6650 3470 6660
rect 3840 6650 3850 6660
rect 3860 6650 3910 6660
rect 9710 6650 9720 6660
rect 9780 6650 9850 6660
rect 1860 6640 2200 6650
rect 2660 6640 3500 6650
rect 3870 6640 3910 6650
rect 9710 6640 9820 6650
rect 1890 6630 2190 6640
rect 2650 6630 3530 6640
rect 3860 6630 3920 6640
rect 9710 6630 9760 6640
rect 9770 6630 9800 6640
rect 1780 6620 1810 6630
rect 1840 6620 2180 6630
rect 2650 6620 3560 6630
rect 3880 6620 3930 6630
rect 9700 6620 9750 6630
rect 1800 6610 2170 6620
rect 2660 6610 3590 6620
rect 3890 6610 3930 6620
rect 9700 6610 9730 6620
rect 1620 6600 1630 6610
rect 1770 6600 2160 6610
rect 2660 6600 3620 6610
rect 3900 6600 3940 6610
rect 9700 6600 9710 6610
rect 1610 6590 1620 6600
rect 1770 6590 2130 6600
rect 2660 6590 3640 6600
rect 3910 6590 3940 6600
rect 1580 6580 1610 6590
rect 1790 6580 2070 6590
rect 2100 6580 2130 6590
rect 2670 6580 3670 6590
rect 3910 6580 3950 6590
rect 1570 6570 1600 6580
rect 1800 6570 2070 6580
rect 2660 6570 3710 6580
rect 3920 6570 3960 6580
rect 1550 6560 1590 6570
rect 1810 6560 1990 6570
rect 2680 6560 3720 6570
rect 3930 6560 3960 6570
rect 1530 6550 1580 6560
rect 1820 6550 2000 6560
rect 2670 6550 3750 6560
rect 3940 6550 3970 6560
rect 1510 6540 1580 6550
rect 1690 6540 1710 6550
rect 1830 6540 2010 6550
rect 2680 6540 3760 6550
rect 3940 6540 3980 6550
rect 1450 6530 1470 6540
rect 1510 6530 1570 6540
rect 1620 6530 1740 6540
rect 1840 6530 2030 6540
rect 2690 6530 3780 6540
rect 3950 6530 3980 6540
rect 1490 6520 1570 6530
rect 1610 6520 1730 6530
rect 1850 6520 2040 6530
rect 2610 6520 3810 6530
rect 3960 6520 3980 6530
rect 1390 6510 1420 6520
rect 1490 6510 1570 6520
rect 1600 6510 1730 6520
rect 1850 6510 2060 6520
rect 2570 6510 3830 6520
rect 3970 6510 3990 6520
rect 9990 6510 9990 6520
rect 1310 6500 1330 6510
rect 1380 6500 1450 6510
rect 1470 6500 1550 6510
rect 1590 6500 1720 6510
rect 1860 6500 2080 6510
rect 2550 6500 3850 6510
rect 3970 6500 3990 6510
rect 9980 6500 9990 6510
rect 1310 6490 1330 6500
rect 1370 6490 1540 6500
rect 1590 6490 1690 6500
rect 1890 6490 2100 6500
rect 2550 6490 3870 6500
rect 3980 6490 4000 6500
rect 9980 6490 9990 6500
rect 1290 6480 1300 6490
rect 1310 6480 1330 6490
rect 1380 6480 1430 6490
rect 1440 6480 1550 6490
rect 1580 6480 1680 6490
rect 1890 6480 2100 6490
rect 2410 6480 2430 6490
rect 2550 6480 3880 6490
rect 3990 6480 4000 6490
rect 9890 6480 9910 6490
rect 9970 6480 9990 6490
rect 1280 6470 1320 6480
rect 1420 6470 1440 6480
rect 1450 6470 1560 6480
rect 1590 6470 1660 6480
rect 1900 6470 1920 6480
rect 1950 6470 2120 6480
rect 2410 6470 2430 6480
rect 2510 6470 2530 6480
rect 2570 6470 3900 6480
rect 4000 6470 4010 6480
rect 9880 6470 9930 6480
rect 9960 6470 9990 6480
rect 1260 6460 1310 6470
rect 1390 6460 1400 6470
rect 1410 6460 1550 6470
rect 1580 6460 1620 6470
rect 1910 6460 1920 6470
rect 1960 6460 2100 6470
rect 2400 6460 2430 6470
rect 2500 6460 2520 6470
rect 2570 6460 3920 6470
rect 9880 6460 9930 6470
rect 9970 6460 9990 6470
rect 1250 6450 1300 6460
rect 1380 6450 1550 6460
rect 1580 6450 1620 6460
rect 2400 6450 2430 6460
rect 2440 6450 2470 6460
rect 2490 6450 2510 6460
rect 2560 6450 3940 6460
rect 9870 6450 9930 6460
rect 9980 6450 9990 6460
rect 1260 6440 1290 6450
rect 1380 6440 1440 6450
rect 1460 6440 1550 6450
rect 1580 6440 1590 6450
rect 2390 6440 2490 6450
rect 2550 6440 3950 6450
rect 9800 6440 9930 6450
rect 9980 6440 9990 6450
rect 1250 6430 1280 6440
rect 1380 6430 1420 6440
rect 1470 6430 1550 6440
rect 2390 6430 2410 6440
rect 2430 6430 2500 6440
rect 2530 6430 3970 6440
rect 6470 6430 6480 6440
rect 9800 6430 9930 6440
rect 9990 6430 9990 6440
rect 1250 6420 1280 6430
rect 1400 6420 1420 6430
rect 1470 6420 1550 6430
rect 2380 6420 2410 6430
rect 2430 6420 2490 6430
rect 2520 6420 3980 6430
rect 6450 6420 6490 6430
rect 9760 6420 9770 6430
rect 9780 6420 9930 6430
rect 1250 6410 1270 6420
rect 1400 6410 1420 6420
rect 1490 6410 1550 6420
rect 2380 6410 2500 6420
rect 2520 6410 4000 6420
rect 6450 6410 6490 6420
rect 9770 6410 9930 6420
rect 1400 6400 1410 6410
rect 1490 6400 1550 6410
rect 2380 6400 2400 6410
rect 2410 6400 2490 6410
rect 2510 6400 4020 6410
rect 6460 6400 6500 6410
rect 9720 6400 9730 6410
rect 9750 6400 9930 6410
rect 1470 6390 1550 6400
rect 2400 6390 2410 6400
rect 2420 6390 4030 6400
rect 6470 6390 6490 6400
rect 9690 6390 9720 6400
rect 9750 6390 9760 6400
rect 9810 6390 9920 6400
rect 1470 6380 1550 6390
rect 2410 6380 2470 6390
rect 2480 6380 4040 6390
rect 9700 6380 9710 6390
rect 9830 6380 9930 6390
rect 1470 6370 1550 6380
rect 1780 6370 1820 6380
rect 2410 6370 2460 6380
rect 2480 6370 4060 6380
rect 9850 6370 9930 6380
rect 9990 6370 9990 6380
rect 1480 6360 1550 6370
rect 1760 6360 1830 6370
rect 2420 6360 2460 6370
rect 2480 6360 4070 6370
rect 9710 6360 9740 6370
rect 9860 6360 9940 6370
rect 1480 6350 1550 6360
rect 1750 6350 1830 6360
rect 2420 6350 4080 6360
rect 9690 6350 9740 6360
rect 9860 6350 9960 6360
rect 1470 6340 1560 6350
rect 1740 6340 1830 6350
rect 2420 6340 2450 6350
rect 2480 6340 4100 6350
rect 9680 6340 9740 6350
rect 9850 6340 9960 6350
rect 1460 6330 1560 6340
rect 1740 6330 1830 6340
rect 2430 6330 2450 6340
rect 2480 6330 4110 6340
rect 9710 6330 9740 6340
rect 9840 6330 9940 6340
rect 1450 6320 1560 6330
rect 1730 6320 1830 6330
rect 2430 6320 2450 6330
rect 2480 6320 4120 6330
rect 9690 6320 9740 6330
rect 9830 6320 9940 6330
rect 1450 6310 1560 6320
rect 1730 6310 1800 6320
rect 2430 6310 2440 6320
rect 2470 6310 4120 6320
rect 9690 6310 9790 6320
rect 9800 6310 9950 6320
rect 1430 6300 1560 6310
rect 1720 6300 1780 6310
rect 2430 6300 2440 6310
rect 2470 6300 4140 6310
rect 5430 6300 5470 6310
rect 9700 6300 9940 6310
rect 1420 6290 1570 6300
rect 1720 6290 1760 6300
rect 2430 6290 2440 6300
rect 2470 6290 4150 6300
rect 5450 6290 5500 6300
rect 9700 6290 9820 6300
rect 9890 6290 9930 6300
rect 1410 6280 1540 6290
rect 1550 6280 1570 6290
rect 1710 6280 1760 6290
rect 2430 6280 2440 6290
rect 2470 6280 4160 6290
rect 5410 6280 5520 6290
rect 9680 6280 9810 6290
rect 1420 6270 1530 6280
rect 1560 6270 1570 6280
rect 1700 6270 1750 6280
rect 2430 6270 2440 6280
rect 2460 6270 4170 6280
rect 5390 6270 5520 6280
rect 6710 6270 6740 6280
rect 9680 6270 9810 6280
rect 1420 6260 1520 6270
rect 1690 6260 1740 6270
rect 2430 6260 2440 6270
rect 2460 6260 4180 6270
rect 5390 6260 5400 6270
rect 5420 6260 5510 6270
rect 6710 6260 6740 6270
rect 9680 6260 9810 6270
rect 1420 6250 1560 6260
rect 1680 6250 1740 6260
rect 2430 6250 2440 6260
rect 2460 6250 4190 6260
rect 5420 6250 5500 6260
rect 6720 6250 6740 6260
rect 9650 6250 9660 6260
rect 9680 6250 9810 6260
rect 1420 6240 1570 6250
rect 1660 6240 1730 6250
rect 2430 6240 2440 6250
rect 2460 6240 4200 6250
rect 5340 6240 5360 6250
rect 5400 6240 5490 6250
rect 9530 6240 9600 6250
rect 9690 6240 9800 6250
rect 1420 6230 1560 6240
rect 1660 6230 1710 6240
rect 2430 6230 2440 6240
rect 2460 6230 4210 6240
rect 5330 6230 5340 6240
rect 5380 6230 5480 6240
rect 9510 6230 9520 6240
rect 9530 6230 9600 6240
rect 9680 6230 9800 6240
rect 1420 6220 1570 6230
rect 1660 6220 1700 6230
rect 2430 6220 2440 6230
rect 2460 6220 4220 6230
rect 5320 6220 5330 6230
rect 5370 6220 5470 6230
rect 9490 6220 9500 6230
rect 9520 6220 9540 6230
rect 9550 6220 9600 6230
rect 9630 6220 9640 6230
rect 9680 6220 9790 6230
rect 1430 6210 1570 6220
rect 1670 6210 1690 6220
rect 2430 6210 2440 6220
rect 2460 6210 4230 6220
rect 5360 6210 5390 6220
rect 5400 6210 5460 6220
rect 9450 6210 9480 6220
rect 9500 6210 9520 6220
rect 9530 6210 9600 6220
rect 9700 6210 9790 6220
rect 1420 6200 1570 6210
rect 1660 6200 1700 6210
rect 2430 6200 2450 6210
rect 2460 6200 4240 6210
rect 5350 6200 5380 6210
rect 5390 6200 5440 6210
rect 9410 6200 9600 6210
rect 9690 6200 9780 6210
rect 1420 6190 1570 6200
rect 1670 6190 1690 6200
rect 2430 6190 2450 6200
rect 2460 6190 4250 6200
rect 5340 6190 5440 6200
rect 9430 6190 9600 6200
rect 9690 6190 9780 6200
rect 1430 6180 1580 6190
rect 1680 6180 1690 6190
rect 2430 6180 4250 6190
rect 5330 6180 5430 6190
rect 9400 6180 9420 6190
rect 9430 6180 9600 6190
rect 9700 6180 9780 6190
rect 1430 6170 1580 6180
rect 2430 6170 4260 6180
rect 5320 6170 5420 6180
rect 9430 6170 9600 6180
rect 9700 6170 9790 6180
rect 1430 6160 1600 6170
rect 2430 6160 4260 6170
rect 5310 6160 5420 6170
rect 9340 6160 9350 6170
rect 9440 6160 9450 6170
rect 9460 6160 9600 6170
rect 9690 6160 9790 6170
rect 1430 6150 1600 6160
rect 2430 6150 2450 6160
rect 2460 6150 4270 6160
rect 5310 6150 5410 6160
rect 9470 6150 9610 6160
rect 9690 6150 9790 6160
rect 1440 6140 1610 6150
rect 2430 6140 4280 6150
rect 5300 6140 5400 6150
rect 9480 6140 9610 6150
rect 9690 6140 9800 6150
rect 1440 6130 1620 6140
rect 2440 6130 4280 6140
rect 5300 6130 5400 6140
rect 9280 6130 9300 6140
rect 9480 6130 9490 6140
rect 9500 6130 9630 6140
rect 9690 6130 9820 6140
rect 1370 6120 1380 6130
rect 1450 6120 1630 6130
rect 2440 6120 4290 6130
rect 5290 6120 5390 6130
rect 9270 6120 9350 6130
rect 9470 6120 9640 6130
rect 9690 6120 9820 6130
rect 1370 6110 1380 6120
rect 1430 6110 1440 6120
rect 1450 6110 1630 6120
rect 2440 6110 3790 6120
rect 3800 6110 4300 6120
rect 5290 6110 5380 6120
rect 9270 6110 9360 6120
rect 9480 6110 9640 6120
rect 9700 6110 9830 6120
rect 1320 6100 1330 6110
rect 1370 6100 1390 6110
rect 1430 6100 1590 6110
rect 2450 6100 3790 6110
rect 3800 6100 3910 6110
rect 3940 6100 4300 6110
rect 5280 6100 5380 6110
rect 9240 6100 9390 6110
rect 9490 6100 9600 6110
rect 9610 6100 9640 6110
rect 9700 6100 9830 6110
rect 1320 6090 1340 6100
rect 1380 6090 1390 6100
rect 1430 6090 1590 6100
rect 2450 6090 2470 6100
rect 2480 6090 3790 6100
rect 3800 6090 3890 6100
rect 3960 6090 4310 6100
rect 5270 6090 5370 6100
rect 9250 6090 9360 6100
rect 9520 6090 9640 6100
rect 9700 6090 9850 6100
rect 1310 6080 1340 6090
rect 1390 6080 1400 6090
rect 1430 6080 1590 6090
rect 2450 6080 2470 6090
rect 2480 6080 3780 6090
rect 3800 6080 3880 6090
rect 3970 6080 4310 6090
rect 5270 6080 5360 6090
rect 9260 6080 9340 6090
rect 9520 6080 9640 6090
rect 9710 6080 9850 6090
rect 1310 6070 1320 6080
rect 1330 6070 1350 6080
rect 1380 6070 1410 6080
rect 1430 6070 1590 6080
rect 2460 6070 3780 6080
rect 3800 6070 3860 6080
rect 3970 6070 4320 6080
rect 5260 6070 5360 6080
rect 9220 6070 9240 6080
rect 9250 6070 9330 6080
rect 9530 6070 9640 6080
rect 9710 6070 9850 6080
rect 1340 6060 1350 6070
rect 1390 6060 1410 6070
rect 1430 6060 1600 6070
rect 2460 6060 2480 6070
rect 2490 6060 3240 6070
rect 3260 6060 3780 6070
rect 3800 6060 3820 6070
rect 3980 6060 4330 6070
rect 5260 6060 5360 6070
rect 9230 6060 9270 6070
rect 9530 6060 9630 6070
rect 9710 6060 9850 6070
rect 1320 6050 1330 6060
rect 1340 6050 1360 6060
rect 1380 6050 1410 6060
rect 1430 6050 1600 6060
rect 2460 6050 3230 6060
rect 3280 6050 3780 6060
rect 3990 6050 4330 6060
rect 5250 6050 5360 6060
rect 9530 6050 9640 6060
rect 9720 6050 9860 6060
rect 1340 6040 1360 6050
rect 1370 6040 1420 6050
rect 1430 6040 1610 6050
rect 2470 6040 2490 6050
rect 2500 6040 3220 6050
rect 3290 6040 3780 6050
rect 4000 6040 4330 6050
rect 5240 6040 5360 6050
rect 9520 6040 9640 6050
rect 9720 6040 9860 6050
rect 1330 6030 1420 6040
rect 1430 6030 1610 6040
rect 2470 6030 3210 6040
rect 3290 6030 3780 6040
rect 4010 6030 4340 6040
rect 5240 6030 5360 6040
rect 9520 6030 9650 6040
rect 9720 6030 9850 6040
rect 1210 6020 1220 6030
rect 1330 6020 1420 6030
rect 1430 6020 1610 6030
rect 2480 6020 3200 6030
rect 3290 6020 3790 6030
rect 4020 6020 4340 6030
rect 5240 6020 5360 6030
rect 9290 6020 9320 6030
rect 9520 6020 9650 6030
rect 9720 6020 9850 6030
rect 1220 6010 1230 6020
rect 1340 6010 1420 6020
rect 1430 6010 1620 6020
rect 2490 6010 3190 6020
rect 3290 6010 3790 6020
rect 4040 6010 4340 6020
rect 5230 6010 5350 6020
rect 9280 6010 9310 6020
rect 9500 6010 9600 6020
rect 9610 6010 9650 6020
rect 9720 6010 9850 6020
rect 1220 6000 1240 6010
rect 1340 6000 1420 6010
rect 1430 6000 1620 6010
rect 2490 6000 3180 6010
rect 3290 6000 3800 6010
rect 4050 6000 4340 6010
rect 5210 6000 5340 6010
rect 9300 6000 9310 6010
rect 9480 6000 9660 6010
rect 9720 6000 9870 6010
rect 860 5990 880 6000
rect 1230 5990 1250 6000
rect 1300 5990 1310 6000
rect 1340 5990 1420 6000
rect 1430 5990 1630 6000
rect 2500 5990 3170 6000
rect 3290 5990 3790 6000
rect 4060 5990 4340 6000
rect 5210 5990 5340 6000
rect 9470 5990 9670 6000
rect 9730 5990 9880 6000
rect 1220 5980 1250 5990
rect 1300 5980 1630 5990
rect 2510 5980 3160 5990
rect 3290 5980 3780 5990
rect 4080 5980 4340 5990
rect 5200 5980 5340 5990
rect 9310 5980 9320 5990
rect 9480 5980 9660 5990
rect 9730 5980 9890 5990
rect 1200 5970 1260 5980
rect 1290 5970 1640 5980
rect 1670 5970 1680 5980
rect 2520 5970 3160 5980
rect 3290 5970 3780 5980
rect 3840 5970 3850 5980
rect 4090 5970 4340 5980
rect 5190 5970 5340 5980
rect 9490 5970 9680 5980
rect 9740 5970 9890 5980
rect 1190 5960 1260 5970
rect 1280 5960 1670 5970
rect 2530 5960 3150 5970
rect 3290 5960 3770 5970
rect 4110 5960 4340 5970
rect 5180 5960 5340 5970
rect 9500 5960 9680 5970
rect 9740 5960 9880 5970
rect 1190 5950 1200 5960
rect 1210 5950 1260 5960
rect 1280 5950 1670 5960
rect 2540 5950 3140 5960
rect 3280 5950 3770 5960
rect 4130 5950 4340 5960
rect 5170 5950 5330 5960
rect 9310 5950 9320 5960
rect 9510 5950 9670 5960
rect 9740 5950 9890 5960
rect 990 5940 1000 5950
rect 1140 5940 1150 5950
rect 1190 5940 1260 5950
rect 1280 5940 1670 5950
rect 2550 5940 3130 5950
rect 3280 5940 3770 5950
rect 4150 5940 4330 5950
rect 5160 5940 5330 5950
rect 9300 5940 9320 5950
rect 9330 5940 9340 5950
rect 9520 5940 9690 5950
rect 9750 5940 9890 5950
rect 980 5930 1000 5940
rect 1130 5930 1160 5940
rect 1190 5930 1270 5940
rect 1280 5930 1670 5940
rect 2560 5930 3120 5940
rect 3280 5930 3760 5940
rect 4170 5930 4330 5940
rect 5160 5930 5330 5940
rect 9320 5930 9350 5940
rect 9520 5930 9690 5940
rect 9750 5930 9890 5940
rect 970 5920 1010 5930
rect 1020 5920 1030 5930
rect 1040 5920 1050 5930
rect 1070 5920 1210 5930
rect 1220 5920 1230 5930
rect 1240 5920 1680 5930
rect 2580 5920 3100 5930
rect 3280 5920 3760 5930
rect 4190 5920 4330 5930
rect 5150 5920 5330 5930
rect 6870 5920 6900 5930
rect 9310 5920 9320 5930
rect 9340 5920 9350 5930
rect 9510 5920 9700 5930
rect 9760 5920 9890 5930
rect 950 5910 1010 5920
rect 1060 5910 1210 5920
rect 1230 5910 1680 5920
rect 2590 5910 3090 5920
rect 3290 5910 3760 5920
rect 4210 5910 4320 5920
rect 5140 5910 5170 5920
rect 5180 5910 5330 5920
rect 6860 5910 6910 5920
rect 8730 5910 8750 5920
rect 9310 5910 9320 5920
rect 9350 5910 9360 5920
rect 9440 5910 9450 5920
rect 9470 5910 9710 5920
rect 9760 5910 9890 5920
rect 970 5900 1050 5910
rect 1070 5900 1130 5910
rect 1140 5900 1160 5910
rect 1180 5900 1190 5910
rect 1210 5900 1700 5910
rect 2610 5900 3070 5910
rect 3300 5900 3750 5910
rect 4230 5900 4280 5910
rect 5160 5900 5320 5910
rect 6860 5900 6910 5910
rect 8730 5900 8750 5910
rect 9350 5900 9360 5910
rect 9430 5900 9440 5910
rect 9460 5900 9720 5910
rect 9750 5900 9890 5910
rect 980 5890 1010 5900
rect 1070 5890 1100 5900
rect 1160 5890 1170 5900
rect 1200 5890 1710 5900
rect 2620 5890 3060 5900
rect 3290 5890 3750 5900
rect 5170 5890 5310 5900
rect 6850 5890 6910 5900
rect 9350 5890 9380 5900
rect 9420 5890 9720 5900
rect 9750 5890 9890 5900
rect 990 5880 1020 5890
rect 1130 5880 1720 5890
rect 2640 5880 3040 5890
rect 3290 5880 3740 5890
rect 5160 5880 5320 5890
rect 6850 5880 6910 5890
rect 9350 5880 9730 5890
rect 9750 5880 9900 5890
rect 990 5870 1040 5880
rect 1050 5870 1130 5880
rect 1140 5870 1740 5880
rect 2660 5870 2990 5880
rect 3290 5870 3740 5880
rect 5150 5870 5320 5880
rect 6850 5870 6910 5880
rect 9360 5870 9730 5880
rect 9740 5870 9910 5880
rect 1000 5860 1040 5870
rect 1050 5860 1750 5870
rect 1830 5860 1840 5870
rect 2690 5860 2980 5870
rect 3290 5860 3740 5870
rect 5130 5860 5310 5870
rect 6850 5860 6920 5870
rect 9360 5860 9910 5870
rect 990 5850 1840 5860
rect 2700 5850 2930 5860
rect 3290 5850 3730 5860
rect 5120 5850 5130 5860
rect 5140 5850 5310 5860
rect 6850 5850 6930 5860
rect 9320 5850 9900 5860
rect 860 5840 870 5850
rect 990 5840 1850 5850
rect 2710 5840 2890 5850
rect 3290 5840 3730 5850
rect 5130 5840 5310 5850
rect 6850 5840 6920 5850
rect 9340 5840 9900 5850
rect 820 5830 880 5840
rect 890 5830 910 5840
rect 950 5830 1850 5840
rect 2710 5830 2860 5840
rect 3290 5830 3730 5840
rect 5130 5830 5300 5840
rect 6840 5830 6920 5840
rect 9330 5830 9910 5840
rect 820 5820 1850 5830
rect 2740 5820 2840 5830
rect 3290 5820 3720 5830
rect 5120 5820 5300 5830
rect 6850 5820 6920 5830
rect 9310 5820 9920 5830
rect 820 5810 840 5820
rect 880 5810 1010 5820
rect 1020 5810 1850 5820
rect 3290 5810 3720 5820
rect 5120 5810 5300 5820
rect 6850 5810 6910 5820
rect 9300 5810 9930 5820
rect 820 5800 840 5810
rect 900 5800 1850 5810
rect 3290 5800 3740 5810
rect 3960 5800 3970 5810
rect 5110 5800 5300 5810
rect 6850 5800 6910 5810
rect 8750 5800 8760 5810
rect 9260 5800 9930 5810
rect 810 5790 830 5800
rect 910 5790 1850 5800
rect 3300 5790 3770 5800
rect 3820 5790 3830 5800
rect 5100 5790 5300 5800
rect 6850 5790 6910 5800
rect 6920 5790 6940 5800
rect 8740 5790 8750 5800
rect 9250 5790 9930 5800
rect 800 5780 810 5790
rect 910 5780 1850 5790
rect 3290 5780 3800 5790
rect 5100 5780 5300 5790
rect 6850 5780 6900 5790
rect 6920 5780 6940 5790
rect 9220 5780 9240 5790
rect 9250 5780 9930 5790
rect 790 5770 800 5780
rect 910 5770 1850 5780
rect 3300 5770 3780 5780
rect 5100 5770 5300 5780
rect 6860 5770 6910 5780
rect 6920 5770 6930 5780
rect 9090 5770 9160 5780
rect 9230 5770 9930 5780
rect 890 5760 1850 5770
rect 3300 5760 3770 5770
rect 5110 5760 5290 5770
rect 6870 5760 6930 5770
rect 8760 5760 8770 5770
rect 9070 5760 9180 5770
rect 9200 5760 9930 5770
rect 880 5750 1850 5760
rect 2710 5750 2740 5760
rect 3300 5750 3720 5760
rect 3890 5750 3910 5760
rect 5110 5750 5290 5760
rect 6900 5750 6930 5760
rect 8760 5750 8780 5760
rect 9070 5750 9930 5760
rect 880 5740 1850 5750
rect 2690 5740 2740 5750
rect 3300 5740 3720 5750
rect 3800 5740 3840 5750
rect 3920 5740 3930 5750
rect 5090 5740 5290 5750
rect 6930 5740 6950 5750
rect 8760 5740 8800 5750
rect 9040 5740 9930 5750
rect 870 5730 1850 5740
rect 2680 5730 2720 5740
rect 3310 5730 3700 5740
rect 3720 5730 3740 5740
rect 3840 5730 3880 5740
rect 3890 5730 3930 5740
rect 3990 5730 4000 5740
rect 5100 5730 5280 5740
rect 6930 5730 6950 5740
rect 8750 5730 8760 5740
rect 8770 5730 8800 5740
rect 9050 5730 9930 5740
rect 770 5720 1230 5730
rect 1250 5720 1860 5730
rect 2660 5720 2710 5730
rect 3320 5720 3700 5730
rect 3710 5720 3750 5730
rect 3850 5720 3960 5730
rect 3980 5720 4010 5730
rect 5100 5720 5130 5730
rect 5140 5720 5280 5730
rect 8750 5720 8810 5730
rect 9030 5720 9930 5730
rect 790 5710 1200 5720
rect 1240 5710 1860 5720
rect 2630 5710 2690 5720
rect 3310 5710 3720 5720
rect 3870 5710 4010 5720
rect 5100 5710 5110 5720
rect 5130 5710 5280 5720
rect 8600 5710 8610 5720
rect 8640 5710 8650 5720
rect 8750 5710 8830 5720
rect 8840 5710 8920 5720
rect 8930 5710 8940 5720
rect 8960 5710 8970 5720
rect 9040 5710 9930 5720
rect 810 5700 1160 5710
rect 1230 5700 1610 5710
rect 1620 5700 1860 5710
rect 2620 5700 2680 5710
rect 3320 5700 3670 5710
rect 3680 5700 3720 5710
rect 3780 5700 3800 5710
rect 3880 5700 4010 5710
rect 5130 5700 5280 5710
rect 8620 5700 8650 5710
rect 8760 5700 8950 5710
rect 9050 5700 9950 5710
rect 820 5690 1050 5700
rect 1060 5690 1120 5700
rect 1220 5690 1610 5700
rect 1620 5690 1860 5700
rect 2590 5690 2660 5700
rect 3310 5690 3670 5700
rect 3680 5690 3710 5700
rect 3770 5690 3800 5700
rect 3820 5690 3840 5700
rect 3900 5690 3910 5700
rect 3920 5690 4000 5700
rect 5150 5690 5280 5700
rect 6910 5690 6930 5700
rect 8630 5690 8650 5700
rect 8760 5690 8950 5700
rect 9040 5690 9950 5700
rect 840 5680 1040 5690
rect 1190 5680 1860 5690
rect 2590 5680 2650 5690
rect 3310 5680 3720 5690
rect 3770 5680 3780 5690
rect 3820 5680 3880 5690
rect 3940 5680 4000 5690
rect 5150 5680 5280 5690
rect 8570 5680 8600 5690
rect 8750 5680 8860 5690
rect 8870 5680 8880 5690
rect 8890 5680 8940 5690
rect 8990 5680 9990 5690
rect 840 5670 1150 5680
rect 1190 5670 1860 5680
rect 2590 5670 2630 5680
rect 3310 5670 3700 5680
rect 3710 5670 3720 5680
rect 3810 5670 3820 5680
rect 3840 5670 3850 5680
rect 3860 5670 3870 5680
rect 3890 5670 3900 5680
rect 3950 5670 3990 5680
rect 5150 5670 5270 5680
rect 8520 5670 8530 5680
rect 8580 5670 8620 5680
rect 8640 5670 8670 5680
rect 8740 5670 8880 5680
rect 8900 5670 8940 5680
rect 8990 5670 9990 5680
rect 830 5660 1860 5670
rect 2580 5660 2590 5670
rect 3310 5660 3660 5670
rect 3670 5660 3690 5670
rect 3770 5660 3780 5670
rect 3790 5660 3800 5670
rect 3840 5660 3870 5670
rect 3950 5660 3990 5670
rect 5140 5660 5270 5670
rect 6890 5660 6920 5670
rect 8560 5660 8650 5670
rect 8680 5660 8700 5670
rect 8710 5660 8720 5670
rect 8730 5660 8970 5670
rect 8980 5660 9990 5670
rect 820 5650 1870 5660
rect 2570 5650 2580 5660
rect 3310 5650 3660 5660
rect 3670 5650 3680 5660
rect 3770 5650 3790 5660
rect 3850 5650 3880 5660
rect 3920 5650 3980 5660
rect 5140 5650 5270 5660
rect 6880 5650 6930 5660
rect 8550 5650 8610 5660
rect 8620 5650 8670 5660
rect 8680 5650 9980 5660
rect 810 5640 1870 5650
rect 3300 5640 3700 5650
rect 3760 5640 3780 5650
rect 3830 5640 3850 5650
rect 3860 5640 3870 5650
rect 3920 5640 3930 5650
rect 5130 5640 5270 5650
rect 6880 5640 6940 5650
rect 8560 5640 8630 5650
rect 8640 5640 9980 5650
rect 790 5630 1860 5640
rect 3300 5630 3700 5640
rect 3750 5630 3770 5640
rect 3850 5630 3860 5640
rect 3910 5630 3920 5640
rect 5130 5630 5270 5640
rect 6890 5630 6940 5640
rect 8550 5630 8700 5640
rect 8710 5630 8720 5640
rect 8730 5630 8920 5640
rect 8940 5630 9960 5640
rect 760 5620 1860 5630
rect 3300 5620 3700 5630
rect 3740 5620 3790 5630
rect 5120 5620 5270 5630
rect 6890 5620 6940 5630
rect 8540 5620 8920 5630
rect 8950 5620 9960 5630
rect 740 5610 1860 5620
rect 3300 5610 3670 5620
rect 3720 5610 3790 5620
rect 5120 5610 5270 5620
rect 6890 5610 6940 5620
rect 8500 5610 8920 5620
rect 8950 5610 9960 5620
rect 720 5600 1860 5610
rect 3310 5600 3420 5610
rect 3430 5600 3650 5610
rect 3660 5600 3670 5610
rect 3710 5600 3790 5610
rect 5120 5600 5270 5610
rect 5670 5600 5700 5610
rect 6890 5600 6930 5610
rect 8460 5600 8950 5610
rect 8960 5600 8980 5610
rect 9070 5600 9960 5610
rect 720 5590 1870 5600
rect 3310 5590 3420 5600
rect 3440 5590 3650 5600
rect 3710 5590 3740 5600
rect 3760 5590 3770 5600
rect 5110 5590 5260 5600
rect 5640 5590 5780 5600
rect 6900 5590 6930 5600
rect 8430 5590 8940 5600
rect 8960 5590 8970 5600
rect 9080 5590 9970 5600
rect 690 5580 1860 5590
rect 3310 5580 3430 5590
rect 3450 5580 3650 5590
rect 3710 5580 3770 5590
rect 5120 5580 5260 5590
rect 5640 5580 5810 5590
rect 6900 5580 6930 5590
rect 8410 5580 8930 5590
rect 9090 5580 9980 5590
rect 690 5570 1870 5580
rect 3310 5570 3440 5580
rect 3460 5570 3640 5580
rect 3710 5570 3770 5580
rect 5110 5570 5260 5580
rect 5640 5570 5830 5580
rect 6900 5570 6920 5580
rect 8400 5570 8900 5580
rect 9100 5570 9990 5580
rect 680 5560 1870 5570
rect 3310 5560 3450 5570
rect 3470 5560 3640 5570
rect 3680 5560 3700 5570
rect 3710 5560 3730 5570
rect 5110 5560 5260 5570
rect 5630 5560 5850 5570
rect 6900 5560 6920 5570
rect 8330 5560 8340 5570
rect 8370 5560 8860 5570
rect 9100 5560 9990 5570
rect 670 5550 1870 5560
rect 2530 5550 2540 5560
rect 3310 5550 3460 5560
rect 3480 5550 3650 5560
rect 3710 5550 3720 5560
rect 5110 5550 5260 5560
rect 5680 5550 5850 5560
rect 6340 5550 6400 5560
rect 6910 5550 6930 5560
rect 8360 5550 8840 5560
rect 8850 5550 8860 5560
rect 9090 5550 9990 5560
rect 660 5540 1880 5550
rect 2490 5540 2500 5550
rect 3310 5540 3470 5550
rect 3500 5540 3650 5550
rect 3710 5540 3720 5550
rect 3770 5540 3780 5550
rect 5150 5540 5260 5550
rect 5760 5540 5860 5550
rect 6300 5540 6440 5550
rect 8300 5540 8780 5550
rect 8790 5540 8850 5550
rect 9050 5540 9060 5550
rect 9070 5540 9990 5550
rect 660 5530 930 5540
rect 960 5530 1890 5540
rect 1920 5530 1930 5540
rect 2480 5530 2530 5540
rect 3310 5530 3480 5540
rect 3510 5530 3650 5540
rect 3710 5530 3740 5540
rect 3760 5530 3770 5540
rect 5140 5530 5250 5540
rect 5810 5530 5850 5540
rect 6290 5530 6470 5540
rect 8230 5530 8240 5540
rect 8280 5530 8760 5540
rect 8810 5530 8840 5540
rect 9070 5530 9990 5540
rect 570 5520 590 5530
rect 650 5520 930 5530
rect 960 5520 1880 5530
rect 1920 5520 1930 5530
rect 2470 5520 2520 5530
rect 2540 5520 2550 5530
rect 2560 5520 2570 5530
rect 3310 5520 3500 5530
rect 3520 5520 3650 5530
rect 3710 5520 3730 5530
rect 5140 5520 5250 5530
rect 6270 5520 6480 5530
rect 8190 5520 8710 5530
rect 8740 5520 8750 5530
rect 9050 5520 9990 5530
rect 570 5510 580 5520
rect 650 5510 930 5520
rect 960 5510 1890 5520
rect 1920 5510 1930 5520
rect 2470 5510 2510 5520
rect 2540 5510 2550 5520
rect 3310 5510 3520 5520
rect 3540 5510 3650 5520
rect 3710 5510 3730 5520
rect 4160 5510 4180 5520
rect 5130 5510 5250 5520
rect 6260 5510 6460 5520
rect 8150 5510 8680 5520
rect 9030 5510 9060 5520
rect 9130 5510 9990 5520
rect 540 5500 570 5510
rect 640 5500 1890 5510
rect 1920 5500 1940 5510
rect 2460 5500 2480 5510
rect 3320 5500 3550 5510
rect 3570 5500 3650 5510
rect 5120 5500 5240 5510
rect 6250 5500 6370 5510
rect 7410 5500 7420 5510
rect 8150 5500 8160 5510
rect 8170 5500 8660 5510
rect 9130 5500 9990 5510
rect 450 5490 470 5500
rect 540 5490 570 5500
rect 640 5490 1890 5500
rect 1930 5490 1940 5500
rect 3320 5490 3590 5500
rect 3600 5490 3610 5500
rect 3630 5490 3660 5500
rect 5130 5490 5240 5500
rect 6240 5490 6350 5500
rect 7410 5490 7420 5500
rect 8150 5490 8610 5500
rect 9120 5490 9990 5500
rect 510 5480 550 5490
rect 630 5480 950 5490
rect 970 5480 1900 5490
rect 3330 5480 3550 5490
rect 3580 5480 3600 5490
rect 5120 5480 5240 5490
rect 6230 5480 6350 5490
rect 7410 5480 7420 5490
rect 8150 5480 8600 5490
rect 9130 5480 9990 5490
rect 490 5470 540 5480
rect 590 5470 610 5480
rect 620 5470 1900 5480
rect 2490 5470 2510 5480
rect 2530 5470 2540 5480
rect 3330 5470 3560 5480
rect 5120 5470 5240 5480
rect 5590 5470 5620 5480
rect 6240 5470 6350 5480
rect 8150 5470 8600 5480
rect 9130 5470 9990 5480
rect 460 5460 540 5470
rect 550 5460 560 5470
rect 590 5460 1900 5470
rect 2470 5460 2550 5470
rect 3330 5460 3570 5470
rect 5120 5460 5130 5470
rect 5140 5460 5240 5470
rect 5540 5460 5610 5470
rect 5660 5460 5750 5470
rect 6240 5460 6360 5470
rect 8150 5460 8520 5470
rect 8570 5460 8590 5470
rect 9130 5460 9990 5470
rect 460 5450 530 5460
rect 590 5450 1900 5460
rect 2460 5450 2550 5460
rect 3320 5450 3580 5460
rect 5140 5450 5240 5460
rect 5510 5450 5570 5460
rect 5690 5450 5770 5460
rect 6240 5450 6250 5460
rect 6270 5450 6360 5460
rect 8150 5450 8510 5460
rect 9020 5450 9030 5460
rect 9130 5450 9990 5460
rect 460 5440 520 5450
rect 590 5440 1910 5450
rect 1930 5440 1940 5450
rect 2440 5440 2540 5450
rect 2550 5440 2580 5450
rect 3320 5440 3580 5450
rect 5130 5440 5240 5450
rect 5490 5440 5540 5450
rect 5710 5440 5790 5450
rect 6240 5440 6360 5450
rect 8160 5440 8500 5450
rect 9030 5440 9040 5450
rect 9120 5440 9990 5450
rect 460 5430 510 5440
rect 580 5430 1910 5440
rect 2430 5430 2580 5440
rect 2600 5430 2620 5440
rect 3300 5430 3580 5440
rect 5130 5430 5240 5440
rect 5480 5430 5520 5440
rect 5740 5430 5800 5440
rect 6230 5430 6480 5440
rect 7470 5430 7480 5440
rect 7990 5430 8010 5440
rect 8160 5430 8430 5440
rect 8450 5430 8490 5440
rect 9120 5430 9550 5440
rect 9570 5430 9990 5440
rect 460 5420 500 5430
rect 580 5420 1920 5430
rect 2420 5420 2520 5430
rect 2530 5420 2610 5430
rect 3280 5420 3580 5430
rect 5120 5420 5230 5430
rect 5470 5420 5500 5430
rect 5580 5420 5700 5430
rect 5740 5420 5840 5430
rect 6230 5420 6530 5430
rect 7470 5420 7480 5430
rect 7980 5420 8010 5430
rect 8150 5420 8390 5430
rect 9120 5420 9550 5430
rect 9580 5420 9990 5430
rect 450 5410 500 5420
rect 580 5410 1920 5420
rect 2420 5410 2520 5420
rect 2530 5410 2600 5420
rect 2920 5410 2960 5420
rect 3270 5410 3570 5420
rect 5120 5410 5230 5420
rect 5460 5410 5490 5420
rect 5540 5410 5730 5420
rect 5750 5410 5860 5420
rect 6220 5410 6410 5420
rect 6430 5410 6560 5420
rect 8160 5410 8360 5420
rect 9100 5410 9480 5420
rect 9500 5410 9540 5420
rect 9590 5410 9990 5420
rect 440 5400 490 5410
rect 570 5400 760 5410
rect 780 5400 830 5410
rect 840 5400 890 5410
rect 950 5400 1920 5410
rect 2420 5400 2580 5410
rect 2910 5400 2990 5410
rect 3230 5400 3570 5410
rect 5110 5400 5230 5410
rect 5450 5400 5470 5410
rect 5520 5400 5870 5410
rect 6210 5400 6600 5410
rect 8150 5400 8340 5410
rect 9080 5400 9480 5410
rect 9520 5400 9540 5410
rect 9580 5400 9990 5410
rect 420 5390 500 5400
rect 570 5390 760 5400
rect 770 5390 820 5400
rect 830 5390 980 5400
rect 990 5390 1920 5400
rect 2420 5390 2580 5400
rect 2930 5390 3050 5400
rect 3210 5390 3570 5400
rect 5100 5390 5230 5400
rect 5440 5390 5460 5400
rect 5490 5390 5880 5400
rect 6210 5390 6620 5400
rect 8140 5390 8310 5400
rect 8320 5390 8340 5400
rect 8960 5390 8980 5400
rect 9050 5390 9410 5400
rect 9430 5390 9480 5400
rect 9580 5390 9990 5400
rect 400 5380 460 5390
rect 570 5380 1920 5390
rect 2430 5380 2480 5390
rect 2490 5380 2580 5390
rect 2950 5380 3080 5390
rect 3190 5380 3570 5390
rect 5100 5380 5230 5390
rect 5480 5380 5880 5390
rect 6210 5380 6630 5390
rect 8180 5380 8240 5390
rect 8950 5380 9400 5390
rect 9440 5380 9480 5390
rect 9580 5380 9990 5390
rect 380 5370 450 5380
rect 570 5370 880 5380
rect 920 5370 1920 5380
rect 2420 5370 2480 5380
rect 2490 5370 2580 5380
rect 3000 5370 3110 5380
rect 3170 5370 3490 5380
rect 3510 5370 3570 5380
rect 5100 5370 5130 5380
rect 5140 5370 5230 5380
rect 5460 5370 5720 5380
rect 5750 5370 5870 5380
rect 6200 5370 6650 5380
rect 7790 5370 7820 5380
rect 8180 5370 8220 5380
rect 8950 5370 9400 5380
rect 9450 5370 9490 5380
rect 9580 5370 9990 5380
rect 360 5360 440 5370
rect 550 5360 880 5370
rect 900 5360 1930 5370
rect 2420 5360 2480 5370
rect 2490 5360 2590 5370
rect 3010 5360 3490 5370
rect 3520 5360 3570 5370
rect 5100 5360 5130 5370
rect 5140 5360 5230 5370
rect 5440 5360 5720 5370
rect 5760 5360 5820 5370
rect 6200 5360 6550 5370
rect 6560 5360 6660 5370
rect 7780 5360 7830 5370
rect 8180 5360 8210 5370
rect 8870 5360 8880 5370
rect 8940 5360 9290 5370
rect 9360 5360 9400 5370
rect 9450 5360 9500 5370
rect 9580 5360 9990 5370
rect 350 5350 400 5360
rect 550 5350 880 5360
rect 900 5350 1930 5360
rect 2420 5350 2460 5360
rect 2510 5350 2600 5360
rect 3020 5350 3490 5360
rect 3520 5350 3560 5360
rect 5100 5350 5220 5360
rect 5430 5350 5460 5360
rect 5570 5350 5580 5360
rect 5590 5350 5600 5360
rect 5650 5350 5710 5360
rect 5750 5350 5830 5360
rect 6200 5350 6370 5360
rect 6390 5350 6540 5360
rect 6570 5350 6680 5360
rect 7760 5350 7840 5360
rect 8180 5350 8200 5360
rect 8850 5350 9270 5360
rect 9370 5350 9400 5360
rect 9450 5350 9510 5360
rect 9580 5350 9990 5360
rect 330 5340 360 5350
rect 560 5340 1930 5350
rect 2420 5340 2460 5350
rect 2520 5340 2600 5350
rect 3030 5340 3490 5350
rect 3510 5340 3560 5350
rect 5090 5340 5140 5350
rect 5150 5340 5220 5350
rect 5750 5340 5840 5350
rect 6210 5340 6280 5350
rect 6300 5340 6360 5350
rect 6390 5340 6540 5350
rect 6570 5340 6690 5350
rect 7720 5340 7740 5350
rect 7750 5340 7840 5350
rect 8490 5340 8510 5350
rect 8850 5340 9270 5350
rect 9380 5340 9410 5350
rect 9450 5340 9520 5350
rect 9580 5340 9990 5350
rect 290 5330 320 5340
rect 570 5330 1930 5340
rect 2420 5330 2450 5340
rect 2530 5330 2590 5340
rect 3050 5330 3480 5340
rect 3500 5330 3560 5340
rect 5130 5330 5140 5340
rect 5160 5330 5220 5340
rect 5770 5330 5850 5340
rect 6210 5330 6250 5340
rect 6290 5330 6350 5340
rect 6400 5330 6690 5340
rect 7480 5330 7490 5340
rect 7730 5330 7840 5340
rect 8480 5330 8510 5340
rect 8830 5330 9260 5340
rect 9370 5330 9410 5340
rect 9460 5330 9520 5340
rect 9590 5330 9990 5340
rect 270 5320 300 5330
rect 580 5320 1930 5330
rect 2430 5320 2440 5330
rect 2540 5320 2590 5330
rect 2790 5320 2800 5330
rect 3050 5320 3550 5330
rect 5170 5320 5210 5330
rect 5840 5320 5850 5330
rect 6220 5320 6240 5330
rect 6290 5320 6340 5330
rect 6400 5320 6700 5330
rect 7700 5320 7840 5330
rect 8490 5320 8520 5330
rect 8790 5320 9260 5330
rect 9330 5320 9420 5330
rect 9460 5320 9520 5330
rect 9600 5320 9990 5330
rect 590 5310 1940 5320
rect 2550 5310 2590 5320
rect 2810 5310 2830 5320
rect 3050 5310 3550 5320
rect 5170 5310 5180 5320
rect 5190 5310 5200 5320
rect 6280 5310 6370 5320
rect 6510 5310 6560 5320
rect 6660 5310 6720 5320
rect 7640 5310 7650 5320
rect 7670 5310 7690 5320
rect 7700 5310 7830 5320
rect 8480 5310 8520 5320
rect 8790 5310 9120 5320
rect 9150 5310 9250 5320
rect 9300 5310 9310 5320
rect 9320 5310 9420 5320
rect 9460 5310 9520 5320
rect 9610 5310 9990 5320
rect 580 5300 1940 5310
rect 2570 5300 2590 5310
rect 3060 5300 3540 5310
rect 5190 5300 5200 5310
rect 6290 5300 6350 5310
rect 6690 5300 6730 5310
rect 7690 5300 7840 5310
rect 8490 5300 8530 5310
rect 8730 5300 8770 5310
rect 8780 5300 9120 5310
rect 9160 5300 9250 5310
rect 9370 5300 9420 5310
rect 9460 5300 9520 5310
rect 9620 5300 9990 5310
rect 590 5290 1940 5300
rect 2580 5290 2590 5300
rect 2840 5290 2860 5300
rect 2990 5290 3540 5300
rect 5190 5290 5200 5300
rect 6320 5290 6330 5300
rect 6720 5290 6740 5300
rect 7640 5290 7680 5300
rect 7690 5290 7840 5300
rect 8500 5290 8530 5300
rect 8680 5290 9110 5300
rect 9160 5290 9250 5300
rect 9380 5290 9430 5300
rect 9470 5290 9510 5300
rect 9620 5290 9940 5300
rect 9980 5290 9990 5300
rect 610 5280 1940 5290
rect 2970 5280 3530 5290
rect 5100 5280 5110 5290
rect 5180 5280 5200 5290
rect 7570 5280 7580 5290
rect 7620 5280 7650 5290
rect 7660 5280 7830 5290
rect 8510 5280 8530 5290
rect 8610 5280 8650 5290
rect 8660 5280 9030 5290
rect 9080 5280 9100 5290
rect 9170 5280 9260 5290
rect 9390 5280 9430 5290
rect 9470 5280 9510 5290
rect 9560 5280 9580 5290
rect 9620 5280 9940 5290
rect 9980 5280 9990 5290
rect 630 5270 1400 5280
rect 1410 5270 1950 5280
rect 2970 5270 3530 5280
rect 5180 5270 5190 5280
rect 5200 5270 5210 5280
rect 7570 5270 7600 5280
rect 7610 5270 7670 5280
rect 7680 5270 7840 5280
rect 8520 5270 8550 5280
rect 8610 5270 9020 5280
rect 9090 5270 9100 5280
rect 9170 5270 9270 5280
rect 9400 5270 9430 5280
rect 9470 5270 9510 5280
rect 9550 5270 9850 5280
rect 9880 5270 9940 5280
rect 9980 5270 9990 5280
rect 610 5260 730 5270
rect 740 5260 1390 5270
rect 1400 5260 1950 5270
rect 2610 5260 2630 5270
rect 2910 5260 2920 5270
rect 2960 5260 3490 5270
rect 3500 5260 3520 5270
rect 7470 5260 7480 5270
rect 7500 5260 7510 5270
rect 7550 5260 7600 5270
rect 7610 5260 7620 5270
rect 7630 5260 7650 5270
rect 7660 5260 7850 5270
rect 8520 5260 8940 5270
rect 8970 5260 9030 5270
rect 9180 5260 9350 5270
rect 9400 5260 9430 5270
rect 9480 5260 9520 5270
rect 9550 5260 9850 5270
rect 9890 5260 9940 5270
rect 9990 5260 9990 5270
rect 620 5250 1380 5260
rect 1390 5250 1950 5260
rect 2620 5250 2640 5260
rect 2910 5250 3500 5260
rect 3510 5250 3520 5260
rect 5080 5250 5090 5260
rect 7450 5250 7460 5260
rect 7480 5250 7490 5260
rect 7500 5250 7580 5260
rect 7600 5250 7610 5260
rect 7630 5250 7650 5260
rect 7680 5250 7850 5260
rect 7860 5250 7870 5260
rect 8520 5250 8920 5260
rect 8980 5250 9030 5260
rect 9180 5250 9350 5260
rect 9400 5250 9440 5260
rect 9480 5250 9760 5260
rect 9790 5250 9850 5260
rect 9900 5250 9950 5260
rect 9990 5250 9990 5260
rect 630 5240 1370 5250
rect 1380 5240 1950 5250
rect 2630 5240 2650 5250
rect 2920 5240 3500 5250
rect 7440 5240 7580 5250
rect 7600 5240 7610 5250
rect 7630 5240 7640 5250
rect 7680 5240 7850 5250
rect 7860 5240 7870 5250
rect 8510 5240 8840 5250
rect 8850 5240 8890 5250
rect 8900 5240 8910 5250
rect 8980 5240 9030 5250
rect 9180 5240 9300 5250
rect 9310 5240 9350 5250
rect 9400 5240 9440 5250
rect 9470 5240 9740 5250
rect 9810 5240 9850 5250
rect 9920 5240 9950 5250
rect 9990 5240 9990 5250
rect 630 5230 1360 5240
rect 1370 5230 1950 5240
rect 2930 5230 3500 5240
rect 7450 5230 7540 5240
rect 7550 5230 7580 5240
rect 7590 5230 7640 5240
rect 7660 5230 7670 5240
rect 7680 5230 7860 5240
rect 8430 5230 8830 5240
rect 8890 5230 8900 5240
rect 8990 5230 9040 5240
rect 9180 5230 9290 5240
rect 9390 5230 9720 5240
rect 9820 5230 9850 5240
rect 9930 5230 9960 5240
rect 9990 5230 9990 5240
rect 620 5220 1950 5230
rect 2950 5220 3500 5230
rect 7440 5220 7450 5230
rect 7460 5220 7520 5230
rect 7550 5220 7560 5230
rect 7600 5220 7620 5230
rect 7640 5220 7650 5230
rect 7660 5220 7670 5230
rect 7680 5220 7850 5230
rect 8420 5220 8830 5230
rect 9000 5220 9040 5230
rect 9180 5220 9290 5230
rect 9390 5220 9720 5230
rect 9830 5220 9850 5230
rect 9950 5220 9960 5230
rect 620 5210 650 5220
rect 670 5210 1960 5220
rect 2720 5210 2730 5220
rect 2960 5210 3500 5220
rect 7440 5210 7530 5220
rect 7600 5210 7610 5220
rect 7640 5210 7650 5220
rect 7670 5210 7860 5220
rect 8380 5210 8750 5220
rect 8780 5210 8820 5220
rect 8880 5210 8900 5220
rect 9000 5210 9040 5220
rect 9190 5210 9290 5220
rect 9380 5210 9710 5220
rect 9760 5210 9790 5220
rect 9840 5210 9860 5220
rect 9950 5210 9970 5220
rect 620 5200 650 5210
rect 690 5200 1960 5210
rect 2680 5200 2730 5210
rect 3000 5200 3490 5210
rect 5120 5200 5130 5210
rect 7440 5200 7530 5210
rect 7540 5200 7550 5210
rect 7620 5200 7630 5210
rect 7640 5200 7650 5210
rect 7660 5200 7860 5210
rect 8360 5200 8750 5210
rect 8790 5200 8810 5210
rect 8890 5200 8910 5210
rect 9010 5200 9050 5210
rect 9190 5200 9310 5210
rect 9360 5200 9710 5210
rect 9750 5200 9790 5210
rect 9840 5200 9860 5210
rect 9900 5200 9910 5210
rect 620 5190 640 5200
rect 700 5190 1830 5200
rect 1840 5190 1960 5200
rect 2690 5190 2730 5200
rect 3010 5190 3350 5200
rect 3360 5190 3480 5200
rect 5120 5190 5130 5200
rect 7440 5190 7540 5200
rect 7550 5190 7560 5200
rect 7590 5190 7610 5200
rect 7670 5190 7860 5200
rect 8330 5190 8680 5200
rect 8730 5190 8740 5200
rect 8810 5190 8820 5200
rect 8880 5190 8900 5200
rect 9010 5190 9040 5200
rect 9100 5190 9110 5200
rect 9190 5190 9550 5200
rect 9600 5190 9710 5200
rect 9750 5190 9790 5200
rect 9840 5190 9870 5200
rect 9900 5190 9930 5200
rect 630 5180 640 5190
rect 710 5180 1810 5190
rect 1850 5180 1960 5190
rect 2700 5180 2740 5190
rect 3020 5180 3480 5190
rect 5080 5180 5090 5190
rect 7440 5180 7540 5190
rect 7600 5180 7610 5190
rect 7630 5180 7870 5190
rect 8270 5180 8650 5190
rect 8880 5180 8900 5190
rect 8910 5180 8920 5190
rect 9020 5180 9050 5190
rect 9110 5180 9130 5190
rect 9190 5180 9520 5190
rect 9610 5180 9710 5190
rect 9750 5180 9800 5190
rect 9840 5180 9870 5190
rect 9910 5180 9940 5190
rect 630 5170 640 5180
rect 700 5170 1800 5180
rect 1860 5170 1960 5180
rect 2720 5170 2760 5180
rect 3010 5170 3330 5180
rect 3340 5170 3470 5180
rect 5080 5170 5110 5180
rect 7440 5170 7540 5180
rect 7590 5170 7680 5180
rect 7690 5170 7870 5180
rect 8260 5170 8620 5180
rect 8800 5170 8820 5180
rect 8890 5170 8910 5180
rect 9030 5170 9060 5180
rect 9110 5170 9150 5180
rect 9190 5170 9510 5180
rect 9620 5170 9710 5180
rect 9760 5170 9800 5180
rect 9840 5170 9870 5180
rect 9910 5170 9960 5180
rect 630 5160 640 5170
rect 710 5160 1800 5170
rect 1860 5160 1960 5170
rect 2730 5160 2790 5170
rect 3010 5160 3470 5170
rect 5090 5160 5100 5170
rect 5130 5160 5140 5170
rect 7450 5160 7550 5170
rect 7560 5160 7890 5170
rect 8230 5160 8610 5170
rect 8720 5160 8740 5170
rect 8890 5160 8910 5170
rect 9030 5160 9060 5170
rect 9110 5160 9440 5170
rect 9470 5160 9500 5170
rect 9620 5160 9710 5170
rect 9760 5160 9810 5170
rect 9850 5160 9880 5170
rect 9920 5160 9970 5170
rect 620 5150 640 5160
rect 720 5150 1790 5160
rect 1830 5150 1850 5160
rect 1860 5150 1960 5160
rect 2740 5150 2800 5160
rect 3010 5150 3460 5160
rect 5130 5150 5140 5160
rect 7450 5150 7890 5160
rect 8230 5150 8600 5160
rect 8700 5150 8740 5160
rect 8890 5150 8910 5160
rect 9040 5150 9070 5160
rect 9110 5150 9400 5160
rect 9480 5150 9500 5160
rect 9550 5150 9580 5160
rect 9630 5150 9720 5160
rect 9760 5150 9810 5160
rect 9850 5150 9880 5160
rect 9920 5150 9980 5160
rect 620 5140 640 5150
rect 740 5140 1800 5150
rect 1840 5140 1960 5150
rect 2750 5140 2810 5150
rect 3040 5140 3450 5150
rect 5120 5140 5140 5150
rect 7450 5140 7570 5150
rect 7610 5140 7620 5150
rect 7640 5140 7880 5150
rect 8170 5140 8180 5150
rect 8210 5140 8600 5150
rect 8700 5140 8740 5150
rect 8890 5140 8900 5150
rect 9050 5140 9080 5150
rect 9100 5140 9370 5150
rect 9480 5140 9500 5150
rect 9550 5140 9580 5150
rect 9630 5140 9720 5150
rect 9760 5140 9810 5150
rect 9850 5140 9880 5150
rect 9920 5140 9990 5150
rect 620 5130 650 5140
rect 740 5130 1800 5140
rect 1840 5130 1970 5140
rect 2760 5130 2830 5140
rect 3040 5130 3450 5140
rect 5120 5130 5140 5140
rect 7450 5130 7560 5140
rect 7590 5130 7610 5140
rect 7640 5130 7880 5140
rect 8200 5130 8470 5140
rect 8520 5130 8650 5140
rect 8700 5130 8750 5140
rect 8830 5130 8850 5140
rect 8900 5130 8910 5140
rect 9050 5130 9370 5140
rect 9470 5130 9500 5140
rect 9550 5130 9590 5140
rect 9630 5130 9720 5140
rect 9770 5130 9810 5140
rect 9850 5130 9890 5140
rect 9930 5130 9990 5140
rect 620 5120 660 5130
rect 740 5120 1800 5130
rect 1880 5120 1890 5130
rect 1900 5120 1970 5130
rect 2780 5120 2860 5130
rect 3000 5120 3010 5130
rect 3030 5120 3310 5130
rect 3320 5120 3440 5130
rect 7450 5120 7520 5130
rect 7530 5120 7580 5130
rect 7590 5120 7600 5130
rect 7620 5120 7630 5130
rect 7640 5120 7870 5130
rect 8080 5120 8090 5130
rect 8130 5120 8140 5130
rect 8220 5120 8430 5130
rect 8520 5120 8650 5130
rect 8700 5120 8760 5130
rect 8810 5120 8850 5130
rect 8900 5120 8910 5130
rect 8970 5120 9010 5130
rect 9040 5120 9280 5130
rect 9340 5120 9360 5130
rect 9430 5120 9510 5130
rect 9550 5120 9590 5130
rect 9630 5120 9720 5130
rect 9770 5120 9810 5130
rect 9850 5120 9890 5130
rect 9920 5120 9990 5130
rect 630 5110 670 5120
rect 740 5110 1780 5120
rect 1860 5110 1890 5120
rect 1900 5110 1970 5120
rect 2800 5110 2900 5120
rect 2990 5110 3000 5120
rect 3030 5110 3430 5120
rect 7450 5110 7870 5120
rect 8030 5110 8110 5120
rect 8220 5110 8420 5120
rect 8520 5110 8650 5120
rect 8700 5110 8770 5120
rect 8810 5110 8850 5120
rect 8910 5110 8920 5120
rect 8960 5110 9250 5120
rect 9340 5110 9360 5120
rect 9410 5110 9510 5120
rect 9550 5110 9600 5120
rect 9640 5110 9730 5120
rect 9850 5110 9990 5120
rect 630 5100 670 5110
rect 750 5100 1800 5110
rect 1860 5100 1970 5110
rect 2820 5100 2930 5110
rect 2990 5100 3000 5110
rect 3030 5100 3430 5110
rect 5180 5100 5190 5110
rect 7450 5100 7460 5110
rect 7470 5100 7540 5110
rect 7550 5100 7560 5110
rect 7570 5100 7880 5110
rect 8030 5100 8110 5110
rect 8210 5100 8410 5110
rect 8500 5100 8660 5110
rect 8700 5100 8770 5110
rect 8810 5100 8860 5110
rect 8900 5100 8930 5110
rect 8960 5100 9230 5110
rect 9340 5100 9370 5110
rect 9410 5100 9520 5110
rect 9560 5100 9600 5110
rect 9640 5100 9730 5110
rect 9840 5100 9990 5110
rect 630 5090 680 5100
rect 750 5090 1800 5100
rect 1860 5090 1880 5100
rect 1890 5090 1980 5100
rect 2850 5090 2960 5100
rect 2980 5090 3010 5100
rect 3030 5090 3420 5100
rect 5180 5090 5190 5100
rect 7450 5090 7880 5100
rect 8040 5090 8130 5100
rect 8170 5090 8180 5100
rect 8210 5090 8220 5100
rect 8230 5090 8320 5100
rect 8380 5090 8400 5100
rect 8470 5090 8660 5100
rect 8710 5090 8770 5100
rect 8820 5090 8860 5100
rect 8900 5090 9220 5100
rect 9320 5090 9370 5100
rect 9480 5090 9520 5100
rect 9560 5090 9600 5100
rect 9640 5090 9740 5100
rect 9830 5090 9990 5100
rect 640 5080 690 5090
rect 750 5080 1790 5090
rect 1810 5080 1820 5090
rect 1880 5080 1980 5090
rect 2870 5080 3410 5090
rect 5180 5080 5200 5090
rect 7450 5080 7880 5090
rect 8040 5080 8110 5090
rect 8120 5080 8130 5090
rect 8140 5080 8150 5090
rect 8170 5080 8190 5090
rect 8220 5080 8290 5090
rect 8470 5080 8670 5090
rect 8710 5080 8760 5090
rect 8820 5080 8880 5090
rect 8890 5080 9130 5090
rect 9200 5080 9230 5090
rect 9310 5080 9370 5090
rect 9480 5080 9520 5090
rect 9560 5080 9610 5090
rect 9640 5080 9770 5090
rect 9800 5080 9990 5090
rect 650 5070 700 5080
rect 740 5070 1770 5080
rect 1870 5070 1970 5080
rect 2870 5070 2880 5080
rect 2890 5070 3410 5080
rect 7450 5070 7880 5080
rect 8040 5070 8120 5080
rect 8140 5070 8160 5080
rect 8210 5070 8270 5080
rect 8520 5070 8660 5080
rect 8710 5070 8770 5080
rect 8820 5070 9110 5080
rect 9210 5070 9270 5080
rect 9310 5070 9370 5080
rect 9470 5070 9530 5080
rect 9560 5070 9600 5080
rect 9640 5070 9990 5080
rect 650 5060 1760 5070
rect 1880 5060 1980 5070
rect 2980 5060 3400 5070
rect 7450 5060 7890 5070
rect 8050 5060 8130 5070
rect 8170 5060 8180 5070
rect 8240 5060 8250 5070
rect 8530 5060 8670 5070
rect 8720 5060 8780 5070
rect 8810 5060 9090 5070
rect 9200 5060 9270 5070
rect 9320 5060 9380 5070
rect 9450 5060 9530 5070
rect 9570 5060 9580 5070
rect 9640 5060 9990 5070
rect 650 5050 1770 5060
rect 1880 5050 1990 5060
rect 3040 5050 3300 5060
rect 3330 5050 3390 5060
rect 7450 5050 7900 5060
rect 8050 5050 8110 5060
rect 8120 5050 8130 5060
rect 8330 5050 8340 5060
rect 8520 5050 8670 5060
rect 8720 5050 9040 5060
rect 9060 5050 9090 5060
rect 9180 5050 9270 5060
rect 9320 5050 9390 5060
rect 9420 5050 9530 5060
rect 9630 5050 9990 5060
rect 480 5040 500 5050
rect 620 5040 1780 5050
rect 1880 5040 1990 5050
rect 3050 5040 3080 5050
rect 3090 5040 3310 5050
rect 3330 5040 3380 5050
rect 7390 5040 7420 5050
rect 7430 5040 7900 5050
rect 8050 5040 8110 5050
rect 8330 5040 8340 5050
rect 8350 5040 8360 5050
rect 8410 5040 8420 5050
rect 8500 5040 8680 5050
rect 8720 5040 9030 5050
rect 9070 5040 9090 5050
rect 9180 5040 9270 5050
rect 9320 5040 9390 5050
rect 9430 5040 9530 5050
rect 9620 5040 9990 5050
rect 470 5030 1760 5040
rect 1780 5030 1790 5040
rect 1890 5030 1990 5040
rect 3050 5030 3330 5040
rect 3340 5030 3370 5040
rect 7440 5030 7900 5040
rect 8090 5030 8100 5040
rect 8330 5030 8350 5040
rect 8480 5030 8690 5040
rect 8710 5030 8970 5040
rect 9000 5030 9020 5040
rect 9070 5030 9130 5040
rect 9180 5030 9280 5040
rect 9320 5030 9390 5040
rect 9430 5030 9470 5040
rect 9500 5030 9540 5040
rect 9600 5030 9990 5040
rect 470 5020 1750 5030
rect 1790 5020 1800 5030
rect 1880 5020 1990 5030
rect 3050 5020 3360 5030
rect 3370 5020 3390 5030
rect 7350 5020 7390 5030
rect 7460 5020 7900 5030
rect 8400 5020 8430 5030
rect 8480 5020 8960 5030
rect 9010 5020 9030 5030
rect 9080 5020 9130 5030
rect 9180 5020 9280 5030
rect 9330 5020 9390 5030
rect 9510 5020 9990 5030
rect 460 5010 1750 5020
rect 1800 5010 1810 5020
rect 1870 5010 2000 5020
rect 3040 5010 3350 5020
rect 3370 5010 3390 5020
rect 7350 5010 7430 5020
rect 7480 5010 7880 5020
rect 8400 5010 8430 5020
rect 8550 5010 8880 5020
rect 8920 5010 8960 5020
rect 9010 5010 9030 5020
rect 9080 5010 9130 5020
rect 9190 5010 9280 5020
rect 9330 5010 9390 5020
rect 9510 5010 9990 5020
rect 430 5000 440 5010
rect 460 5000 1760 5010
rect 1820 5000 2020 5010
rect 3030 5000 3340 5010
rect 4170 5000 4180 5010
rect 7340 5000 7370 5010
rect 7380 5000 7470 5010
rect 7500 5000 7890 5010
rect 7910 5000 7930 5010
rect 8380 5000 8430 5010
rect 8550 5000 8860 5010
rect 8940 5000 8950 5010
rect 9010 5000 9030 5010
rect 9080 5000 9140 5010
rect 9190 5000 9290 5010
rect 9330 5000 9400 5010
rect 9490 5000 9990 5010
rect 430 4990 450 5000
rect 460 4990 1770 5000
rect 1820 4990 1830 5000
rect 1840 4990 2020 5000
rect 2030 4990 2040 5000
rect 2050 4990 2060 5000
rect 3000 4990 3330 5000
rect 3350 4990 3360 5000
rect 7350 4990 7500 5000
rect 7530 4990 7890 5000
rect 8400 4990 8440 5000
rect 8550 4990 8870 5000
rect 9080 4990 9150 5000
rect 9190 4990 9300 5000
rect 9330 4990 9400 5000
rect 9450 4990 9990 5000
rect 440 4980 450 4990
rect 480 4980 1780 4990
rect 1830 4980 2060 4990
rect 2990 4980 3260 4990
rect 3270 4980 3330 4990
rect 3350 4980 3360 4990
rect 7350 4980 7860 4990
rect 7870 4980 7890 4990
rect 8410 4980 8440 4990
rect 8530 4980 8760 4990
rect 8840 4980 8870 4990
rect 9020 4980 9030 4990
rect 9080 4980 9140 4990
rect 9190 4980 9300 4990
rect 9330 4980 9690 4990
rect 9700 4980 9990 4990
rect 440 4970 450 4980
rect 500 4970 1800 4980
rect 1830 4970 2060 4980
rect 2970 4970 3340 4980
rect 4330 4970 4350 4980
rect 4540 4970 4550 4980
rect 7350 4970 7840 4980
rect 8420 4970 8460 4980
rect 8490 4970 8740 4980
rect 8850 4970 8870 4980
rect 9020 4970 9030 4980
rect 9090 4970 9150 4980
rect 9200 4970 9300 4980
rect 9330 4970 9650 4980
rect 9720 4970 9990 4980
rect 440 4960 450 4970
rect 550 4960 1820 4970
rect 1830 4960 2100 4970
rect 2950 4960 3340 4970
rect 4010 4960 4060 4970
rect 4210 4960 4310 4970
rect 4350 4960 4370 4970
rect 7350 4960 7840 4970
rect 8350 4960 8360 4970
rect 8410 4960 8670 4970
rect 8710 4960 8740 4970
rect 8860 4960 8870 4970
rect 9020 4960 9040 4970
rect 9090 4960 9150 4970
rect 9200 4960 9310 4970
rect 9330 4960 9620 4970
rect 9710 4960 9990 4970
rect 440 4950 450 4960
rect 560 4950 1850 4960
rect 1890 4950 2120 4960
rect 2910 4950 2920 4960
rect 2940 4950 3230 4960
rect 3250 4950 3340 4960
rect 4010 4950 4040 4960
rect 4050 4950 4060 4960
rect 4200 4950 4330 4960
rect 7340 4950 7840 4960
rect 8350 4950 8380 4960
rect 8410 4950 8640 4960
rect 8720 4950 8730 4960
rect 8860 4950 8880 4960
rect 9020 4950 9050 4960
rect 9090 4950 9150 4960
rect 9210 4950 9610 4960
rect 9710 4950 9990 4960
rect 430 4940 440 4950
rect 590 4940 1040 4950
rect 1050 4940 1860 4950
rect 1890 4940 2130 4950
rect 2900 4940 2920 4950
rect 2930 4940 3220 4950
rect 3240 4940 3330 4950
rect 4010 4940 4080 4950
rect 4200 4940 4410 4950
rect 7340 4940 7830 4950
rect 8350 4940 8620 4950
rect 8710 4940 8730 4950
rect 8780 4940 8800 4950
rect 8860 4940 8880 4950
rect 9030 4940 9050 4950
rect 9090 4940 9140 4950
rect 9260 4940 9540 4950
rect 9580 4940 9610 4950
rect 9680 4940 9990 4950
rect 610 4930 1040 4940
rect 1060 4930 1860 4940
rect 1890 4930 2150 4940
rect 2890 4930 3220 4940
rect 3230 4930 3330 4940
rect 4010 4930 4060 4940
rect 4190 4930 4350 4940
rect 4380 4930 4430 4940
rect 7340 4930 7760 4940
rect 8280 4930 8310 4940
rect 8340 4930 8600 4940
rect 8710 4930 8740 4940
rect 8800 4930 8810 4940
rect 8860 4930 8890 4940
rect 9030 4930 9060 4940
rect 9100 4930 9130 4940
rect 9280 4930 9540 4940
rect 9580 4930 9610 4940
rect 9660 4930 9990 4940
rect 640 4920 1040 4930
rect 1060 4920 2160 4930
rect 2280 4920 2290 4930
rect 2880 4920 3210 4930
rect 3220 4920 3300 4930
rect 3310 4920 3330 4930
rect 4010 4920 4040 4930
rect 4200 4920 4350 4930
rect 4410 4920 4450 4930
rect 5690 4920 5700 4930
rect 5840 4920 5900 4930
rect 7340 4920 7760 4930
rect 8270 4920 8600 4930
rect 8690 4920 8740 4930
rect 8860 4920 8900 4930
rect 9030 4920 9060 4930
rect 9100 4920 9120 4930
rect 9290 4920 9460 4930
rect 9480 4920 9540 4930
rect 9580 4920 9610 4930
rect 9660 4920 9990 4930
rect 670 4910 680 4920
rect 690 4910 1040 4920
rect 1070 4910 2160 4920
rect 2280 4910 2290 4920
rect 2880 4910 3210 4920
rect 3220 4910 3300 4920
rect 3310 4910 3320 4920
rect 4020 4910 4050 4920
rect 4120 4910 4140 4920
rect 4210 4910 4390 4920
rect 4410 4910 4430 4920
rect 4440 4910 4470 4920
rect 5840 4910 5920 4920
rect 6230 4910 6290 4920
rect 7340 4910 7690 4920
rect 7730 4910 7750 4920
rect 8260 4910 8500 4920
rect 8560 4910 8590 4920
rect 8650 4910 8740 4920
rect 8850 4910 8900 4920
rect 8990 4910 9000 4920
rect 9030 4910 9060 4920
rect 9100 4910 9110 4920
rect 9300 4910 9450 4920
rect 9490 4910 9530 4920
rect 9590 4910 9620 4920
rect 9660 4910 9670 4920
rect 9720 4910 9990 4920
rect 720 4900 1070 4910
rect 1090 4900 2170 4910
rect 2270 4900 2300 4910
rect 2860 4900 3190 4910
rect 3220 4900 3300 4910
rect 3310 4900 3320 4910
rect 4010 4900 4020 4910
rect 4090 4900 4160 4910
rect 4200 4900 4490 4910
rect 5860 4900 5940 4910
rect 6200 4900 6290 4910
rect 7350 4900 7680 4910
rect 8260 4900 8470 4910
rect 8650 4900 8740 4910
rect 8850 4900 8900 4910
rect 8980 4900 9000 4910
rect 9040 4900 9070 4910
rect 9300 4900 9390 4910
rect 9410 4900 9450 4910
rect 9500 4900 9530 4910
rect 9590 4900 9620 4910
rect 9720 4900 9990 4910
rect 740 4890 1070 4900
rect 1080 4890 2180 4900
rect 2260 4890 2310 4900
rect 2830 4890 3170 4900
rect 3210 4890 3290 4900
rect 3310 4890 3320 4900
rect 3980 4890 4010 4900
rect 4070 4890 4160 4900
rect 4200 4890 4470 4900
rect 4700 4890 4740 4900
rect 5880 4890 5950 4900
rect 6180 4890 6300 4900
rect 7360 4890 7670 4900
rect 8150 4890 8200 4900
rect 8210 4890 8470 4900
rect 8580 4890 8590 4900
rect 8710 4890 8750 4900
rect 8840 4890 8910 4900
rect 8950 4890 9000 4900
rect 9030 4890 9100 4900
rect 9310 4890 9380 4900
rect 9420 4890 9450 4900
rect 9510 4890 9530 4900
rect 9590 4890 9620 4900
rect 9720 4890 9990 4900
rect 740 4880 1040 4890
rect 1050 4880 1060 4890
rect 1080 4880 2190 4890
rect 2260 4880 2280 4890
rect 2810 4880 3160 4890
rect 3200 4880 3310 4890
rect 3890 4880 3900 4890
rect 3980 4880 4000 4890
rect 4050 4880 4170 4890
rect 4200 4880 4510 4890
rect 4620 4880 4640 4890
rect 4650 4880 4670 4890
rect 4680 4880 4740 4890
rect 5890 4880 5960 4890
rect 6160 4880 6300 4890
rect 7370 4880 7670 4890
rect 8080 4880 8100 4890
rect 8140 4880 8460 4890
rect 8710 4880 8750 4890
rect 8850 4880 8910 4890
rect 8950 4880 9090 4890
rect 9360 4880 9380 4890
rect 9420 4880 9450 4890
rect 9510 4880 9530 4890
rect 9590 4880 9620 4890
rect 9700 4880 9990 4890
rect 760 4870 1060 4880
rect 1090 4870 2200 4880
rect 2210 4870 2220 4880
rect 2260 4870 2270 4880
rect 2300 4870 2340 4880
rect 2800 4870 3150 4880
rect 3190 4870 3320 4880
rect 3890 4870 3910 4880
rect 3970 4870 3990 4880
rect 4030 4870 4180 4880
rect 4200 4870 4570 4880
rect 4610 4870 4780 4880
rect 6140 4870 6300 4880
rect 6410 4870 6440 4880
rect 7350 4870 7670 4880
rect 8090 4870 8100 4880
rect 8110 4870 8460 4880
rect 8590 4870 8600 4880
rect 8710 4870 8750 4880
rect 8800 4870 8810 4880
rect 8870 4870 8910 4880
rect 8950 4870 9080 4880
rect 9360 4870 9380 4880
rect 9430 4870 9450 4880
rect 9600 4870 9620 4880
rect 9670 4870 9990 4880
rect 760 4860 1010 4870
rect 1020 4860 1060 4870
rect 1100 4860 2240 4870
rect 2250 4860 2260 4870
rect 2280 4860 2330 4870
rect 2790 4860 3100 4870
rect 3120 4860 3140 4870
rect 3190 4860 3320 4870
rect 3710 4860 3720 4870
rect 3870 4860 3920 4870
rect 3930 4860 3970 4870
rect 4010 4860 4190 4870
rect 4200 4860 4850 4870
rect 6120 4860 6220 4870
rect 6230 4860 6300 4870
rect 6420 4860 6440 4870
rect 7390 4860 7470 4870
rect 7480 4860 7680 4870
rect 8090 4860 8320 4870
rect 8360 4860 8460 4870
rect 8590 4860 8600 4870
rect 8690 4860 8760 4870
rect 8800 4860 8820 4870
rect 8880 4860 8920 4870
rect 8940 4860 9080 4870
rect 9350 4860 9390 4870
rect 9430 4860 9460 4870
rect 9600 4860 9630 4870
rect 9670 4860 9990 4870
rect 750 4850 1070 4860
rect 1120 4850 2330 4860
rect 2780 4850 3100 4860
rect 3180 4850 3320 4860
rect 3690 4850 3720 4860
rect 3830 4850 3840 4860
rect 3870 4850 3960 4860
rect 4000 4850 4890 4860
rect 6120 4850 6160 4860
rect 6230 4850 6280 4860
rect 6420 4850 6430 4860
rect 7410 4850 7680 4860
rect 8080 4850 8250 4860
rect 8280 4850 8290 4860
rect 8370 4850 8470 4860
rect 8590 4850 8620 4860
rect 8660 4850 8760 4860
rect 8800 4850 8830 4860
rect 8880 4850 9060 4860
rect 9340 4850 9390 4860
rect 9430 4850 9460 4860
rect 9600 4850 9630 4860
rect 9680 4850 9720 4860
rect 9750 4850 9990 4860
rect 790 4840 1030 4850
rect 1100 4840 1110 4850
rect 1120 4840 2330 4850
rect 2780 4840 3090 4850
rect 3130 4840 3150 4850
rect 3170 4840 3240 4850
rect 3270 4840 3320 4850
rect 3680 4840 3710 4850
rect 3820 4840 3850 4850
rect 3870 4840 3950 4850
rect 3990 4840 4260 4850
rect 4270 4840 4910 4850
rect 6120 4840 6140 4850
rect 6220 4840 6270 4850
rect 7350 4840 7680 4850
rect 8090 4840 8250 4850
rect 8380 4840 8470 4850
rect 8580 4840 8620 4850
rect 8660 4840 8760 4850
rect 8800 4840 8850 4850
rect 8870 4840 9060 4850
rect 9330 4840 9390 4850
rect 9430 4840 9460 4850
rect 9610 4840 9630 4850
rect 9760 4840 9990 4850
rect 350 4830 390 4840
rect 790 4830 1030 4840
rect 1070 4830 1100 4840
rect 1110 4830 2340 4840
rect 2790 4830 3080 4840
rect 3130 4830 3140 4840
rect 3170 4830 3230 4840
rect 3270 4830 3320 4840
rect 3660 4830 3670 4840
rect 3680 4830 3700 4840
rect 3820 4830 3850 4840
rect 3860 4830 3940 4840
rect 3980 4830 4910 4840
rect 4960 4830 4970 4840
rect 5600 4830 5620 4840
rect 6230 4830 6250 4840
rect 7350 4830 7680 4840
rect 8090 4830 8200 4840
rect 8230 4830 8240 4840
rect 8370 4830 8470 4840
rect 8570 4830 8620 4840
rect 8660 4830 8680 4840
rect 8740 4830 8770 4840
rect 8800 4830 9060 4840
rect 9330 4830 9390 4840
rect 9440 4830 9470 4840
rect 9610 4830 9640 4840
rect 9760 4830 9990 4840
rect 330 4820 470 4830
rect 490 4820 510 4830
rect 730 4820 1020 4830
rect 1090 4820 1140 4830
rect 1150 4820 2350 4830
rect 2790 4820 3070 4830
rect 3120 4820 3140 4830
rect 3160 4820 3230 4830
rect 3270 4820 3330 4830
rect 3350 4820 3360 4830
rect 3660 4820 3700 4830
rect 3810 4820 3930 4830
rect 3970 4820 4910 4830
rect 4940 4820 4950 4830
rect 4970 4820 4990 4830
rect 5600 4820 5620 4830
rect 7350 4820 7360 4830
rect 7370 4820 7570 4830
rect 7590 4820 7690 4830
rect 8080 4820 8190 4830
rect 8320 4820 8480 4830
rect 8560 4820 8620 4830
rect 8740 4820 9060 4830
rect 9330 4820 9400 4830
rect 9440 4820 9470 4830
rect 9510 4820 9520 4830
rect 9550 4820 9570 4830
rect 9610 4820 9640 4830
rect 9740 4820 9990 4830
rect 310 4810 540 4820
rect 680 4810 840 4820
rect 870 4810 980 4820
rect 990 4810 1030 4820
rect 1100 4810 2350 4820
rect 2810 4810 3050 4820
rect 3150 4810 3210 4820
rect 3270 4810 3320 4820
rect 3650 4810 3690 4820
rect 3710 4810 3720 4820
rect 3770 4810 3780 4820
rect 3810 4810 3910 4820
rect 3950 4810 4910 4820
rect 4930 4810 4960 4820
rect 4980 4810 5000 4820
rect 5590 4810 5620 4820
rect 7370 4810 7450 4820
rect 7460 4810 7690 4820
rect 7910 4810 7930 4820
rect 7940 4810 7950 4820
rect 7970 4810 7980 4820
rect 8090 4810 8120 4820
rect 8150 4810 8190 4820
rect 8320 4810 8480 4820
rect 8540 4810 8620 4820
rect 8740 4810 9040 4820
rect 9340 4810 9400 4820
rect 9440 4810 9470 4820
rect 9520 4810 9570 4820
rect 9610 4810 9640 4820
rect 9710 4810 9990 4820
rect 290 4800 330 4810
rect 460 4800 550 4810
rect 580 4800 600 4810
rect 630 4800 740 4810
rect 880 4800 1030 4810
rect 1040 4800 1050 4810
rect 1100 4800 1140 4810
rect 1150 4800 2350 4810
rect 2840 4800 3040 4810
rect 3150 4800 3220 4810
rect 3280 4800 3310 4810
rect 3640 4800 3680 4810
rect 3690 4800 3780 4810
rect 3790 4800 3900 4810
rect 3930 4800 4910 4810
rect 5000 4800 5010 4810
rect 5560 4800 5620 4810
rect 7370 4800 7520 4810
rect 7540 4800 7690 4810
rect 7830 4800 7930 4810
rect 7940 4800 7980 4810
rect 8360 4800 8480 4810
rect 8530 4800 8630 4810
rect 8720 4800 9000 4810
rect 9030 4800 9040 4810
rect 9340 4800 9400 4810
rect 9440 4800 9480 4810
rect 9520 4800 9570 4810
rect 9610 4800 9990 4810
rect 250 4790 300 4800
rect 480 4790 550 4800
rect 580 4790 600 4800
rect 880 4790 890 4800
rect 900 4790 1030 4800
rect 1100 4790 2360 4800
rect 2920 4790 3040 4800
rect 3140 4790 3240 4800
rect 3260 4790 3270 4800
rect 3280 4790 3320 4800
rect 3630 4790 3880 4800
rect 3910 4790 4930 4800
rect 4950 4790 4990 4800
rect 5000 4790 5030 4800
rect 5230 4790 5240 4800
rect 5560 4790 5610 4800
rect 7370 4790 7510 4800
rect 7520 4790 7690 4800
rect 7780 4790 7790 4800
rect 7820 4790 7920 4800
rect 7940 4790 7980 4800
rect 8380 4790 8490 4800
rect 8530 4790 8630 4800
rect 8680 4790 8990 4800
rect 9340 4790 9410 4800
rect 9450 4790 9480 4800
rect 9520 4790 9580 4800
rect 9610 4790 9990 4800
rect 320 4780 460 4790
rect 520 4780 600 4790
rect 880 4780 900 4790
rect 920 4780 1040 4790
rect 1100 4780 2360 4790
rect 2370 4780 2390 4790
rect 2930 4780 3030 4790
rect 3130 4780 3320 4790
rect 3610 4780 3870 4790
rect 3900 4780 5030 4790
rect 5220 4780 5240 4790
rect 5550 4780 5610 4790
rect 7370 4780 7500 4790
rect 7510 4780 7700 4790
rect 7750 4780 7990 4790
rect 8390 4780 8490 4790
rect 8530 4780 8920 4790
rect 8940 4780 9000 4790
rect 9340 4780 9410 4790
rect 9450 4780 9480 4790
rect 9520 4780 9990 4790
rect 310 4770 480 4780
rect 550 4770 590 4780
rect 850 4770 880 4780
rect 900 4770 1050 4780
rect 1060 4770 1070 4780
rect 1110 4770 2390 4780
rect 2930 4770 3020 4780
rect 3130 4770 3240 4780
rect 3290 4770 3330 4780
rect 3600 4770 3620 4780
rect 3630 4770 3800 4780
rect 3810 4770 3860 4780
rect 3890 4770 5040 4780
rect 5530 4770 5600 4780
rect 7360 4770 7480 4780
rect 7500 4770 7710 4780
rect 7740 4770 7960 4780
rect 8400 4770 8490 4780
rect 8540 4770 8910 4780
rect 8950 4770 9000 4780
rect 9350 4770 9410 4780
rect 9450 4770 9490 4780
rect 9520 4770 9990 4780
rect 320 4760 500 4770
rect 960 4760 990 4770
rect 1010 4760 1080 4770
rect 1130 4760 2380 4770
rect 2940 4760 3000 4770
rect 3120 4760 3250 4770
rect 3300 4760 3330 4770
rect 3600 4760 3610 4770
rect 3620 4760 3790 4770
rect 3810 4760 3840 4770
rect 3870 4760 5060 4770
rect 5530 4760 5580 4770
rect 7360 4760 7470 4770
rect 7480 4760 7930 4770
rect 7950 4760 7960 4770
rect 8260 4760 8300 4770
rect 8400 4760 8500 4770
rect 8530 4760 8820 4770
rect 8860 4760 8910 4770
rect 8960 4760 9000 4770
rect 9350 4760 9410 4770
rect 9450 4760 9990 4770
rect 350 4750 530 4760
rect 950 4750 990 4760
rect 1010 4750 1070 4760
rect 1140 4750 2380 4760
rect 2410 4750 2420 4760
rect 3120 4750 3250 4760
rect 3290 4750 3340 4760
rect 3590 4750 3780 4760
rect 3800 4750 3830 4760
rect 3880 4750 5070 4760
rect 5510 4750 5580 4760
rect 7400 4750 7450 4760
rect 7470 4750 7890 4760
rect 8260 4750 8300 4760
rect 8310 4750 8350 4760
rect 8400 4750 8510 4760
rect 8520 4750 8800 4760
rect 8880 4750 8910 4760
rect 8970 4750 9000 4760
rect 9350 4750 9420 4760
rect 9450 4750 9920 4760
rect 9960 4750 9990 4760
rect 370 4740 550 4750
rect 960 4740 980 4750
rect 1000 4740 1010 4750
rect 1020 4740 1090 4750
rect 1110 4740 1140 4750
rect 1170 4740 2400 4750
rect 2410 4740 2420 4750
rect 3110 4740 3260 4750
rect 3300 4740 3340 4750
rect 3580 4740 3780 4750
rect 3800 4740 3820 4750
rect 3850 4740 3910 4750
rect 3930 4740 3980 4750
rect 3990 4740 5080 4750
rect 5510 4740 5570 4750
rect 7380 4740 7440 4750
rect 7460 4740 7870 4750
rect 8330 4740 8340 4750
rect 8400 4740 8790 4750
rect 8890 4740 8910 4750
rect 8990 4740 9000 4750
rect 9300 4740 9310 4750
rect 9350 4740 9870 4750
rect 410 4730 570 4740
rect 650 4730 670 4740
rect 1000 4730 1010 4740
rect 1030 4730 1090 4740
rect 1120 4730 1140 4740
rect 1150 4730 2410 4740
rect 2420 4730 2430 4740
rect 3100 4730 3260 4740
rect 3300 4730 3340 4740
rect 3580 4730 3790 4740
rect 3800 4730 3820 4740
rect 3830 4730 5080 4740
rect 5090 4730 5110 4740
rect 5510 4730 5550 4740
rect 7370 4730 7440 4740
rect 7450 4730 7860 4740
rect 8390 4730 8780 4740
rect 8890 4730 8920 4740
rect 9300 4730 9320 4740
rect 9350 4730 9850 4740
rect 430 4720 620 4730
rect 640 4720 690 4730
rect 1020 4720 1030 4730
rect 1040 4720 1060 4730
rect 1070 4720 1090 4730
rect 1160 4720 2430 4730
rect 3090 4720 3270 4730
rect 3300 4720 3350 4730
rect 3560 4720 3580 4730
rect 3600 4720 3780 4730
rect 3800 4720 5090 4730
rect 5110 4720 5120 4730
rect 5500 4720 5550 4730
rect 7370 4720 7430 4730
rect 7440 4720 7770 4730
rect 7800 4720 7850 4730
rect 8380 4720 8780 4730
rect 8830 4720 8850 4730
rect 8900 4720 8920 4730
rect 9290 4720 9330 4730
rect 9350 4720 9840 4730
rect 450 4710 630 4720
rect 650 4710 710 4720
rect 1040 4710 1100 4720
rect 1170 4710 2430 4720
rect 3090 4710 3270 4720
rect 3310 4710 3350 4720
rect 3560 4710 3580 4720
rect 3600 4710 3770 4720
rect 3800 4710 5100 4720
rect 5500 4710 5550 4720
rect 7370 4710 7410 4720
rect 7440 4710 7730 4720
rect 7820 4710 7830 4720
rect 8130 4710 8140 4720
rect 8370 4710 8640 4720
rect 8670 4710 8780 4720
rect 8820 4710 8850 4720
rect 8900 4710 8920 4720
rect 9290 4710 9840 4720
rect 470 4700 660 4710
rect 670 4700 730 4710
rect 990 4700 1000 4710
rect 1030 4700 1080 4710
rect 1090 4700 1100 4710
rect 1170 4700 2440 4710
rect 2450 4700 2470 4710
rect 3100 4700 3170 4710
rect 3180 4700 3270 4710
rect 3320 4700 3350 4710
rect 3550 4700 3770 4710
rect 3790 4700 5100 4710
rect 5130 4700 5140 4710
rect 5500 4700 5570 4710
rect 7370 4700 7400 4710
rect 7430 4700 7720 4710
rect 8270 4700 8300 4710
rect 8350 4700 8600 4710
rect 8680 4700 8780 4710
rect 8820 4700 8860 4710
rect 8900 4700 8930 4710
rect 9290 4700 9830 4710
rect 500 4690 670 4700
rect 680 4690 740 4700
rect 1030 4690 1060 4700
rect 1090 4690 1110 4700
rect 1170 4690 2440 4700
rect 2460 4690 2480 4700
rect 3080 4690 3090 4700
rect 3110 4690 3170 4700
rect 3190 4690 3270 4700
rect 3310 4690 3350 4700
rect 3490 4690 3500 4700
rect 3550 4690 3620 4700
rect 3640 4690 5110 4700
rect 5130 4690 5150 4700
rect 5500 4690 5580 4700
rect 7390 4690 7400 4700
rect 7420 4690 7660 4700
rect 7690 4690 7700 4700
rect 8270 4690 8570 4700
rect 8670 4690 8780 4700
rect 8820 4690 8860 4700
rect 8900 4690 8930 4700
rect 9280 4690 9820 4700
rect 510 4680 750 4690
rect 1040 4680 1120 4690
rect 1170 4680 2450 4690
rect 2470 4680 2480 4690
rect 2530 4680 2540 4690
rect 3060 4680 3100 4690
rect 3110 4680 3130 4690
rect 3190 4680 3270 4690
rect 3290 4680 3350 4690
rect 3540 4680 3600 4690
rect 3610 4680 3630 4690
rect 3640 4680 5120 4690
rect 5140 4680 5160 4690
rect 5510 4680 5580 4690
rect 6530 4680 6550 4690
rect 7410 4680 7630 4690
rect 8210 4680 8240 4690
rect 8260 4680 8560 4690
rect 8660 4680 8780 4690
rect 8830 4680 8860 4690
rect 8910 4680 8930 4690
rect 9280 4680 9810 4690
rect 520 4670 760 4680
rect 1010 4670 1030 4680
rect 1050 4670 1160 4680
rect 1180 4670 2510 4680
rect 2520 4670 2540 4680
rect 3060 4670 3100 4680
rect 3190 4670 3260 4680
rect 3290 4670 3340 4680
rect 3500 4670 3600 4680
rect 3610 4670 3700 4680
rect 3720 4670 5120 4680
rect 5150 4670 5170 4680
rect 5520 4670 5590 4680
rect 6540 4670 6550 4680
rect 7400 4670 7610 4680
rect 8130 4670 8140 4680
rect 8190 4670 8500 4680
rect 8540 4670 8560 4680
rect 8640 4670 8790 4680
rect 8830 4670 8870 4680
rect 8910 4670 8930 4680
rect 9270 4670 9800 4680
rect 540 4660 800 4670
rect 1040 4660 1170 4670
rect 1180 4660 2500 4670
rect 2510 4660 2550 4670
rect 2730 4660 2760 4670
rect 3060 4660 3100 4670
rect 3180 4660 3250 4670
rect 3280 4660 3340 4670
rect 3500 4660 3610 4670
rect 3620 4660 3780 4670
rect 3790 4660 5130 4670
rect 5160 4660 5180 4670
rect 5520 4660 5590 4670
rect 6520 4660 6560 4670
rect 7390 4660 7600 4670
rect 8120 4660 8150 4670
rect 8180 4660 8500 4670
rect 8540 4660 8590 4670
rect 8650 4660 8790 4670
rect 8830 4660 8870 4670
rect 8910 4660 8930 4670
rect 8980 4660 8990 4670
rect 9270 4660 9790 4670
rect 560 4650 830 4660
rect 1070 4650 1140 4660
rect 1180 4650 2480 4660
rect 2490 4650 2500 4660
rect 2510 4650 2540 4660
rect 2720 4650 2780 4660
rect 3060 4650 3090 4660
rect 3120 4650 3130 4660
rect 3180 4650 3340 4660
rect 3500 4650 5140 4660
rect 5160 4650 5190 4660
rect 5520 4650 5730 4660
rect 6520 4650 6560 4660
rect 7390 4650 7510 4660
rect 7560 4650 7600 4660
rect 7670 4650 7700 4660
rect 7830 4650 7910 4660
rect 8120 4650 8500 4660
rect 8550 4650 8610 4660
rect 8650 4650 8790 4660
rect 8830 4650 8870 4660
rect 8910 4650 8940 4660
rect 9260 4650 9780 4660
rect 580 4640 840 4650
rect 1090 4640 1100 4650
rect 1110 4640 2490 4650
rect 2500 4640 2540 4650
rect 2550 4640 2560 4650
rect 2720 4640 2770 4650
rect 3070 4640 3090 4650
rect 3180 4640 3320 4650
rect 3490 4640 5140 4650
rect 5170 4640 5190 4650
rect 5530 4640 5760 4650
rect 6510 4640 6560 4650
rect 7390 4640 7490 4650
rect 7580 4640 7590 4650
rect 7650 4640 7710 4650
rect 7830 4640 7920 4650
rect 8110 4640 8500 4650
rect 8550 4640 8610 4650
rect 8650 4640 8790 4650
rect 8840 4640 8870 4650
rect 8910 4640 8940 4650
rect 9260 4640 9770 4650
rect 600 4630 840 4640
rect 1120 4630 1180 4640
rect 1190 4630 2490 4640
rect 2500 4630 2590 4640
rect 2720 4630 2780 4640
rect 2800 4630 2810 4640
rect 2820 4630 2830 4640
rect 3000 4630 3010 4640
rect 3030 4630 3040 4640
rect 3050 4630 3080 4640
rect 3110 4630 3130 4640
rect 3160 4630 3170 4640
rect 3180 4630 3320 4640
rect 3480 4630 5150 4640
rect 5180 4630 5200 4640
rect 5540 4630 5750 4640
rect 5760 4630 5790 4640
rect 6500 4630 6560 4640
rect 7390 4630 7480 4640
rect 7590 4630 7600 4640
rect 7700 4630 7720 4640
rect 7820 4630 7870 4640
rect 7990 4630 8010 4640
rect 8120 4630 8300 4640
rect 8370 4630 8490 4640
rect 8560 4630 8610 4640
rect 8650 4630 8800 4640
rect 8910 4630 8950 4640
rect 9260 4630 9760 4640
rect 620 4620 850 4630
rect 1120 4620 1130 4630
rect 1200 4620 2600 4630
rect 2710 4620 2720 4630
rect 2800 4620 2880 4630
rect 3000 4620 3010 4630
rect 3030 4620 3120 4630
rect 3130 4620 3140 4630
rect 3160 4620 3300 4630
rect 3480 4620 5160 4630
rect 5180 4620 5200 4630
rect 5540 4620 5610 4630
rect 5630 4620 5750 4630
rect 5770 4620 5800 4630
rect 6490 4620 6560 4630
rect 7400 4620 7470 4630
rect 7700 4620 7720 4630
rect 7820 4620 7870 4630
rect 7990 4620 8080 4630
rect 8120 4620 8280 4630
rect 8380 4620 8490 4630
rect 8570 4620 8620 4630
rect 8660 4620 8800 4630
rect 8910 4620 8980 4630
rect 9250 4620 9750 4630
rect 630 4610 860 4620
rect 1220 4610 2730 4620
rect 2750 4610 2840 4620
rect 2960 4610 2970 4620
rect 3020 4610 3130 4620
rect 3170 4610 3230 4620
rect 3240 4610 3290 4620
rect 3480 4610 5170 4620
rect 5180 4610 5210 4620
rect 5540 4610 5600 4620
rect 5640 4610 5750 4620
rect 5770 4610 5780 4620
rect 6110 4610 6160 4620
rect 6360 4610 6380 4620
rect 6480 4610 6530 4620
rect 7400 4610 7470 4620
rect 7700 4610 7730 4620
rect 7840 4610 7860 4620
rect 7980 4610 8070 4620
rect 8120 4610 8230 4620
rect 8240 4610 8270 4620
rect 8390 4610 8490 4620
rect 8570 4610 8620 4620
rect 8660 4610 8810 4620
rect 8900 4610 8970 4620
rect 9250 4610 9740 4620
rect 650 4600 870 4610
rect 1220 4600 2850 4610
rect 2930 4600 2990 4610
rect 3020 4600 3030 4610
rect 3040 4600 3050 4610
rect 3060 4600 3130 4610
rect 3160 4600 3220 4610
rect 3240 4600 3280 4610
rect 3470 4600 5180 4610
rect 5190 4600 5210 4610
rect 5540 4600 5570 4610
rect 5650 4600 5750 4610
rect 6080 4600 6180 4610
rect 6190 4600 6510 4610
rect 7410 4600 7470 4610
rect 7520 4600 7540 4610
rect 7600 4600 7610 4610
rect 7690 4600 7730 4610
rect 7850 4600 7870 4610
rect 7960 4600 7970 4610
rect 7980 4600 8070 4610
rect 8130 4600 8190 4610
rect 8390 4600 8490 4610
rect 8580 4600 8620 4610
rect 8660 4600 8830 4610
rect 8880 4600 8970 4610
rect 9250 4600 9730 4610
rect 660 4590 870 4600
rect 1210 4590 2820 4600
rect 2830 4590 2850 4600
rect 2870 4590 3030 4600
rect 3050 4590 3130 4600
rect 3170 4590 3200 4600
rect 3240 4590 3270 4600
rect 3470 4590 5180 4600
rect 5190 4590 5220 4600
rect 5540 4590 5570 4600
rect 5650 4590 5750 4600
rect 6200 4590 6510 4600
rect 7420 4590 7470 4600
rect 7590 4590 7610 4600
rect 7670 4590 7730 4600
rect 7850 4590 7910 4600
rect 7930 4590 8080 4600
rect 8130 4590 8160 4600
rect 8390 4590 8490 4600
rect 8580 4590 8620 4600
rect 8660 4590 8960 4600
rect 9240 4590 9720 4600
rect 670 4580 890 4590
rect 1210 4580 2810 4590
rect 2830 4580 3110 4590
rect 3120 4580 3140 4590
rect 3230 4580 3270 4590
rect 3470 4580 5220 4590
rect 5550 4580 5570 4590
rect 5660 4580 5760 4590
rect 6260 4580 6500 4590
rect 7390 4580 7480 4590
rect 7590 4580 7610 4590
rect 7660 4580 7720 4590
rect 7850 4580 8070 4590
rect 8130 4580 8150 4590
rect 8400 4580 8490 4590
rect 8590 4580 8620 4590
rect 8670 4580 8960 4590
rect 9240 4580 9710 4590
rect 700 4570 910 4580
rect 1220 4570 3020 4580
rect 3040 4570 3130 4580
rect 3230 4570 3260 4580
rect 3460 4570 5230 4580
rect 5550 4570 5570 4580
rect 5660 4570 5760 4580
rect 6290 4570 6310 4580
rect 6320 4570 6480 4580
rect 7390 4570 7470 4580
rect 7580 4570 7610 4580
rect 7660 4570 7690 4580
rect 7720 4570 7730 4580
rect 7830 4570 8070 4580
rect 8240 4570 8260 4580
rect 8400 4570 8490 4580
rect 8600 4570 8630 4580
rect 8670 4570 8960 4580
rect 9240 4570 9700 4580
rect 700 4560 920 4570
rect 1230 4560 3030 4570
rect 3040 4560 3130 4570
rect 3230 4560 3250 4570
rect 3450 4560 5230 4570
rect 5550 4560 5570 4570
rect 5680 4560 5780 4570
rect 6330 4560 6480 4570
rect 7390 4560 7480 4570
rect 7570 4560 7610 4570
rect 7740 4560 7750 4570
rect 7810 4560 8080 4570
rect 8200 4560 8270 4570
rect 8400 4560 8490 4570
rect 8600 4560 8630 4570
rect 8670 4560 8950 4570
rect 9240 4560 9690 4570
rect 710 4550 930 4560
rect 1200 4550 1210 4560
rect 1240 4550 2800 4560
rect 2820 4550 2980 4560
rect 2990 4550 3030 4560
rect 3080 4550 3130 4560
rect 3160 4550 3170 4560
rect 3230 4550 3250 4560
rect 3440 4550 5240 4560
rect 5550 4550 5560 4560
rect 5680 4550 5790 4560
rect 6330 4550 6470 4560
rect 7390 4550 7490 4560
rect 7550 4550 7610 4560
rect 7740 4550 8010 4560
rect 8050 4550 8060 4560
rect 8200 4550 8260 4560
rect 8390 4550 8480 4560
rect 8610 4550 8640 4560
rect 8660 4550 8950 4560
rect 9240 4550 9690 4560
rect 720 4540 940 4550
rect 1170 4540 2810 4550
rect 2820 4540 2980 4550
rect 2990 4540 3040 4550
rect 3060 4540 3150 4550
rect 3160 4540 3180 4550
rect 3230 4540 3240 4550
rect 3440 4540 5250 4550
rect 5690 4540 5790 4550
rect 6320 4540 6450 4550
rect 7390 4540 7490 4550
rect 7540 4540 7610 4550
rect 7720 4540 8000 4550
rect 8380 4540 8480 4550
rect 8550 4540 8570 4550
rect 8600 4540 8950 4550
rect 9230 4540 9680 4550
rect 730 4530 950 4540
rect 1160 4530 2970 4540
rect 2990 4530 3030 4540
rect 3060 4530 3070 4540
rect 3080 4530 3190 4540
rect 3430 4530 5240 4540
rect 5690 4530 5800 4540
rect 6310 4530 6460 4540
rect 7400 4530 7490 4540
rect 7540 4530 7620 4540
rect 7690 4530 7910 4540
rect 8380 4530 8480 4540
rect 8530 4530 8580 4540
rect 8590 4530 8940 4540
rect 9230 4530 9670 4540
rect 770 4520 980 4530
rect 1160 4520 2980 4530
rect 2990 4520 3010 4530
rect 3020 4520 3040 4530
rect 3060 4520 3070 4530
rect 3090 4520 3200 4530
rect 3430 4520 5250 4530
rect 5700 4520 5810 4530
rect 6300 4520 6470 4530
rect 7400 4520 7480 4530
rect 7540 4520 7640 4530
rect 7650 4520 7890 4530
rect 8250 4520 8280 4530
rect 8400 4520 8490 4530
rect 8520 4520 8940 4530
rect 9230 4520 9660 4530
rect 680 4510 690 4520
rect 770 4510 980 4520
rect 1170 4510 1180 4520
rect 1200 4510 2980 4520
rect 3030 4510 3040 4520
rect 3060 4510 3070 4520
rect 3090 4510 3210 4520
rect 3420 4510 3870 4520
rect 3920 4510 5260 4520
rect 5700 4510 5770 4520
rect 5850 4510 5860 4520
rect 6290 4510 6420 4520
rect 7410 4510 7500 4520
rect 7540 4510 7830 4520
rect 7850 4510 7880 4520
rect 8250 4510 8280 4520
rect 8400 4510 8500 4520
rect 8510 4510 8940 4520
rect 9230 4510 9650 4520
rect 780 4500 990 4510
rect 1170 4500 1190 4510
rect 1200 4500 2990 4510
rect 3030 4500 3240 4510
rect 3420 4500 3870 4510
rect 3940 4500 5260 4510
rect 5720 4500 5770 4510
rect 5840 4500 5860 4510
rect 6290 4500 6410 4510
rect 7350 4500 7360 4510
rect 7410 4500 7500 4510
rect 7540 4500 7780 4510
rect 8220 4500 8280 4510
rect 8410 4500 8930 4510
rect 9230 4500 9640 4510
rect 9990 4500 9990 4510
rect 600 4490 610 4500
rect 650 4490 670 4500
rect 690 4490 730 4500
rect 770 4490 1000 4500
rect 1160 4490 1180 4500
rect 1190 4490 3000 4500
rect 3030 4490 3060 4500
rect 3090 4490 3250 4500
rect 3410 4490 3860 4500
rect 3950 4490 5270 4500
rect 5720 4490 5760 4500
rect 6280 4490 6410 4500
rect 7420 4490 7510 4500
rect 7530 4490 7760 4500
rect 8220 4490 8290 4500
rect 8410 4490 8930 4500
rect 9220 4490 9630 4500
rect 9980 4490 9990 4500
rect 590 4480 610 4490
rect 640 4480 1010 4490
rect 1140 4480 1150 4490
rect 1160 4480 1170 4490
rect 1180 4480 2880 4490
rect 2890 4480 2990 4490
rect 3040 4480 3050 4490
rect 3110 4480 3260 4490
rect 3400 4480 3860 4490
rect 3950 4480 5280 4490
rect 5740 4480 5760 4490
rect 6240 4480 6400 4490
rect 7430 4480 7750 4490
rect 8370 4480 8920 4490
rect 9220 4480 9620 4490
rect 9970 4480 9990 4490
rect 580 4470 600 4480
rect 620 4470 1010 4480
rect 1100 4470 1120 4480
rect 1170 4470 2990 4480
rect 3040 4470 3050 4480
rect 3110 4470 3270 4480
rect 3400 4470 3860 4480
rect 3950 4470 5280 4480
rect 5740 4470 5790 4480
rect 6190 4470 6200 4480
rect 6240 4470 6390 4480
rect 7420 4470 7750 4480
rect 7850 4470 7860 4480
rect 8340 4470 8920 4480
rect 9220 4470 9610 4480
rect 9960 4470 9990 4480
rect 470 4460 520 4470
rect 580 4460 590 4470
rect 620 4460 1030 4470
rect 1130 4460 1140 4470
rect 1170 4460 2990 4470
rect 3040 4460 3050 4470
rect 3130 4460 3140 4470
rect 3150 4460 3160 4470
rect 3180 4460 3270 4470
rect 3400 4460 3870 4470
rect 3950 4460 5280 4470
rect 5750 4460 5780 4470
rect 6190 4460 6210 4470
rect 6220 4460 6380 4470
rect 7420 4460 7760 4470
rect 7840 4460 7870 4470
rect 8290 4460 8910 4470
rect 9220 4460 9600 4470
rect 9950 4460 9990 4470
rect 440 4450 460 4460
rect 470 4450 520 4460
rect 570 4450 600 4460
rect 610 4450 690 4460
rect 700 4450 1040 4460
rect 1160 4450 2850 4460
rect 2860 4450 2980 4460
rect 3040 4450 3050 4460
rect 3200 4450 3230 4460
rect 3250 4450 3270 4460
rect 3390 4450 5290 4460
rect 5760 4450 5780 4460
rect 6200 4450 6360 4460
rect 7420 4450 7790 4460
rect 7840 4450 7870 4460
rect 8270 4450 8910 4460
rect 9210 4450 9590 4460
rect 9950 4450 9990 4460
rect 460 4440 540 4450
rect 600 4440 680 4450
rect 690 4440 1060 4450
rect 1160 4440 2840 4450
rect 2860 4440 2990 4450
rect 3040 4440 3060 4450
rect 3070 4440 3090 4450
rect 3190 4440 3220 4450
rect 3230 4440 3240 4450
rect 3390 4440 3900 4450
rect 3910 4440 4620 4450
rect 4630 4440 5290 4450
rect 6210 4440 6220 4450
rect 6250 4440 6340 4450
rect 7420 4440 7780 4450
rect 7850 4440 7880 4450
rect 8240 4440 8880 4450
rect 9210 4440 9580 4450
rect 9940 4440 9990 4450
rect 450 4430 500 4440
rect 510 4430 560 4440
rect 580 4430 1070 4440
rect 1110 4430 1140 4440
rect 1170 4430 2820 4440
rect 2860 4430 2980 4440
rect 3050 4430 3070 4440
rect 3190 4430 3230 4440
rect 3390 4430 3860 4440
rect 3950 4430 4610 4440
rect 4650 4430 5300 4440
rect 6250 4430 6340 4440
rect 7420 4430 7780 4440
rect 7850 4430 7870 4440
rect 8020 4430 8030 4440
rect 8180 4430 8850 4440
rect 9210 4430 9570 4440
rect 9930 4430 9990 4440
rect 290 4420 310 4430
rect 410 4420 460 4430
rect 490 4420 1080 4430
rect 1110 4420 1140 4430
rect 1150 4420 2630 4430
rect 2640 4420 2750 4430
rect 2760 4420 2970 4430
rect 3050 4420 3070 4430
rect 3200 4420 3230 4430
rect 3380 4420 3850 4430
rect 3950 4420 4230 4430
rect 4280 4420 4610 4430
rect 4670 4420 4780 4430
rect 4790 4420 5300 4430
rect 6250 4420 6320 4430
rect 7420 4420 7790 4430
rect 7850 4420 7880 4430
rect 8020 4420 8030 4430
rect 8100 4420 8110 4430
rect 8170 4420 8850 4430
rect 9210 4420 9560 4430
rect 9920 4420 9990 4430
rect 280 4410 320 4420
rect 350 4410 360 4420
rect 400 4410 410 4420
rect 420 4410 460 4420
rect 480 4410 1090 4420
rect 1100 4410 2740 4420
rect 2760 4410 2840 4420
rect 2850 4410 2960 4420
rect 3060 4410 3070 4420
rect 3210 4410 3220 4420
rect 3300 4410 3310 4420
rect 3380 4410 3830 4420
rect 3950 4410 4230 4420
rect 4300 4410 4600 4420
rect 4690 4410 4780 4420
rect 4790 4410 5310 4420
rect 6250 4410 6300 4420
rect 7430 4410 7790 4420
rect 7860 4410 7880 4420
rect 8020 4410 8030 4420
rect 8040 4410 8050 4420
rect 8090 4410 8120 4420
rect 8170 4410 8850 4420
rect 9200 4410 9550 4420
rect 9910 4410 9990 4420
rect 280 4400 330 4410
rect 360 4400 2650 4410
rect 2670 4400 2840 4410
rect 2860 4400 2870 4410
rect 2880 4400 2960 4410
rect 3300 4400 3310 4410
rect 3370 4400 3820 4410
rect 3910 4400 3920 4410
rect 3940 4400 4240 4410
rect 4310 4400 4600 4410
rect 4710 4400 5310 4410
rect 6250 4400 6290 4410
rect 7430 4400 7790 4410
rect 7860 4400 7890 4410
rect 8010 4400 8130 4410
rect 8170 4400 8850 4410
rect 9200 4400 9540 4410
rect 9900 4400 9990 4410
rect 220 4390 230 4400
rect 260 4390 350 4400
rect 370 4390 380 4400
rect 400 4390 2640 4400
rect 2670 4390 2800 4400
rect 2820 4390 2830 4400
rect 2850 4390 2940 4400
rect 2950 4390 2960 4400
rect 3210 4390 3220 4400
rect 3300 4390 3320 4400
rect 3370 4390 3820 4400
rect 3920 4390 4250 4400
rect 4310 4390 4590 4400
rect 4730 4390 4820 4400
rect 4860 4390 4880 4400
rect 4890 4390 5310 4400
rect 6240 4390 6280 4400
rect 7430 4390 7790 4400
rect 7860 4390 7890 4400
rect 8000 4390 8120 4400
rect 8170 4390 8680 4400
rect 8710 4390 8850 4400
rect 9200 4390 9530 4400
rect 9890 4390 9990 4400
rect 220 4380 370 4390
rect 380 4380 2640 4390
rect 2650 4380 2700 4390
rect 2710 4380 2800 4390
rect 2840 4380 2860 4390
rect 2880 4380 2930 4390
rect 2940 4380 2960 4390
rect 3220 4380 3230 4390
rect 3300 4380 3320 4390
rect 3360 4380 3820 4390
rect 3920 4380 4260 4390
rect 4320 4380 4590 4390
rect 4740 4380 4800 4390
rect 4900 4380 5320 4390
rect 6210 4380 6270 4390
rect 7430 4380 7790 4390
rect 7860 4380 7890 4390
rect 7900 4380 7910 4390
rect 7990 4380 8130 4390
rect 8170 4380 8660 4390
rect 8730 4380 8850 4390
rect 9200 4380 9510 4390
rect 9880 4380 9990 4390
rect 220 4370 2630 4380
rect 2650 4370 2700 4380
rect 2720 4370 2820 4380
rect 2830 4370 2840 4380
rect 2880 4370 2950 4380
rect 3130 4370 3170 4380
rect 3300 4370 3330 4380
rect 3360 4370 3830 4380
rect 3930 4370 4270 4380
rect 4320 4370 4580 4380
rect 4780 4370 4790 4380
rect 4900 4370 5330 4380
rect 6190 4370 6220 4380
rect 7430 4370 7800 4380
rect 7860 4370 8130 4380
rect 8170 4370 8600 4380
rect 8620 4370 8650 4380
rect 8730 4370 8850 4380
rect 9190 4370 9500 4380
rect 9870 4370 9990 4380
rect 220 4360 2590 4370
rect 2600 4360 2620 4370
rect 2630 4360 2700 4370
rect 2710 4360 2820 4370
rect 2840 4360 2930 4370
rect 3090 4360 3170 4370
rect 3210 4360 3220 4370
rect 3310 4360 3330 4370
rect 3360 4360 3840 4370
rect 3920 4360 4280 4370
rect 4330 4360 4570 4370
rect 4900 4360 5330 4370
rect 7430 4360 7800 4370
rect 7860 4360 8140 4370
rect 8170 4360 8540 4370
rect 8560 4360 8590 4370
rect 8620 4360 8650 4370
rect 8680 4360 8850 4370
rect 9190 4360 9490 4370
rect 9860 4360 9990 4370
rect 240 4350 2820 4360
rect 2840 4350 2940 4360
rect 3080 4350 3180 4360
rect 3200 4350 3230 4360
rect 3310 4350 3330 4360
rect 3360 4350 3850 4360
rect 3900 4350 4280 4360
rect 4320 4350 4570 4360
rect 4920 4350 5330 4360
rect 7430 4350 7820 4360
rect 7860 4350 8140 4360
rect 8170 4350 8540 4360
rect 8570 4350 8590 4360
rect 8620 4350 8650 4360
rect 8680 4350 8860 4360
rect 9190 4350 9480 4360
rect 9860 4350 9970 4360
rect 240 4340 2580 4350
rect 2590 4340 2740 4350
rect 2750 4340 2820 4350
rect 2840 4340 2920 4350
rect 3060 4340 3160 4350
rect 3210 4340 3240 4350
rect 3310 4340 3330 4350
rect 3340 4340 3850 4350
rect 3860 4340 4170 4350
rect 4190 4340 4200 4350
rect 4230 4340 4300 4350
rect 4320 4340 4560 4350
rect 4930 4340 5340 4350
rect 7430 4340 8140 4350
rect 8180 4340 8490 4350
rect 8510 4340 8540 4350
rect 8620 4340 8650 4350
rect 8730 4340 8860 4350
rect 9190 4340 9470 4350
rect 9850 4340 9900 4350
rect 80 4330 90 4340
rect 240 4330 260 4340
rect 270 4330 2580 4340
rect 2590 4330 2630 4340
rect 2640 4330 2740 4340
rect 2750 4330 2840 4340
rect 2850 4330 2920 4340
rect 3040 4330 3090 4340
rect 3100 4330 3140 4340
rect 3210 4330 3240 4340
rect 3310 4330 4170 4340
rect 4240 4330 4300 4340
rect 4330 4330 4560 4340
rect 4940 4330 5340 4340
rect 7410 4330 8140 4340
rect 8180 4330 8440 4340
rect 8460 4330 8490 4340
rect 8520 4330 8550 4340
rect 8610 4330 8660 4340
rect 8740 4330 8870 4340
rect 9190 4330 9460 4340
rect 9840 4330 9860 4340
rect 70 4320 90 4330
rect 120 4320 130 4330
rect 270 4320 2810 4330
rect 2820 4320 2840 4330
rect 2860 4320 2920 4330
rect 3030 4320 3100 4330
rect 3110 4320 3120 4330
rect 3210 4320 3240 4330
rect 3310 4320 4150 4330
rect 4160 4320 4170 4330
rect 4260 4320 4320 4330
rect 4340 4320 4550 4330
rect 4940 4320 5350 4330
rect 7360 4320 8150 4330
rect 8180 4320 8430 4330
rect 8470 4320 8490 4330
rect 8520 4320 8560 4330
rect 8610 4320 8680 4330
rect 8700 4320 8710 4330
rect 8740 4320 8870 4330
rect 9190 4320 9450 4330
rect 140 4310 150 4320
rect 170 4310 180 4320
rect 210 4310 230 4320
rect 260 4310 2690 4320
rect 2700 4310 2800 4320
rect 2860 4310 2920 4320
rect 3020 4310 3090 4320
rect 3210 4310 3220 4320
rect 3250 4310 3260 4320
rect 3300 4310 4150 4320
rect 4270 4310 4330 4320
rect 4340 4310 4550 4320
rect 4940 4310 5320 4320
rect 5330 4310 5350 4320
rect 7340 4310 8160 4320
rect 8180 4310 8430 4320
rect 8480 4310 8490 4320
rect 8520 4310 8570 4320
rect 8610 4310 8670 4320
rect 8680 4310 8720 4320
rect 8740 4310 8860 4320
rect 9190 4310 9440 4320
rect 80 4300 100 4310
rect 120 4300 2560 4310
rect 2570 4300 2800 4310
rect 2830 4300 2850 4310
rect 2860 4300 2910 4310
rect 3010 4300 3050 4310
rect 3250 4300 3260 4310
rect 3300 4300 4140 4310
rect 4280 4300 4540 4310
rect 4950 4300 5320 4310
rect 5330 4300 5350 4310
rect 7290 4300 8160 4310
rect 8180 4300 8440 4310
rect 8520 4300 8580 4310
rect 8610 4300 8660 4310
rect 8740 4300 8860 4310
rect 9190 4300 9440 4310
rect 70 4290 2560 4300
rect 2590 4290 2830 4300
rect 2850 4290 2910 4300
rect 3000 4290 3040 4300
rect 3080 4290 3100 4300
rect 3200 4290 3210 4300
rect 3250 4290 3260 4300
rect 3270 4290 3280 4300
rect 3300 4290 4140 4300
rect 4290 4290 4530 4300
rect 4960 4290 5350 4300
rect 7250 4290 7350 4300
rect 7370 4290 8160 4300
rect 8180 4290 8440 4300
rect 8530 4290 8580 4300
rect 8610 4290 8660 4300
rect 8740 4290 8860 4300
rect 9190 4290 9430 4300
rect 80 4280 2580 4290
rect 2590 4280 2810 4290
rect 2820 4280 2880 4290
rect 2900 4280 2910 4290
rect 3000 4280 3030 4290
rect 3120 4280 3130 4290
rect 3260 4280 3280 4290
rect 3300 4280 4130 4290
rect 4310 4280 4530 4290
rect 4960 4280 5350 4290
rect 7220 4280 8160 4290
rect 8180 4280 8440 4290
rect 8530 4280 8580 4290
rect 8610 4280 8680 4290
rect 8720 4280 8850 4290
rect 9190 4280 9420 4290
rect 80 4270 2830 4280
rect 2860 4270 2870 4280
rect 2990 4270 3030 4280
rect 3190 4270 3200 4280
rect 3260 4270 3280 4280
rect 3300 4270 4140 4280
rect 4310 4270 4520 4280
rect 4980 4270 5360 4280
rect 7180 4270 7200 4280
rect 7220 4270 8170 4280
rect 8190 4270 8440 4280
rect 8530 4270 8580 4280
rect 8610 4270 8850 4280
rect 9190 4270 9410 4280
rect 80 4260 2810 4270
rect 2860 4260 2890 4270
rect 2980 4260 3020 4270
rect 3190 4260 3200 4270
rect 3290 4260 4140 4270
rect 4330 4260 4510 4270
rect 4970 4260 5360 4270
rect 7240 4260 7400 4270
rect 7440 4260 8170 4270
rect 8190 4260 8440 4270
rect 8530 4260 8590 4270
rect 8610 4260 8850 4270
rect 9190 4260 9400 4270
rect 9790 4260 9800 4270
rect 90 4250 2800 4260
rect 2850 4250 2880 4260
rect 2980 4250 3010 4260
rect 3190 4250 3200 4260
rect 3280 4250 4130 4260
rect 4340 4250 4510 4260
rect 4990 4250 5370 4260
rect 7230 4250 7350 4260
rect 7450 4250 8170 4260
rect 8200 4250 8440 4260
rect 8480 4250 8490 4260
rect 8530 4250 8840 4260
rect 9190 4250 9400 4260
rect 9780 4250 9810 4260
rect 120 4240 2540 4250
rect 2550 4240 2740 4250
rect 2760 4240 2790 4250
rect 2800 4240 2820 4250
rect 2990 4240 3010 4250
rect 3180 4240 3190 4250
rect 3230 4240 3240 4250
rect 3270 4240 4120 4250
rect 4350 4240 4490 4250
rect 5000 4240 5370 4250
rect 7190 4240 7280 4250
rect 7450 4240 8160 4250
rect 8200 4240 8450 4250
rect 8480 4240 8510 4250
rect 8520 4240 8840 4250
rect 9190 4240 9390 4250
rect 9760 4240 9810 4250
rect 0 4230 10 4240
rect 110 4230 2510 4240
rect 2520 4230 2530 4240
rect 2550 4230 2690 4240
rect 2700 4230 2830 4240
rect 2990 4230 3060 4240
rect 3160 4230 3190 4240
rect 3260 4230 4120 4240
rect 4360 4230 4480 4240
rect 5000 4230 5380 4240
rect 7170 4230 7250 4240
rect 7450 4230 8170 4240
rect 8200 4230 8460 4240
rect 8480 4230 8840 4240
rect 9190 4230 9390 4240
rect 9750 4230 9800 4240
rect 0 4220 10 4230
rect 110 4220 2530 4230
rect 2550 4220 2600 4230
rect 2610 4220 2790 4230
rect 2810 4220 2860 4230
rect 2990 4220 3010 4230
rect 3110 4220 3130 4230
rect 3150 4220 3180 4230
rect 3220 4220 3230 4230
rect 3260 4220 4110 4230
rect 4370 4220 4460 4230
rect 5010 4220 5390 4230
rect 7140 4220 7210 4230
rect 7460 4220 8160 4230
rect 8200 4220 8830 4230
rect 9180 4220 9360 4230
rect 9740 4220 9840 4230
rect 0 4210 20 4220
rect 130 4210 2770 4220
rect 2810 4210 2840 4220
rect 2890 4210 2910 4220
rect 2970 4210 3000 4220
rect 3160 4210 3170 4220
rect 3220 4210 3230 4220
rect 3260 4210 4110 4220
rect 4370 4210 4450 4220
rect 5010 4210 5400 4220
rect 7470 4210 8170 4220
rect 8200 4210 8830 4220
rect 9180 4210 9320 4220
rect 9750 4210 9810 4220
rect 0 4200 60 4210
rect 120 4200 2780 4210
rect 2800 4200 2950 4210
rect 2960 4200 3010 4210
rect 3140 4200 3160 4210
rect 3250 4200 4110 4210
rect 4390 4200 4440 4210
rect 5010 4200 5390 4210
rect 7470 4200 8180 4210
rect 8210 4200 8830 4210
rect 9180 4200 9310 4210
rect 9770 4200 9810 4210
rect 9980 4200 9990 4210
rect 10 4190 70 4200
rect 130 4190 150 4200
rect 200 4190 2550 4200
rect 2560 4190 2570 4200
rect 2600 4190 2650 4200
rect 2660 4190 2760 4200
rect 2790 4190 2870 4200
rect 2910 4190 2990 4200
rect 3050 4190 3080 4200
rect 3250 4190 4100 4200
rect 4400 4190 4440 4200
rect 5020 4190 5390 4200
rect 5500 4190 5510 4200
rect 7480 4190 8180 4200
rect 8200 4190 8830 4200
rect 9180 4190 9220 4200
rect 9280 4190 9310 4200
rect 9800 4190 9810 4200
rect 20 4180 30 4190
rect 40 4180 80 4190
rect 130 4180 2570 4190
rect 2610 4180 2640 4190
rect 2660 4180 2760 4190
rect 2790 4180 2820 4190
rect 2930 4180 3000 4190
rect 3240 4180 4100 4190
rect 4410 4180 4440 4190
rect 5030 4180 5390 4190
rect 5500 4180 5540 4190
rect 7240 4180 7290 4190
rect 7480 4180 8180 4190
rect 8210 4180 8820 4190
rect 30 4170 70 4180
rect 130 4170 2570 4180
rect 2600 4170 2630 4180
rect 2660 4170 2670 4180
rect 2690 4170 2700 4180
rect 2710 4170 2760 4180
rect 2790 4170 2810 4180
rect 2950 4170 3000 4180
rect 3230 4170 4090 4180
rect 5030 4170 5380 4180
rect 5500 4170 5540 4180
rect 7270 4170 7310 4180
rect 7480 4170 8180 4180
rect 8210 4170 8820 4180
rect 9830 4170 9860 4180
rect 30 4160 60 4170
rect 130 4160 2580 4170
rect 2610 4160 2650 4170
rect 2660 4160 2680 4170
rect 2780 4160 2810 4170
rect 2970 4160 2990 4170
rect 3170 4160 3180 4170
rect 3210 4160 4090 4170
rect 5040 4160 5400 4170
rect 5500 4160 5560 4170
rect 7270 4160 7310 4170
rect 7480 4160 8190 4170
rect 8200 4160 8820 4170
rect 9280 4160 9310 4170
rect 9840 4160 9870 4170
rect 0 4150 10 4160
rect 40 4150 50 4160
rect 110 4150 2580 4160
rect 2620 4150 2670 4160
rect 2690 4150 2700 4160
rect 2730 4150 2740 4160
rect 2760 4150 2770 4160
rect 2780 4150 2810 4160
rect 3120 4150 3170 4160
rect 3210 4150 3230 4160
rect 3240 4150 3270 4160
rect 3280 4150 4080 4160
rect 5040 4150 5430 4160
rect 5500 4150 5570 4160
rect 7260 4150 7350 4160
rect 7480 4150 8820 4160
rect 9290 4150 9310 4160
rect 9860 4150 9880 4160
rect 0 4140 50 4150
rect 150 4140 2580 4150
rect 2590 4140 2600 4150
rect 2630 4140 2670 4150
rect 2680 4140 2690 4150
rect 2720 4140 2740 4150
rect 2790 4140 2810 4150
rect 3110 4140 3140 4150
rect 3230 4140 3260 4150
rect 3290 4140 4080 4150
rect 5060 4140 5430 4150
rect 5500 4140 5590 4150
rect 7250 4140 7370 4150
rect 7480 4140 8200 4150
rect 8210 4140 8810 4150
rect 9880 4140 9910 4150
rect 0 4130 60 4140
rect 150 4130 2480 4140
rect 2490 4130 2580 4140
rect 2620 4130 2680 4140
rect 2790 4130 2810 4140
rect 3060 4130 3070 4140
rect 3220 4130 3230 4140
rect 3280 4130 4080 4140
rect 4800 4130 4880 4140
rect 5090 4130 5440 4140
rect 5500 4130 5600 4140
rect 7250 4130 7390 4140
rect 7480 4130 8200 4140
rect 8210 4130 8810 4140
rect 9890 4130 9940 4140
rect 0 4120 90 4130
rect 120 4120 130 4130
rect 150 4120 2590 4130
rect 2630 4120 2680 4130
rect 2790 4120 2820 4130
rect 3000 4120 3010 4130
rect 3210 4120 3220 4130
rect 3280 4120 4070 4130
rect 4760 4120 4920 4130
rect 5100 4120 5440 4130
rect 5500 4120 5610 4130
rect 7250 4120 7440 4130
rect 7460 4120 8200 4130
rect 8210 4120 8810 4130
rect 9900 4120 9950 4130
rect 0 4110 90 4120
rect 150 4110 2600 4120
rect 2640 4110 2680 4120
rect 2790 4110 2810 4120
rect 3280 4110 4070 4120
rect 4730 4110 4940 4120
rect 5110 4110 5450 4120
rect 5500 4110 5620 4120
rect 7240 4110 7430 4120
rect 7440 4110 7450 4120
rect 7470 4110 8810 4120
rect 9920 4110 9960 4120
rect 0 4100 100 4110
rect 150 4100 2610 4110
rect 2650 4100 2680 4110
rect 2790 4100 2820 4110
rect 3280 4100 4070 4110
rect 4700 4100 4920 4110
rect 5120 4100 5450 4110
rect 5500 4100 5630 4110
rect 7240 4100 7450 4110
rect 7490 4100 8800 4110
rect 9930 4100 9980 4110
rect 0 4090 110 4100
rect 150 4090 2610 4100
rect 2800 4090 2810 4100
rect 3030 4090 3050 4100
rect 3060 4090 3070 4100
rect 3280 4090 4060 4100
rect 4680 4090 4890 4100
rect 5130 4090 5430 4100
rect 5500 4090 5640 4100
rect 7230 4090 7470 4100
rect 7520 4090 8800 4100
rect 9950 4090 9990 4100
rect 0 4080 110 4090
rect 140 4080 2600 4090
rect 2610 4080 2620 4090
rect 2800 4080 2820 4090
rect 3020 4080 3030 4090
rect 3280 4080 4060 4090
rect 4670 4080 4850 4090
rect 5130 4080 5430 4090
rect 5500 4080 5660 4090
rect 7230 4080 7500 4090
rect 7580 4080 8780 4090
rect 9970 4080 9990 4090
rect 0 4070 130 4080
rect 150 4070 2610 4080
rect 2650 4070 2660 4080
rect 2810 4070 2820 4080
rect 3060 4070 3080 4080
rect 3280 4070 4050 4080
rect 4660 4070 4830 4080
rect 5140 4070 5420 4080
rect 5500 4070 5660 4080
rect 7220 4070 7550 4080
rect 7610 4070 8730 4080
rect 8750 4070 8770 4080
rect 9980 4070 9990 4080
rect 0 4060 140 4070
rect 160 4060 2620 4070
rect 2650 4060 2660 4070
rect 2810 4060 2820 4070
rect 3090 4060 3110 4070
rect 3270 4060 4050 4070
rect 4650 4060 4810 4070
rect 5140 4060 5420 4070
rect 5500 4060 5670 4070
rect 7220 4060 7590 4070
rect 7650 4060 8730 4070
rect 8750 4060 8760 4070
rect 8770 4060 8790 4070
rect 0 4050 2620 4060
rect 2820 4050 2830 4060
rect 3280 4050 4040 4060
rect 4640 4050 4800 4060
rect 5150 4050 5420 4060
rect 5510 4050 5690 4060
rect 7210 4050 7620 4060
rect 7670 4050 8630 4060
rect 8670 4050 8690 4060
rect 8700 4050 8750 4060
rect 8770 4050 8790 4060
rect 0 4040 150 4050
rect 160 4040 2620 4050
rect 3270 4040 4030 4050
rect 4640 4040 4780 4050
rect 5150 4040 5410 4050
rect 5510 4040 5700 4050
rect 7210 4040 7650 4050
rect 7700 4040 8580 4050
rect 8620 4040 8630 4050
rect 8670 4040 8760 4050
rect 0 4030 150 4040
rect 160 4030 2600 4040
rect 2640 4030 2650 4040
rect 3280 4030 4030 4040
rect 4630 4030 4760 4040
rect 5160 4030 5410 4040
rect 5510 4030 5710 4040
rect 7210 4030 7670 4040
rect 7720 4030 8530 4040
rect 8630 4030 8640 4040
rect 8670 4030 8730 4040
rect 8750 4030 8780 4040
rect 0 4020 150 4030
rect 180 4020 2600 4030
rect 3280 4020 4030 4030
rect 4630 4020 4750 4030
rect 5160 4020 5410 4030
rect 5510 4020 5720 4030
rect 7200 4020 7700 4030
rect 7750 4020 8480 4030
rect 8500 4020 8530 4030
rect 8650 4020 8670 4030
rect 8690 4020 8730 4030
rect 8740 4020 8780 4030
rect 0 4010 160 4020
rect 180 4010 2590 4020
rect 3280 4010 4020 4020
rect 4630 4010 4730 4020
rect 5160 4010 5410 4020
rect 5510 4010 5730 4020
rect 7200 4010 7720 4020
rect 7770 4010 8440 4020
rect 8510 4010 8530 4020
rect 8650 4010 8680 4020
rect 8710 4010 8760 4020
rect 0 4000 160 4010
rect 180 4000 2600 4010
rect 3270 4000 4010 4010
rect 4630 4000 4710 4010
rect 5170 4000 5410 4010
rect 5510 4000 5740 4010
rect 7190 4000 7750 4010
rect 7800 4000 8380 4010
rect 8400 4000 8430 4010
rect 8660 4000 8690 4010
rect 8730 4000 8760 4010
rect 0 3990 2610 4000
rect 3270 3990 4000 4000
rect 4630 3990 4680 4000
rect 5170 3990 5410 4000
rect 5510 3990 5760 4000
rect 7190 3990 7780 4000
rect 7820 3990 8340 4000
rect 8410 3990 8430 4000
rect 8500 3990 8510 4000
rect 8540 3990 8560 4000
rect 8680 3990 8700 4000
rect 8740 3990 8760 4000
rect 0 3980 2610 3990
rect 3280 3980 4000 3990
rect 4630 3980 4660 3990
rect 5180 3980 5410 3990
rect 5500 3980 5780 3990
rect 7180 3980 7800 3990
rect 7850 3980 8310 3990
rect 0 3970 2610 3980
rect 3280 3970 3980 3980
rect 4630 3970 4640 3980
rect 5180 3970 5410 3980
rect 5500 3970 5790 3980
rect 7180 3970 7820 3980
rect 7880 3970 8240 3980
rect 8280 3970 8300 3980
rect 8520 3970 8540 3980
rect 0 3960 2610 3970
rect 3280 3960 3960 3970
rect 5200 3960 5410 3970
rect 5500 3960 5820 3970
rect 7170 3960 7850 3970
rect 7900 3960 8200 3970
rect 8530 3960 8560 3970
rect 0 3950 2610 3960
rect 3280 3950 3950 3960
rect 5210 3950 5410 3960
rect 5500 3950 5860 3960
rect 7170 3950 7880 3960
rect 7920 3950 8160 3960
rect 8420 3950 8440 3960
rect 8540 3950 8570 3960
rect 0 3940 2610 3950
rect 3280 3940 3930 3950
rect 5220 3940 5410 3950
rect 5500 3940 5910 3950
rect 5920 3940 5960 3950
rect 7160 3940 7900 3950
rect 7940 3940 8120 3950
rect 8420 3940 8450 3950
rect 8510 3940 8520 3950
rect 8550 3940 8570 3950
rect 9700 3940 9720 3950
rect 0 3930 2610 3940
rect 3280 3930 3910 3940
rect 5220 3930 5420 3940
rect 5490 3930 6010 3940
rect 7160 3930 7920 3940
rect 7960 3930 8100 3940
rect 8430 3930 8450 3940
rect 8520 3930 8530 3940
rect 8640 3930 8660 3940
rect 9690 3930 9730 3940
rect 0 3920 2610 3930
rect 3280 3920 3910 3930
rect 5230 3920 5420 3930
rect 5440 3920 5460 3930
rect 5480 3920 6050 3930
rect 6080 3920 6090 3930
rect 6130 3920 6160 3930
rect 7150 3920 7940 3930
rect 7980 3920 8020 3930
rect 8060 3920 8090 3930
rect 8520 3920 8550 3930
rect 8580 3920 8680 3930
rect 9680 3920 9720 3930
rect 9730 3920 9750 3930
rect 0 3910 2610 3920
rect 3280 3910 3900 3920
rect 5230 3910 5420 3920
rect 5440 3910 6160 3920
rect 7150 3910 7950 3920
rect 8070 3910 8100 3920
rect 8110 3910 8120 3920
rect 8530 3910 8550 3920
rect 8590 3910 8640 3920
rect 8660 3910 8700 3920
rect 9630 3910 9650 3920
rect 9670 3910 9710 3920
rect 9730 3910 9740 3920
rect 9760 3910 9770 3920
rect 0 3900 2590 3910
rect 3280 3900 3900 3910
rect 5230 3900 6000 3910
rect 6010 3900 6140 3910
rect 7140 3900 7970 3910
rect 8070 3900 8190 3910
rect 8300 3900 8320 3910
rect 8550 3900 8590 3910
rect 8600 3900 8650 3910
rect 8670 3900 8700 3910
rect 9620 3900 9650 3910
rect 9660 3900 9740 3910
rect 9760 3900 9780 3910
rect 0 3890 2570 3900
rect 3280 3890 3890 3900
rect 5240 3890 6020 3900
rect 6030 3890 6040 3900
rect 7140 3890 7970 3900
rect 8080 3890 8190 3900
rect 8300 3890 8340 3900
rect 8520 3890 8530 3900
rect 8560 3890 8600 3900
rect 8640 3890 8650 3900
rect 9610 3890 9640 3900
rect 9650 3890 9730 3900
rect 0 3880 2550 3890
rect 3110 3880 3120 3890
rect 3280 3880 3890 3890
rect 5240 3880 6040 3890
rect 7130 3880 7970 3890
rect 8070 3880 8200 3890
rect 8310 3880 8320 3890
rect 8330 3880 8340 3890
rect 8580 3880 8600 3890
rect 9560 3880 9720 3890
rect 0 3870 2530 3880
rect 3100 3870 3110 3880
rect 3280 3870 3880 3880
rect 5250 3870 5990 3880
rect 6000 3870 6020 3880
rect 6040 3870 6060 3880
rect 7130 3870 7970 3880
rect 8010 3870 8020 3880
rect 8050 3870 8210 3880
rect 8540 3870 8550 3880
rect 9490 3870 9520 3880
rect 9550 3870 9720 3880
rect 9820 3870 9830 3880
rect 0 3860 2230 3870
rect 2300 3860 2430 3870
rect 2460 3860 2540 3870
rect 3280 3860 3880 3870
rect 5250 3860 5990 3870
rect 7120 3860 7980 3870
rect 8010 3860 8030 3870
rect 8060 3860 8210 3870
rect 9490 3860 9520 3870
rect 9560 3860 9730 3870
rect 9820 3860 9850 3870
rect 0 3850 2020 3860
rect 2050 3850 2230 3860
rect 2290 3850 2310 3860
rect 2330 3850 2390 3860
rect 2460 3850 2540 3860
rect 3280 3850 3870 3860
rect 4180 3850 4230 3860
rect 5250 3850 5980 3860
rect 7120 3850 7980 3860
rect 8010 3850 8040 3860
rect 8070 3850 8210 3860
rect 9580 3850 9730 3860
rect 9810 3850 9860 3860
rect 0 3840 2020 3850
rect 2040 3840 2240 3850
rect 2300 3840 2320 3850
rect 2340 3840 2400 3850
rect 2470 3840 2570 3850
rect 3280 3840 3860 3850
rect 4150 3840 4250 3850
rect 5260 3840 5970 3850
rect 5980 3840 5990 3850
rect 7110 3840 7990 3850
rect 8020 3840 8060 3850
rect 8080 3840 8210 3850
rect 9590 3840 9720 3850
rect 9800 3840 9860 3850
rect 0 3830 2040 3840
rect 2050 3830 2410 3840
rect 2470 3830 2580 3840
rect 3280 3830 3860 3840
rect 4130 3830 4280 3840
rect 5260 3830 5980 3840
rect 7110 3830 8000 3840
rect 8020 3830 8080 3840
rect 8100 3830 8170 3840
rect 9610 3830 9720 3840
rect 9800 3830 9840 3840
rect 0 3820 2420 3830
rect 2450 3820 2590 3830
rect 2970 3820 2980 3830
rect 3280 3820 3850 3830
rect 4110 3820 4290 3830
rect 5260 3820 5980 3830
rect 7100 3820 8010 3830
rect 8020 3820 8070 3830
rect 8120 3820 8170 3830
rect 9610 3820 9730 3830
rect 0 3810 2600 3820
rect 2950 3810 2970 3820
rect 3280 3810 3860 3820
rect 4090 3810 4290 3820
rect 5270 3810 5970 3820
rect 7090 3810 8080 3820
rect 8090 3810 8100 3820
rect 8140 3810 8170 3820
rect 8630 3810 8640 3820
rect 9600 3810 9750 3820
rect 9780 3810 9810 3820
rect 0 3800 2620 3810
rect 3280 3800 3860 3810
rect 4070 3800 4290 3810
rect 5270 3800 5960 3810
rect 7080 3800 8020 3810
rect 8030 3800 8110 3810
rect 8150 3800 8180 3810
rect 9610 3800 9820 3810
rect 0 3790 2540 3800
rect 2560 3790 2600 3800
rect 2610 3790 2620 3800
rect 3290 3790 3870 3800
rect 4060 3790 4270 3800
rect 5280 3790 5970 3800
rect 7080 3790 8020 3800
rect 8030 3790 8110 3800
rect 8150 3790 8180 3800
rect 8250 3790 8260 3800
rect 8470 3790 8480 3800
rect 9620 3790 9750 3800
rect 9760 3790 9820 3800
rect 0 3780 2530 3790
rect 2570 3780 2620 3790
rect 3290 3780 3870 3790
rect 4050 3780 4240 3790
rect 5280 3780 5980 3790
rect 7070 3780 8020 3790
rect 8030 3780 8120 3790
rect 8160 3780 8190 3790
rect 8480 3780 8500 3790
rect 9620 3780 9740 3790
rect 9770 3780 9810 3790
rect 0 3770 1700 3780
rect 1720 3770 2540 3780
rect 2580 3770 2630 3780
rect 3280 3770 3290 3780
rect 3300 3770 3870 3780
rect 4040 3770 4220 3780
rect 5290 3770 6010 3780
rect 6050 3770 6060 3780
rect 7060 3770 8140 3780
rect 8160 3770 8180 3780
rect 9640 3770 9720 3780
rect 9770 3770 9800 3780
rect 0 3760 1680 3770
rect 1720 3760 2550 3770
rect 2590 3760 2640 3770
rect 3300 3760 3880 3770
rect 4020 3760 4180 3770
rect 5290 3760 6000 3770
rect 6010 3760 6020 3770
rect 7060 3760 8140 3770
rect 9660 3760 9710 3770
rect 9770 3760 9790 3770
rect 9820 3760 9860 3770
rect 0 3750 1660 3760
rect 1720 3750 2560 3760
rect 2600 3750 2650 3760
rect 2730 3750 2740 3760
rect 3300 3750 3880 3760
rect 4010 3750 4140 3760
rect 5300 3750 6020 3760
rect 7050 3750 8150 3760
rect 8360 3750 8370 3760
rect 9670 3750 9710 3760
rect 9730 3750 9750 3760
rect 9760 3750 9780 3760
rect 9830 3750 9850 3760
rect 0 3740 1640 3750
rect 1710 3740 2560 3750
rect 2600 3740 2670 3750
rect 3280 3740 3290 3750
rect 3310 3740 3880 3750
rect 4000 3740 4090 3750
rect 5300 3740 6040 3750
rect 7040 3740 8160 3750
rect 8350 3740 8380 3750
rect 9690 3740 9780 3750
rect 9830 3740 9850 3750
rect 0 3730 1630 3740
rect 1700 3730 2570 3740
rect 2600 3730 2680 3740
rect 2710 3730 2740 3740
rect 3310 3730 3880 3740
rect 3990 3730 4070 3740
rect 5300 3730 6070 3740
rect 7040 3730 8170 3740
rect 8350 3730 8380 3740
rect 9700 3730 9780 3740
rect 9800 3730 9810 3740
rect 0 3720 1610 3730
rect 1690 3720 2580 3730
rect 2590 3720 2770 3730
rect 3310 3720 3870 3730
rect 3990 3720 4050 3730
rect 5300 3720 6070 3730
rect 7030 3720 8170 3730
rect 9700 3720 9760 3730
rect 9800 3720 9820 3730
rect 9880 3720 9910 3730
rect 9920 3720 9960 3730
rect 0 3710 1620 3720
rect 1680 3710 2860 3720
rect 3310 3710 3870 3720
rect 3980 3710 4030 3720
rect 5310 3710 6070 3720
rect 7020 3710 8180 3720
rect 8580 3710 8600 3720
rect 9880 3710 9950 3720
rect 10 3700 1620 3710
rect 1710 3700 2870 3710
rect 3320 3700 3870 3710
rect 3970 3700 4010 3710
rect 5310 3700 6070 3710
rect 7020 3700 8190 3710
rect 8400 3700 8410 3710
rect 8580 3700 8610 3710
rect 9880 3700 9950 3710
rect 30 3690 1610 3700
rect 1690 3690 1700 3700
rect 1710 3690 2850 3700
rect 3320 3690 3870 3700
rect 3960 3690 4000 3700
rect 5310 3690 6070 3700
rect 7010 3690 8200 3700
rect 8400 3690 8450 3700
rect 8570 3690 8620 3700
rect 9890 3690 9930 3700
rect 30 3680 1610 3690
rect 1690 3680 2860 3690
rect 2870 3680 2910 3690
rect 2920 3680 3030 3690
rect 3330 3680 3870 3690
rect 3960 3680 3990 3690
rect 5320 3680 6070 3690
rect 7000 3680 8200 3690
rect 8410 3680 8450 3690
rect 8460 3680 8470 3690
rect 8570 3680 8610 3690
rect 9850 3680 9870 3690
rect 9880 3680 9920 3690
rect 40 3670 1610 3680
rect 1690 3670 1700 3680
rect 1710 3670 3040 3680
rect 3330 3670 3870 3680
rect 3940 3670 3980 3680
rect 5320 3670 6070 3680
rect 6990 3670 8200 3680
rect 8410 3670 8470 3680
rect 8570 3670 8590 3680
rect 9850 3670 9900 3680
rect 50 3660 1630 3670
rect 1650 3660 1660 3670
rect 1670 3660 1700 3670
rect 1720 3660 3070 3670
rect 3340 3660 3880 3670
rect 3940 3660 3970 3670
rect 5320 3660 6070 3670
rect 6990 3660 8200 3670
rect 8410 3660 8460 3670
rect 8470 3660 8480 3670
rect 8510 3660 8520 3670
rect 9860 3660 9880 3670
rect 0 3650 1690 3660
rect 1720 3650 3090 3660
rect 3340 3650 3960 3660
rect 5320 3650 6140 3660
rect 6980 3650 8210 3660
rect 8410 3650 8530 3660
rect 0 3640 1670 3650
rect 1690 3640 1700 3650
rect 1710 3640 3070 3650
rect 3120 3640 3130 3650
rect 3350 3640 3950 3650
rect 5330 3640 6150 3650
rect 6970 3640 8220 3650
rect 8410 3640 8510 3650
rect 8520 3640 8530 3650
rect 0 3630 1640 3640
rect 1650 3630 1700 3640
rect 1710 3630 3150 3640
rect 3350 3630 3950 3640
rect 5330 3630 6160 3640
rect 6960 3630 8230 3640
rect 8390 3630 8410 3640
rect 8430 3630 8500 3640
rect 9880 3630 9890 3640
rect 0 3620 1690 3630
rect 1710 3620 3170 3630
rect 3360 3620 3940 3630
rect 5330 3620 6170 3630
rect 6960 3620 8250 3630
rect 8390 3620 8410 3630
rect 8430 3620 8490 3630
rect 9910 3620 9920 3630
rect 0 3610 1680 3620
rect 1690 3610 1700 3620
rect 1710 3610 3170 3620
rect 3360 3610 3930 3620
rect 5330 3610 6180 3620
rect 6950 3610 8260 3620
rect 8390 3610 8500 3620
rect 9910 3610 9930 3620
rect 0 3600 1490 3610
rect 1500 3600 1690 3610
rect 1720 3600 3210 3610
rect 3370 3600 3920 3610
rect 5330 3600 6190 3610
rect 6940 3600 8260 3610
rect 8380 3600 8410 3610
rect 8430 3600 8500 3610
rect 9920 3600 9940 3610
rect 0 3590 1480 3600
rect 1490 3590 1700 3600
rect 1710 3590 3230 3600
rect 3370 3590 3910 3600
rect 5340 3590 6180 3600
rect 6930 3590 8280 3600
rect 8440 3590 8490 3600
rect 0 3580 1470 3590
rect 1490 3580 1690 3590
rect 1720 3580 3240 3590
rect 3370 3580 3910 3590
rect 5340 3580 6180 3590
rect 6920 3580 8300 3590
rect 8450 3580 8490 3590
rect 0 3570 1470 3580
rect 1480 3570 1690 3580
rect 1710 3570 3240 3580
rect 3380 3570 3900 3580
rect 5340 3570 6180 3580
rect 6920 3570 8310 3580
rect 8420 3570 8430 3580
rect 8460 3570 8480 3580
rect 0 3560 1460 3570
rect 1480 3560 1680 3570
rect 1710 3560 3250 3570
rect 3380 3560 3900 3570
rect 5340 3560 6180 3570
rect 6910 3560 8320 3570
rect 8420 3560 8440 3570
rect 8470 3560 8490 3570
rect 0 3550 1450 3560
rect 1480 3550 1690 3560
rect 1700 3550 3260 3560
rect 3390 3550 3900 3560
rect 4750 3550 4760 3560
rect 5340 3550 6170 3560
rect 6900 3550 8320 3560
rect 8420 3550 8440 3560
rect 8460 3550 8490 3560
rect 0 3540 1450 3550
rect 1480 3540 1690 3550
rect 1700 3540 3270 3550
rect 3390 3540 3900 3550
rect 4740 3540 4750 3550
rect 5340 3540 6170 3550
rect 6890 3540 8330 3550
rect 8450 3540 8480 3550
rect 0 3530 1440 3540
rect 1480 3530 1690 3540
rect 1700 3530 2710 3540
rect 2720 3530 3280 3540
rect 3400 3530 3910 3540
rect 5340 3530 6170 3540
rect 6880 3530 8340 3540
rect 8450 3530 8480 3540
rect 0 3520 1430 3530
rect 1480 3520 1690 3530
rect 1700 3520 3280 3530
rect 3400 3520 3920 3530
rect 5340 3520 6160 3530
rect 6880 3520 8340 3530
rect 8470 3520 8490 3530
rect 0 3510 1430 3520
rect 1470 3510 2570 3520
rect 2580 3510 3290 3520
rect 3320 3510 3330 3520
rect 3410 3510 3920 3520
rect 5340 3510 6160 3520
rect 6870 3510 8350 3520
rect 8470 3510 8490 3520
rect 0 3500 1420 3510
rect 1470 3500 2500 3510
rect 2600 3500 3300 3510
rect 3320 3500 3350 3510
rect 3410 3500 3920 3510
rect 5340 3500 6160 3510
rect 6860 3500 8350 3510
rect 8450 3500 8480 3510
rect 0 3490 1420 3500
rect 1470 3490 2440 3500
rect 2680 3490 3310 3500
rect 3330 3490 3360 3500
rect 3410 3490 3920 3500
rect 5010 3490 5040 3500
rect 5340 3490 6160 3500
rect 6850 3490 8350 3500
rect 8380 3490 8390 3500
rect 8460 3490 8510 3500
rect 9350 3490 9360 3500
rect 0 3480 1410 3490
rect 1460 3480 2390 3490
rect 2400 3480 2410 3490
rect 2760 3480 3310 3490
rect 3360 3480 3370 3490
rect 3420 3480 3920 3490
rect 4990 3480 5040 3490
rect 5340 3480 6160 3490
rect 6850 3480 8360 3490
rect 8380 3480 8400 3490
rect 8480 3480 8520 3490
rect 9280 3480 9340 3490
rect 0 3470 1410 3480
rect 1460 3470 2370 3480
rect 2810 3470 3320 3480
rect 3360 3470 3380 3480
rect 3420 3470 3920 3480
rect 4970 3470 5040 3480
rect 5340 3470 6150 3480
rect 6840 3470 8420 3480
rect 8490 3470 8530 3480
rect 9270 3470 9310 3480
rect 0 3460 1400 3470
rect 1450 3460 2350 3470
rect 2820 3460 3340 3470
rect 3390 3460 3400 3470
rect 3440 3460 3920 3470
rect 4950 3460 5030 3470
rect 5340 3460 6140 3470
rect 6830 3460 8420 3470
rect 8490 3460 8530 3470
rect 9260 3460 9290 3470
rect 0 3450 1400 3460
rect 1450 3450 2300 3460
rect 2310 3450 2320 3460
rect 2870 3450 3350 3460
rect 3400 3450 3410 3460
rect 3440 3450 3920 3460
rect 4520 3450 4590 3460
rect 4940 3450 5030 3460
rect 5340 3450 5870 3460
rect 5880 3450 6140 3460
rect 6820 3450 8430 3460
rect 8490 3450 8520 3460
rect 9240 3450 9270 3460
rect 0 3440 1390 3450
rect 1450 3440 2280 3450
rect 2900 3440 3380 3450
rect 3390 3440 3430 3450
rect 3450 3440 3930 3450
rect 4480 3440 4610 3450
rect 4930 3440 5020 3450
rect 5340 3440 5850 3450
rect 5890 3440 5900 3450
rect 5910 3440 5940 3450
rect 5950 3440 5960 3450
rect 5970 3440 6140 3450
rect 6810 3440 8450 3450
rect 8500 3440 8520 3450
rect 9220 3440 9260 3450
rect 0 3430 1390 3440
rect 1450 3430 2270 3440
rect 2940 3430 3440 3440
rect 3450 3430 3930 3440
rect 4460 3430 4560 3440
rect 4910 3430 5020 3440
rect 5340 3430 5850 3440
rect 5990 3430 6020 3440
rect 6030 3430 6130 3440
rect 6800 3430 8450 3440
rect 8510 3430 8540 3440
rect 9210 3430 9240 3440
rect 0 3420 1380 3430
rect 1450 3420 2240 3430
rect 2960 3420 3410 3430
rect 3420 3420 3940 3430
rect 4440 3420 4510 3430
rect 4900 3420 4970 3430
rect 4990 3420 5020 3430
rect 5340 3420 5860 3430
rect 6020 3420 6050 3430
rect 6060 3420 6130 3430
rect 6790 3420 8490 3430
rect 8510 3420 8540 3430
rect 9190 3420 9230 3430
rect 0 3410 1380 3420
rect 1440 3410 2230 3420
rect 2970 3410 3940 3420
rect 4880 3410 4940 3420
rect 5000 3410 5020 3420
rect 5340 3410 5840 3420
rect 6020 3410 6040 3420
rect 6060 3410 6130 3420
rect 6770 3410 8490 3420
rect 8510 3410 8530 3420
rect 9180 3410 9210 3420
rect 0 3400 1370 3410
rect 1440 3400 2210 3410
rect 2990 3400 3950 3410
rect 4860 3400 4920 3410
rect 5010 3400 5020 3410
rect 5330 3400 5680 3410
rect 5690 3400 5860 3410
rect 6060 3400 6130 3410
rect 6760 3400 8500 3410
rect 8510 3400 8520 3410
rect 9110 3400 9200 3410
rect 0 3390 1370 3400
rect 1430 3390 2190 3400
rect 3010 3390 3950 3400
rect 4300 3390 4310 3400
rect 4850 3390 4910 3400
rect 5330 3390 5680 3400
rect 5710 3390 5850 3400
rect 6050 3390 6140 3400
rect 6750 3390 8500 3400
rect 9110 3390 9190 3400
rect 0 3380 1360 3390
rect 1430 3380 2180 3390
rect 3040 3380 3490 3390
rect 3520 3380 3960 3390
rect 4290 3380 4300 3390
rect 4830 3380 4900 3390
rect 5330 3380 5680 3390
rect 5730 3380 5850 3390
rect 6040 3380 6140 3390
rect 6740 3380 8500 3390
rect 9120 3380 9180 3390
rect 0 3370 1360 3380
rect 1420 3370 2160 3380
rect 3040 3370 3490 3380
rect 3540 3370 3960 3380
rect 4290 3370 4300 3380
rect 4800 3370 4890 3380
rect 5330 3370 5630 3380
rect 5650 3370 5670 3380
rect 5740 3370 5830 3380
rect 5840 3370 5850 3380
rect 6050 3370 6140 3380
rect 6730 3370 8500 3380
rect 9120 3370 9170 3380
rect 0 3360 1360 3370
rect 1420 3360 2160 3370
rect 3060 3360 3490 3370
rect 3550 3360 3970 3370
rect 4280 3360 4300 3370
rect 4790 3360 4880 3370
rect 5330 3360 5640 3370
rect 5740 3360 5850 3370
rect 6050 3360 6130 3370
rect 6720 3360 8500 3370
rect 9120 3360 9160 3370
rect 9740 3360 9810 3370
rect 0 3350 1350 3360
rect 1410 3350 2160 3360
rect 3070 3350 3480 3360
rect 3560 3350 3960 3360
rect 4280 3350 4290 3360
rect 4780 3350 4870 3360
rect 5330 3350 5640 3360
rect 5760 3350 5850 3360
rect 6050 3350 6130 3360
rect 6700 3350 8500 3360
rect 9100 3350 9150 3360
rect 9730 3350 9810 3360
rect 0 3340 1350 3350
rect 1410 3340 2140 3350
rect 3080 3340 3480 3350
rect 3580 3340 3970 3350
rect 4270 3340 4290 3350
rect 4760 3340 4850 3350
rect 5320 3340 5630 3350
rect 5760 3340 5850 3350
rect 6080 3340 6130 3350
rect 6700 3340 8490 3350
rect 9090 3340 9140 3350
rect 9730 3340 9790 3350
rect 0 3330 1340 3340
rect 1410 3330 2120 3340
rect 3100 3330 3490 3340
rect 3590 3330 3980 3340
rect 4270 3330 4280 3340
rect 4750 3330 4790 3340
rect 4820 3330 4840 3340
rect 5320 3330 5620 3340
rect 5770 3330 5850 3340
rect 6060 3330 6130 3340
rect 6680 3330 8490 3340
rect 9060 3330 9130 3340
rect 9760 3330 9790 3340
rect 0 3320 1340 3330
rect 1410 3320 2120 3330
rect 3110 3320 3500 3330
rect 3590 3320 3980 3330
rect 4270 3320 4280 3330
rect 4740 3320 4770 3330
rect 4810 3320 4840 3330
rect 5320 3320 5620 3330
rect 5780 3320 5840 3330
rect 6080 3320 6130 3330
rect 6680 3320 8490 3330
rect 9070 3320 9130 3330
rect 9720 3320 9730 3330
rect 9760 3320 9780 3330
rect 0 3310 1330 3320
rect 1400 3310 2110 3320
rect 3120 3310 3500 3320
rect 3520 3310 3530 3320
rect 3590 3310 3990 3320
rect 4260 3310 4280 3320
rect 4670 3310 4690 3320
rect 4720 3310 4750 3320
rect 5320 3310 5620 3320
rect 5780 3310 5840 3320
rect 6000 3310 6010 3320
rect 6090 3310 6120 3320
rect 6680 3310 8490 3320
rect 9080 3310 9120 3320
rect 9710 3310 9740 3320
rect 0 3300 1330 3310
rect 1400 3300 2100 3310
rect 3120 3300 3510 3310
rect 3590 3300 3990 3310
rect 4650 3300 4740 3310
rect 5310 3300 5620 3310
rect 5790 3300 5820 3310
rect 6680 3300 8480 3310
rect 9080 3300 9110 3310
rect 9710 3300 9730 3310
rect 9740 3300 9760 3310
rect 0 3290 1320 3300
rect 1400 3290 2100 3300
rect 3130 3290 3520 3300
rect 3580 3290 4000 3300
rect 4600 3290 4740 3300
rect 5310 3290 5620 3300
rect 5790 3290 5800 3300
rect 6670 3290 8470 3300
rect 9070 3290 9090 3300
rect 9700 3290 9710 3300
rect 9740 3290 9750 3300
rect 0 3280 1320 3290
rect 1390 3280 2090 3290
rect 3140 3280 3530 3290
rect 3540 3280 3560 3290
rect 3600 3280 4010 3290
rect 4580 3280 4690 3290
rect 5310 3280 5620 3290
rect 6670 3280 8470 3290
rect 0 3270 1320 3280
rect 1390 3270 2080 3280
rect 3150 3270 3570 3280
rect 3590 3270 4020 3280
rect 4530 3270 4690 3280
rect 5310 3270 5620 3280
rect 6670 3270 8470 3280
rect 9990 3270 9990 3280
rect 0 3260 1310 3270
rect 1390 3260 2070 3270
rect 3130 3260 3140 3270
rect 3150 3260 3570 3270
rect 3600 3260 4030 3270
rect 4470 3260 4650 3270
rect 5300 3260 5630 3270
rect 6560 3260 6590 3270
rect 6670 3260 8460 3270
rect 9650 3260 9680 3270
rect 9980 3260 9990 3270
rect 0 3250 1310 3260
rect 1380 3250 2070 3260
rect 3160 3250 3570 3260
rect 3600 3250 4030 3260
rect 4440 3250 4630 3260
rect 5300 3250 5630 3260
rect 6540 3250 6590 3260
rect 6660 3250 8460 3260
rect 9390 3250 9410 3260
rect 9640 3250 9690 3260
rect 9960 3250 9990 3260
rect 0 3240 1300 3250
rect 1380 3240 2060 3250
rect 3170 3240 3570 3250
rect 3610 3240 4040 3250
rect 4420 3240 4600 3250
rect 5300 3240 5640 3250
rect 6520 3240 6580 3250
rect 6660 3240 8450 3250
rect 9110 3240 9120 3250
rect 9380 3240 9400 3250
rect 9630 3240 9670 3250
rect 9960 3240 9990 3250
rect 0 3230 1300 3240
rect 1380 3230 2060 3240
rect 3150 3230 3580 3240
rect 3620 3230 4050 3240
rect 4380 3230 4620 3240
rect 4950 3230 4960 3240
rect 5300 3230 5630 3240
rect 6500 3230 6580 3240
rect 6660 3230 8450 3240
rect 9100 3230 9120 3240
rect 9370 3230 9380 3240
rect 9980 3230 9990 3240
rect 0 3220 1290 3230
rect 1370 3220 2060 3230
rect 3160 3220 3560 3230
rect 3570 3220 3580 3230
rect 3620 3220 4050 3230
rect 4370 3220 4630 3230
rect 5290 3220 5650 3230
rect 6480 3220 6580 3230
rect 6660 3220 8440 3230
rect 9090 3220 9130 3230
rect 0 3210 1290 3220
rect 1370 3210 2060 3220
rect 3160 3210 3590 3220
rect 3620 3210 4070 3220
rect 4360 3210 4580 3220
rect 4940 3210 4950 3220
rect 4960 3210 4970 3220
rect 5290 3210 5650 3220
rect 6470 3210 6580 3220
rect 6660 3210 8440 3220
rect 9080 3210 9140 3220
rect 9350 3210 9360 3220
rect 9950 3210 9960 3220
rect 0 3200 1290 3210
rect 1360 3200 2050 3210
rect 3170 3200 3600 3210
rect 3610 3200 4060 3210
rect 4350 3200 4520 3210
rect 4930 3200 4960 3210
rect 5290 3200 5670 3210
rect 6450 3200 6580 3210
rect 6660 3200 8430 3210
rect 9080 3200 9150 3210
rect 9340 3200 9360 3210
rect 0 3190 1280 3200
rect 1360 3190 2040 3200
rect 3170 3190 4070 3200
rect 4340 3190 4490 3200
rect 4920 3190 4960 3200
rect 5280 3190 5690 3200
rect 6420 3190 6580 3200
rect 6650 3190 8430 3200
rect 9060 3190 9170 3200
rect 9330 3190 9360 3200
rect 9570 3190 9580 3200
rect 9910 3190 9920 3200
rect 0 3180 1280 3190
rect 1360 3180 2040 3190
rect 3170 3180 4060 3190
rect 4110 3180 4120 3190
rect 4350 3180 4470 3190
rect 4910 3180 4950 3190
rect 5280 3180 5710 3190
rect 6390 3180 6580 3190
rect 6650 3180 8430 3190
rect 9060 3180 9190 3190
rect 9330 3180 9350 3190
rect 9910 3180 9940 3190
rect 0 3170 1270 3180
rect 1350 3170 2030 3180
rect 3180 3170 4070 3180
rect 4380 3170 4460 3180
rect 4920 3170 4940 3180
rect 5280 3170 5720 3180
rect 6360 3170 6580 3180
rect 6650 3170 8420 3180
rect 9110 3170 9220 3180
rect 9590 3170 9620 3180
rect 9900 3170 9940 3180
rect 0 3160 1270 3170
rect 1350 3160 2030 3170
rect 3180 3160 4070 3170
rect 4400 3160 4460 3170
rect 4900 3160 4930 3170
rect 5270 3160 5740 3170
rect 6320 3160 6570 3170
rect 6650 3160 8420 3170
rect 9100 3160 9250 3170
rect 9600 3160 9620 3170
rect 9900 3160 9930 3170
rect 9940 3160 9960 3170
rect 0 3150 1270 3160
rect 1350 3150 2030 3160
rect 3180 3150 3750 3160
rect 3760 3150 4070 3160
rect 4420 3150 4460 3160
rect 4900 3150 4920 3160
rect 5270 3150 5770 3160
rect 6290 3150 6570 3160
rect 6650 3150 8410 3160
rect 9100 3150 9260 3160
rect 9600 3150 9620 3160
rect 9900 3150 9920 3160
rect 9930 3150 9970 3160
rect 0 3140 1260 3150
rect 1340 3140 2030 3150
rect 3190 3140 3720 3150
rect 3730 3140 3740 3150
rect 3780 3140 4070 3150
rect 4440 3140 4460 3150
rect 4890 3140 4910 3150
rect 5270 3140 5800 3150
rect 6200 3140 6210 3150
rect 6220 3140 6570 3150
rect 6640 3140 8410 3150
rect 9100 3140 9250 3150
rect 9930 3140 9990 3150
rect 0 3130 1260 3140
rect 1340 3130 2030 3140
rect 3190 3130 3720 3140
rect 3740 3130 3760 3140
rect 3790 3130 4080 3140
rect 4450 3130 4470 3140
rect 4880 3130 4900 3140
rect 5260 3130 5850 3140
rect 6170 3130 6570 3140
rect 6640 3130 8400 3140
rect 9100 3130 9210 3140
rect 9860 3130 9870 3140
rect 9930 3130 9990 3140
rect 0 3120 1250 3130
rect 1340 3120 2030 3130
rect 3190 3120 3720 3130
rect 3730 3120 3770 3130
rect 3830 3120 4080 3130
rect 4160 3120 4170 3130
rect 4470 3120 4490 3130
rect 4860 3120 4890 3130
rect 5260 3120 5910 3130
rect 6060 3120 6080 3130
rect 6090 3120 6100 3130
rect 6110 3120 6570 3130
rect 6640 3120 8390 3130
rect 9100 3120 9200 3130
rect 9450 3120 9460 3130
rect 9860 3120 9870 3130
rect 9940 3120 9990 3130
rect 0 3110 1250 3120
rect 1340 3110 2020 3120
rect 3190 3110 3770 3120
rect 3830 3110 3860 3120
rect 3890 3110 4030 3120
rect 4040 3110 4090 3120
rect 4160 3110 4170 3120
rect 4480 3110 4500 3120
rect 4850 3110 4880 3120
rect 5260 3110 6570 3120
rect 6630 3110 8380 3120
rect 9100 3110 9200 3120
rect 9440 3110 9460 3120
rect 9840 3110 9850 3120
rect 9860 3110 9880 3120
rect 9950 3110 9990 3120
rect 0 3100 1250 3110
rect 1340 3100 2020 3110
rect 3190 3100 3790 3110
rect 3830 3100 3850 3110
rect 3900 3100 4100 3110
rect 4170 3100 4180 3110
rect 4490 3100 4520 3110
rect 4840 3100 4870 3110
rect 5250 3100 6560 3110
rect 6630 3100 8380 3110
rect 9100 3100 9200 3110
rect 9440 3100 9460 3110
rect 9830 3100 9870 3110
rect 9960 3100 9990 3110
rect 0 3090 1240 3100
rect 1330 3090 2020 3100
rect 3190 3090 3780 3100
rect 3820 3090 3850 3100
rect 3940 3090 4040 3100
rect 4050 3090 4100 3100
rect 4190 3090 4200 3100
rect 4500 3090 4550 3100
rect 4820 3090 4870 3100
rect 5250 3090 6560 3100
rect 6630 3090 8380 3100
rect 9100 3090 9200 3100
rect 9440 3090 9460 3100
rect 9830 3090 9870 3100
rect 9990 3090 9990 3100
rect 0 3080 1240 3090
rect 1330 3080 2020 3090
rect 3200 3080 3660 3090
rect 3670 3080 3780 3090
rect 3950 3080 4110 3090
rect 4520 3080 4570 3090
rect 4810 3080 4850 3090
rect 5240 3080 6560 3090
rect 6630 3080 8380 3090
rect 8400 3080 8430 3090
rect 9090 3080 9210 3090
rect 9440 3080 9460 3090
rect 9810 3080 9890 3090
rect 9950 3080 9960 3090
rect 0 3070 1230 3080
rect 1320 3070 2010 3080
rect 3200 3070 3780 3080
rect 3990 3070 4120 3080
rect 4200 3070 4220 3080
rect 4530 3070 4610 3080
rect 4760 3070 4830 3080
rect 5240 3070 6560 3080
rect 6630 3070 8370 3080
rect 8400 3070 8420 3080
rect 9080 3070 9220 3080
rect 9450 3070 9470 3080
rect 9800 3070 9890 3080
rect 0 3060 1230 3070
rect 1320 3060 2010 3070
rect 3190 3060 3760 3070
rect 4030 3060 4060 3070
rect 4070 3060 4130 3070
rect 4220 3060 4230 3070
rect 4550 3060 4690 3070
rect 4700 3060 4710 3070
rect 4720 3060 4810 3070
rect 5230 3060 6560 3070
rect 6630 3060 8370 3070
rect 8400 3060 8410 3070
rect 9090 3060 9230 3070
rect 9460 3060 9480 3070
rect 9800 3060 9890 3070
rect 0 3050 1230 3060
rect 1320 3050 2010 3060
rect 3190 3050 3740 3060
rect 4030 3050 4140 3060
rect 4220 3050 4240 3060
rect 4570 3050 4800 3060
rect 5230 3050 6560 3060
rect 6620 3050 8360 3060
rect 9090 3050 9250 3060
rect 9790 3050 9890 3060
rect 0 3040 1220 3050
rect 1310 3040 2010 3050
rect 3190 3040 3740 3050
rect 4030 3040 4040 3050
rect 4050 3040 4140 3050
rect 4590 3040 4780 3050
rect 5230 3040 6550 3050
rect 6610 3040 8360 3050
rect 9080 3040 9240 3050
rect 9780 3040 9830 3050
rect 9840 3040 9890 3050
rect 0 3030 1220 3040
rect 1310 3030 2010 3040
rect 3190 3030 3740 3040
rect 4040 3030 4160 3040
rect 4630 3030 4750 3040
rect 5220 3030 6550 3040
rect 6610 3030 8350 3040
rect 9080 3030 9230 3040
rect 9780 3030 9900 3040
rect 0 3020 1210 3030
rect 1310 3020 2010 3030
rect 3200 3020 3740 3030
rect 3850 3020 3860 3030
rect 4040 3020 4090 3030
rect 4100 3020 4160 3030
rect 5220 3020 6550 3030
rect 6620 3020 8350 3030
rect 9080 3020 9140 3030
rect 9150 3020 9220 3030
rect 9760 3020 9900 3030
rect 0 3010 1210 3020
rect 1300 3010 2010 3020
rect 3200 3010 3730 3020
rect 3800 3010 3820 3020
rect 3850 3010 3860 3020
rect 4050 3010 4100 3020
rect 4110 3010 4180 3020
rect 5210 3010 6550 3020
rect 6610 3010 8340 3020
rect 8410 3010 8430 3020
rect 9080 3010 9130 3020
rect 9170 3010 9210 3020
rect 9760 3010 9790 3020
rect 9890 3010 9900 3020
rect 0 3000 1200 3010
rect 1300 3000 2010 3010
rect 3200 3000 3740 3010
rect 3790 3000 3810 3010
rect 4070 3000 4190 3010
rect 5210 3000 6550 3010
rect 6610 3000 8340 3010
rect 8410 3000 8440 3010
rect 9080 3000 9130 3010
rect 9180 3000 9200 3010
rect 0 2990 1200 3000
rect 1300 2990 2010 3000
rect 3200 2990 3770 3000
rect 3780 2990 3790 3000
rect 3800 2990 3820 3000
rect 3840 2990 3860 3000
rect 4020 2990 4050 3000
rect 4070 2990 4200 3000
rect 5200 2990 6550 3000
rect 6610 2990 8330 3000
rect 8410 2990 8440 3000
rect 9090 2990 9120 3000
rect 9180 2990 9200 3000
rect 0 2980 1200 2990
rect 1300 2980 2000 2990
rect 3200 2980 3860 2990
rect 4010 2980 4050 2990
rect 4070 2980 4080 2990
rect 4100 2980 4210 2990
rect 5200 2980 6550 2990
rect 6610 2980 8330 2990
rect 8410 2980 8440 2990
rect 9080 2980 9120 2990
rect 0 2970 1190 2980
rect 1290 2970 2000 2980
rect 3200 2970 3860 2980
rect 3870 2970 3880 2980
rect 4010 2970 4040 2980
rect 4110 2970 4140 2980
rect 4150 2970 4230 2980
rect 5190 2970 6550 2980
rect 6600 2970 8320 2980
rect 8410 2970 8440 2980
rect 9080 2970 9110 2980
rect 0 2960 1190 2970
rect 1290 2960 2000 2970
rect 3190 2960 3790 2970
rect 3800 2960 3880 2970
rect 4010 2960 4040 2970
rect 4120 2960 4150 2970
rect 4160 2960 4250 2970
rect 5190 2960 6550 2970
rect 6600 2960 8310 2970
rect 8410 2960 8450 2970
rect 9070 2960 9110 2970
rect 0 2950 1180 2960
rect 1280 2950 2000 2960
rect 3170 2950 3780 2960
rect 3810 2950 3850 2960
rect 3860 2950 3890 2960
rect 4010 2950 4050 2960
rect 4140 2950 4150 2960
rect 4170 2950 4250 2960
rect 5180 2950 6540 2960
rect 6600 2950 8310 2960
rect 9070 2950 9100 2960
rect 0 2940 1180 2950
rect 1280 2940 2000 2950
rect 3170 2940 3820 2950
rect 3880 2940 3890 2950
rect 3980 2940 4000 2950
rect 4020 2940 4050 2950
rect 4180 2940 4270 2950
rect 5180 2940 6540 2950
rect 6600 2940 8300 2950
rect 9070 2940 9100 2950
rect 0 2930 1180 2940
rect 1280 2930 2000 2940
rect 3170 2930 3810 2940
rect 3880 2930 3900 2940
rect 3970 2930 4000 2940
rect 4020 2930 4040 2940
rect 4190 2930 4280 2940
rect 5180 2930 6540 2940
rect 6590 2930 8300 2940
rect 9060 2930 9090 2940
rect 9710 2930 9730 2940
rect 0 2920 1170 2930
rect 1270 2920 2000 2930
rect 3160 2920 3810 2930
rect 3860 2920 3910 2930
rect 3960 2920 3990 2930
rect 4010 2920 4030 2930
rect 4210 2920 4290 2930
rect 5170 2920 6540 2930
rect 6590 2920 8290 2930
rect 9060 2920 9090 2930
rect 9720 2920 9730 2930
rect 0 2910 1170 2920
rect 1260 2910 2000 2920
rect 3160 2910 3810 2920
rect 3850 2910 3880 2920
rect 3890 2910 3990 2920
rect 4000 2910 4020 2920
rect 4220 2910 4310 2920
rect 5170 2910 6540 2920
rect 6590 2910 8280 2920
rect 9060 2910 9080 2920
rect 0 2900 1160 2910
rect 1260 2900 2000 2910
rect 3160 2900 3780 2910
rect 3790 2900 3880 2910
rect 3910 2900 3920 2910
rect 3950 2900 4010 2910
rect 4230 2900 4330 2910
rect 5160 2900 6540 2910
rect 6590 2900 8270 2910
rect 9060 2900 9070 2910
rect 9990 2900 9990 2910
rect 0 2890 1160 2900
rect 1250 2890 1990 2900
rect 3160 2890 3890 2900
rect 3900 2890 3920 2900
rect 3950 2890 4010 2900
rect 4240 2890 4350 2900
rect 5170 2890 6540 2900
rect 6590 2890 8270 2900
rect 9990 2890 9990 2900
rect 0 2880 1160 2890
rect 1250 2880 1990 2890
rect 3160 2880 3590 2890
rect 3600 2880 3890 2890
rect 3900 2880 4000 2890
rect 4250 2880 4360 2890
rect 5170 2880 6540 2890
rect 6580 2880 8260 2890
rect 0 2870 1150 2880
rect 1250 2870 1990 2880
rect 3160 2870 3600 2880
rect 3610 2870 3850 2880
rect 3870 2870 3890 2880
rect 3900 2870 3990 2880
rect 4260 2870 4380 2880
rect 5170 2870 6540 2880
rect 6590 2870 8250 2880
rect 0 2860 1150 2870
rect 1240 2860 1990 2870
rect 3160 2860 3860 2870
rect 3900 2860 3910 2870
rect 3920 2860 3990 2870
rect 4250 2860 4400 2870
rect 5170 2860 6530 2870
rect 6580 2860 7420 2870
rect 7490 2860 8250 2870
rect 9990 2860 9990 2870
rect 0 2850 1140 2860
rect 1230 2850 1990 2860
rect 3160 2850 3810 2860
rect 3830 2850 3860 2860
rect 3880 2850 3900 2860
rect 3940 2850 3980 2860
rect 4250 2850 4410 2860
rect 5170 2850 6530 2860
rect 6570 2850 7270 2860
rect 7350 2850 7380 2860
rect 7510 2850 8240 2860
rect 0 2840 1140 2850
rect 1230 2840 1990 2850
rect 3160 2840 3860 2850
rect 3870 2840 3900 2850
rect 3940 2840 3980 2850
rect 4250 2840 4430 2850
rect 5170 2840 6530 2850
rect 6570 2840 7250 2850
rect 7520 2840 8230 2850
rect 0 2830 1130 2840
rect 1230 2830 1990 2840
rect 3160 2830 3890 2840
rect 3900 2830 3920 2840
rect 3930 2830 3980 2840
rect 4260 2830 4450 2840
rect 5170 2830 6530 2840
rect 6570 2830 7230 2840
rect 7530 2830 8220 2840
rect 9370 2830 9380 2840
rect 0 2820 1130 2830
rect 1230 2820 1990 2830
rect 3160 2820 3910 2830
rect 3930 2820 3960 2830
rect 3970 2820 3980 2830
rect 4260 2820 4460 2830
rect 5170 2820 6530 2830
rect 6570 2820 7210 2830
rect 7540 2820 8210 2830
rect 9370 2820 9410 2830
rect 0 2810 1120 2820
rect 1220 2810 1990 2820
rect 3160 2810 3980 2820
rect 4260 2810 4480 2820
rect 5170 2810 5840 2820
rect 5850 2810 5870 2820
rect 5880 2810 5910 2820
rect 6080 2810 6530 2820
rect 6570 2810 7190 2820
rect 7550 2810 8210 2820
rect 9380 2810 9420 2820
rect 0 2800 1120 2810
rect 1210 2800 1980 2810
rect 3150 2800 3960 2810
rect 4260 2800 4490 2810
rect 5170 2800 5790 2810
rect 5820 2800 5830 2810
rect 6110 2800 6520 2810
rect 6570 2800 7180 2810
rect 7560 2800 8200 2810
rect 9400 2800 9450 2810
rect 9560 2800 9580 2810
rect 0 2790 1120 2800
rect 1210 2790 1980 2800
rect 3150 2790 3970 2800
rect 4270 2790 4500 2800
rect 5170 2790 5740 2800
rect 6120 2790 6530 2800
rect 6560 2790 7160 2800
rect 7570 2790 8190 2800
rect 9420 2790 9470 2800
rect 9580 2790 9590 2800
rect 9930 2790 9940 2800
rect 0 2780 1110 2790
rect 1210 2780 1980 2790
rect 3150 2780 3950 2790
rect 4270 2780 4520 2790
rect 5180 2780 5560 2790
rect 5680 2780 5700 2790
rect 5760 2780 5770 2790
rect 6130 2780 6520 2790
rect 6560 2780 7150 2790
rect 7590 2780 8180 2790
rect 8850 2780 8870 2790
rect 9430 2780 9480 2790
rect 9930 2780 9960 2790
rect 0 2770 1110 2780
rect 1200 2770 1990 2780
rect 3150 2770 3860 2780
rect 3870 2770 3900 2780
rect 3910 2770 3940 2780
rect 4270 2770 4540 2780
rect 5170 2770 5550 2780
rect 6130 2770 6520 2780
rect 6550 2770 7140 2780
rect 7610 2770 8170 2780
rect 8780 2770 8860 2780
rect 9460 2770 9500 2780
rect 9640 2770 9670 2780
rect 9930 2770 9980 2780
rect 0 2760 1100 2770
rect 1190 2760 1980 2770
rect 3160 2760 3860 2770
rect 4270 2760 4560 2770
rect 5180 2760 5540 2770
rect 6130 2760 6530 2770
rect 6560 2760 7120 2770
rect 7620 2760 8170 2770
rect 8750 2760 8850 2770
rect 9480 2760 9520 2770
rect 9630 2760 9680 2770
rect 9930 2760 9990 2770
rect 0 2750 1100 2760
rect 1190 2750 1980 2760
rect 3160 2750 3920 2760
rect 4270 2750 4590 2760
rect 5180 2750 5530 2760
rect 6130 2750 6520 2760
rect 6550 2750 7100 2760
rect 7630 2750 8160 2760
rect 8740 2750 8840 2760
rect 9410 2750 9420 2760
rect 9500 2750 9530 2760
rect 9640 2750 9690 2760
rect 9920 2750 9990 2760
rect 0 2740 1090 2750
rect 1180 2740 1980 2750
rect 3160 2740 3920 2750
rect 4270 2740 4620 2750
rect 5180 2740 5520 2750
rect 6130 2740 6520 2750
rect 6550 2740 7070 2750
rect 7640 2740 8150 2750
rect 8730 2740 8800 2750
rect 9410 2740 9420 2750
rect 9530 2740 9560 2750
rect 9640 2740 9710 2750
rect 9920 2740 9990 2750
rect 0 2730 1090 2740
rect 1180 2730 1980 2740
rect 3160 2730 3880 2740
rect 3900 2730 3910 2740
rect 4270 2730 4670 2740
rect 5180 2730 5510 2740
rect 6140 2730 6520 2740
rect 6550 2730 7050 2740
rect 7640 2730 8140 2740
rect 8740 2730 8770 2740
rect 8860 2730 8890 2740
rect 9400 2730 9410 2740
rect 9550 2730 9580 2740
rect 9640 2730 9690 2740
rect 9920 2730 9990 2740
rect 0 2720 1080 2730
rect 1170 2720 1970 2730
rect 3160 2720 3880 2730
rect 4270 2720 4690 2730
rect 4700 2720 4710 2730
rect 5190 2720 5310 2730
rect 5340 2720 5500 2730
rect 6150 2720 6520 2730
rect 6550 2720 7030 2730
rect 7650 2720 8140 2730
rect 8740 2720 8750 2730
rect 9400 2720 9410 2730
rect 9570 2720 9600 2730
rect 9650 2720 9690 2730
rect 9920 2720 9990 2730
rect 0 2710 1080 2720
rect 1150 2710 1980 2720
rect 3160 2710 3890 2720
rect 4270 2710 4730 2720
rect 5190 2710 5240 2720
rect 5370 2710 5490 2720
rect 6160 2710 6510 2720
rect 6540 2710 7010 2720
rect 7660 2710 8130 2720
rect 9380 2710 9400 2720
rect 9590 2710 9620 2720
rect 9940 2710 9990 2720
rect 0 2700 1070 2710
rect 1140 2700 1980 2710
rect 3160 2700 3890 2710
rect 4280 2700 4770 2710
rect 5180 2700 5220 2710
rect 5380 2700 5470 2710
rect 6170 2700 6510 2710
rect 6540 2700 7000 2710
rect 7660 2700 8120 2710
rect 9610 2700 9640 2710
rect 9980 2700 9990 2710
rect 0 2690 1070 2700
rect 1130 2690 1980 2700
rect 3150 2690 3890 2700
rect 3900 2690 3910 2700
rect 4280 2690 4860 2700
rect 5170 2690 5220 2700
rect 5380 2690 5460 2700
rect 6180 2690 6510 2700
rect 6540 2690 6980 2700
rect 7670 2690 8110 2700
rect 9630 2690 9660 2700
rect 9990 2690 9990 2700
rect 0 2680 1070 2690
rect 1130 2680 1980 2690
rect 3150 2680 3890 2690
rect 4280 2680 4840 2690
rect 5160 2680 5210 2690
rect 5380 2680 5450 2690
rect 6190 2680 6510 2690
rect 6540 2680 6960 2690
rect 7670 2680 8100 2690
rect 9650 2680 9680 2690
rect 0 2670 1060 2680
rect 1120 2670 1980 2680
rect 3150 2670 3890 2680
rect 4230 2670 4240 2680
rect 4270 2670 4840 2680
rect 5150 2670 5190 2680
rect 5370 2670 5440 2680
rect 6200 2670 6510 2680
rect 6540 2670 6950 2680
rect 7680 2670 8090 2680
rect 9670 2670 9700 2680
rect 0 2660 1060 2670
rect 1110 2660 1970 2670
rect 2950 2660 3020 2670
rect 3150 2660 3890 2670
rect 4220 2660 4240 2670
rect 4270 2660 4830 2670
rect 4900 2660 4910 2670
rect 5140 2660 5180 2670
rect 5370 2660 5430 2670
rect 6210 2660 6510 2670
rect 6540 2660 6940 2670
rect 7690 2660 8080 2670
rect 9690 2660 9720 2670
rect 0 2650 1050 2660
rect 1100 2650 1960 2660
rect 2220 2650 2330 2660
rect 2910 2650 3090 2660
rect 3150 2650 3890 2660
rect 4210 2650 4240 2660
rect 4270 2650 4820 2660
rect 4870 2650 4900 2660
rect 5120 2650 5160 2660
rect 5370 2650 5420 2660
rect 6220 2650 6510 2660
rect 6530 2650 6920 2660
rect 7690 2650 8070 2660
rect 9710 2650 9740 2660
rect 0 2640 1050 2650
rect 1100 2640 1960 2650
rect 2170 2640 2350 2650
rect 2880 2640 2950 2650
rect 3060 2640 3120 2650
rect 3150 2640 3890 2650
rect 4210 2640 4240 2650
rect 4270 2640 4810 2650
rect 4820 2640 4830 2650
rect 4840 2640 4880 2650
rect 5100 2640 5130 2650
rect 5360 2640 5410 2650
rect 6220 2640 6510 2650
rect 6530 2640 6910 2650
rect 7700 2640 8060 2650
rect 9080 2640 9190 2650
rect 9730 2640 9760 2650
rect 0 2630 1040 2640
rect 1090 2630 1960 2640
rect 2150 2630 2190 2640
rect 2280 2630 2370 2640
rect 2870 2630 2930 2640
rect 3080 2630 3900 2640
rect 4210 2630 4230 2640
rect 4270 2630 4730 2640
rect 4740 2630 4800 2640
rect 4810 2630 4860 2640
rect 5080 2630 5110 2640
rect 5360 2630 5400 2640
rect 6240 2630 6510 2640
rect 6530 2630 6900 2640
rect 7710 2630 8050 2640
rect 9080 2630 9180 2640
rect 9750 2630 9780 2640
rect 9850 2630 9990 2640
rect 0 2620 1040 2630
rect 1090 2620 1950 2630
rect 2120 2620 2160 2630
rect 2310 2620 2380 2630
rect 2860 2620 2910 2630
rect 3110 2620 3230 2630
rect 3240 2620 3900 2630
rect 4210 2620 4230 2630
rect 4270 2620 4830 2630
rect 5060 2620 5090 2630
rect 5350 2620 5380 2630
rect 6240 2620 6510 2630
rect 6520 2620 6890 2630
rect 7710 2620 8050 2630
rect 9080 2620 9170 2630
rect 9770 2620 9800 2630
rect 9860 2620 9990 2630
rect 0 2610 1030 2620
rect 1090 2610 1950 2620
rect 2100 2610 2130 2620
rect 2270 2610 2290 2620
rect 2340 2610 2390 2620
rect 2860 2610 2910 2620
rect 2940 2610 3040 2620
rect 3120 2610 3890 2620
rect 4210 2610 4230 2620
rect 4270 2610 4800 2620
rect 5040 2610 5080 2620
rect 5340 2610 5360 2620
rect 6250 2610 6510 2620
rect 6520 2610 6880 2620
rect 7720 2610 8030 2620
rect 9080 2610 9160 2620
rect 9790 2610 9820 2620
rect 9870 2610 9990 2620
rect 0 2600 1030 2610
rect 1080 2600 1940 2610
rect 2080 2600 2120 2610
rect 2190 2600 2320 2610
rect 2360 2600 2390 2610
rect 2860 2600 3110 2610
rect 3130 2600 3250 2610
rect 3260 2600 3890 2610
rect 4210 2600 4230 2610
rect 4270 2600 4780 2610
rect 5010 2600 5050 2610
rect 6250 2600 6510 2610
rect 6520 2600 6870 2610
rect 7730 2600 8030 2610
rect 9080 2600 9160 2610
rect 9800 2600 9840 2610
rect 9890 2600 9990 2610
rect 0 2590 1020 2600
rect 1080 2590 1940 2600
rect 2070 2590 2090 2600
rect 2160 2590 2390 2600
rect 2860 2590 3130 2600
rect 3160 2590 3900 2600
rect 4210 2590 4230 2600
rect 4260 2590 4740 2600
rect 4970 2590 5030 2600
rect 6260 2590 6510 2600
rect 6520 2590 6860 2600
rect 7740 2590 8020 2600
rect 9080 2590 9160 2600
rect 9830 2590 9870 2600
rect 9910 2590 9990 2600
rect 0 2580 1020 2590
rect 1060 2580 1940 2590
rect 2060 2580 2080 2590
rect 2130 2580 2390 2590
rect 2850 2580 3900 2590
rect 4260 2580 4690 2590
rect 4920 2580 5010 2590
rect 6270 2580 6510 2590
rect 6520 2580 6860 2590
rect 7740 2580 8000 2590
rect 9100 2580 9110 2590
rect 9840 2580 9890 2590
rect 9930 2580 9990 2590
rect 0 2570 1010 2580
rect 1060 2570 1930 2580
rect 2050 2570 2070 2580
rect 2120 2570 2400 2580
rect 2840 2570 2970 2580
rect 2980 2570 3270 2580
rect 3280 2570 3900 2580
rect 4250 2570 4540 2580
rect 4870 2570 4990 2580
rect 6270 2570 6850 2580
rect 7750 2570 7990 2580
rect 9500 2570 9520 2580
rect 9870 2570 9910 2580
rect 9950 2570 9990 2580
rect 0 2560 1010 2570
rect 1060 2560 1930 2570
rect 2040 2560 2330 2570
rect 2350 2560 2410 2570
rect 2840 2560 2890 2570
rect 2910 2560 3270 2570
rect 3280 2560 3910 2570
rect 4250 2560 4500 2570
rect 4800 2560 4950 2570
rect 4960 2560 4970 2570
rect 4980 2560 4990 2570
rect 6280 2560 6840 2570
rect 7760 2560 7980 2570
rect 9490 2560 9540 2570
rect 9880 2560 9930 2570
rect 9970 2560 9990 2570
rect 0 2550 1000 2560
rect 1060 2550 1930 2560
rect 2020 2550 2330 2560
rect 2360 2550 2410 2560
rect 2830 2550 2880 2560
rect 2910 2550 3960 2560
rect 3980 2550 3990 2560
rect 4180 2550 4230 2560
rect 4270 2550 4500 2560
rect 4690 2550 4730 2560
rect 4740 2550 4920 2560
rect 4930 2550 4940 2560
rect 6280 2550 6830 2560
rect 7770 2550 7970 2560
rect 9390 2550 9410 2560
rect 9440 2550 9470 2560
rect 9500 2550 9560 2560
rect 9900 2550 9950 2560
rect 0 2540 1000 2550
rect 1060 2540 1930 2550
rect 2030 2540 2330 2550
rect 2390 2540 2420 2550
rect 2830 2540 2870 2550
rect 2910 2540 3920 2550
rect 4170 2540 4230 2550
rect 4240 2540 4260 2550
rect 4300 2540 4510 2550
rect 4600 2540 4850 2550
rect 4870 2540 4880 2550
rect 6290 2540 6820 2550
rect 7780 2540 7960 2550
rect 9430 2540 9460 2550
rect 9520 2540 9580 2550
rect 9920 2540 9970 2550
rect 0 2530 990 2540
rect 1040 2530 1920 2540
rect 2020 2530 2330 2540
rect 2390 2530 2420 2540
rect 2840 2530 2860 2540
rect 2910 2530 2920 2540
rect 3150 2530 3920 2540
rect 4160 2530 4840 2540
rect 6300 2530 6810 2540
rect 7780 2530 7940 2540
rect 9350 2530 9370 2540
rect 9390 2530 9420 2540
rect 9440 2530 9480 2540
rect 9520 2530 9560 2540
rect 9580 2530 9590 2540
rect 9940 2530 9980 2540
rect 0 2520 990 2530
rect 1040 2520 1920 2530
rect 2010 2520 2330 2530
rect 3190 2520 3920 2530
rect 4160 2520 4720 2530
rect 6300 2520 6800 2530
rect 7790 2520 7930 2530
rect 9340 2520 9420 2530
rect 9430 2520 9480 2530
rect 9520 2520 9610 2530
rect 9960 2520 9990 2530
rect 0 2510 980 2520
rect 1050 2510 1920 2520
rect 3190 2510 3920 2520
rect 3940 2510 3950 2520
rect 3960 2510 3970 2520
rect 4160 2510 4670 2520
rect 4690 2510 4700 2520
rect 6310 2510 6790 2520
rect 7280 2510 7310 2520
rect 7790 2510 7920 2520
rect 9330 2510 9410 2520
rect 9440 2510 9470 2520
rect 9500 2510 9610 2520
rect 9620 2510 9640 2520
rect 9980 2510 9990 2520
rect 0 2500 980 2510
rect 1040 2500 1920 2510
rect 3200 2500 3930 2510
rect 3960 2500 3970 2510
rect 4120 2500 4150 2510
rect 4160 2500 4650 2510
rect 4800 2500 4830 2510
rect 6310 2500 6790 2510
rect 7290 2500 7310 2510
rect 7800 2500 7900 2510
rect 9290 2500 9410 2510
rect 9440 2500 9470 2510
rect 9480 2500 9570 2510
rect 9610 2500 9670 2510
rect 0 2490 970 2500
rect 1040 2490 1910 2500
rect 3210 2490 3940 2500
rect 3960 2490 3980 2500
rect 4130 2490 4650 2500
rect 6320 2490 6780 2500
rect 7300 2490 7320 2500
rect 7800 2490 7880 2500
rect 9270 2490 9560 2500
rect 9610 2490 9680 2500
rect 0 2480 970 2490
rect 1040 2480 1910 2490
rect 3210 2480 3980 2490
rect 4130 2480 4600 2490
rect 4610 2480 4650 2490
rect 6320 2480 6770 2490
rect 7300 2480 7330 2490
rect 7810 2480 7860 2490
rect 9260 2480 9700 2490
rect 0 2470 960 2480
rect 1040 2470 1910 2480
rect 3220 2470 3910 2480
rect 3920 2470 3940 2480
rect 3950 2470 3990 2480
rect 4080 2470 4100 2480
rect 4110 2470 4590 2480
rect 4630 2470 4650 2480
rect 6330 2470 6770 2480
rect 7310 2470 7340 2480
rect 7820 2470 7840 2480
rect 9250 2470 9450 2480
rect 9460 2470 9720 2480
rect 0 2460 960 2470
rect 1030 2460 1910 2470
rect 3230 2460 3910 2470
rect 3920 2460 3940 2470
rect 3950 2460 3980 2470
rect 3990 2460 4020 2470
rect 4080 2460 4590 2470
rect 6330 2460 6760 2470
rect 7310 2460 7340 2470
rect 9240 2460 9450 2470
rect 9490 2460 9500 2470
rect 9510 2460 9730 2470
rect 0 2450 950 2460
rect 1030 2450 1900 2460
rect 3240 2450 3910 2460
rect 3920 2450 3950 2460
rect 3960 2450 3980 2460
rect 4010 2450 4020 2460
rect 4090 2450 4580 2460
rect 6340 2450 6760 2460
rect 7290 2450 7350 2460
rect 9230 2450 9290 2460
rect 9300 2450 9460 2460
rect 9500 2450 9730 2460
rect 0 2440 950 2450
rect 1040 2440 1900 2450
rect 3250 2440 3950 2450
rect 3960 2440 3980 2450
rect 4040 2440 4060 2450
rect 4080 2440 4560 2450
rect 4570 2440 4600 2450
rect 4610 2440 4620 2450
rect 6350 2440 6750 2450
rect 7290 2440 7360 2450
rect 9230 2440 9270 2450
rect 9300 2440 9430 2450
rect 9450 2440 9470 2450
rect 9520 2440 9680 2450
rect 9700 2440 9730 2450
rect 0 2430 940 2440
rect 1040 2430 1900 2440
rect 3250 2430 3920 2440
rect 3930 2430 3980 2440
rect 4040 2430 4580 2440
rect 4590 2430 4610 2440
rect 4890 2430 4900 2440
rect 6350 2430 6750 2440
rect 7310 2430 7370 2440
rect 9230 2430 9260 2440
rect 9300 2430 9430 2440
rect 9450 2430 9480 2440
rect 9520 2430 9670 2440
rect 9710 2430 9790 2440
rect 0 2420 940 2430
rect 1030 2420 1900 2430
rect 3260 2420 3980 2430
rect 4000 2420 4010 2430
rect 4040 2420 4570 2430
rect 4590 2420 4600 2430
rect 6360 2420 6750 2430
rect 7330 2420 7380 2430
rect 9240 2420 9270 2430
rect 9300 2420 9380 2430
rect 9400 2420 9470 2430
rect 9530 2420 9540 2430
rect 9560 2420 9650 2430
rect 9710 2420 9790 2430
rect 0 2410 930 2420
rect 1030 2410 1900 2420
rect 3270 2410 4580 2420
rect 4680 2410 4690 2420
rect 4820 2410 4840 2420
rect 6360 2410 6740 2420
rect 7350 2410 7390 2420
rect 9160 2410 9170 2420
rect 9310 2410 9330 2420
rect 9400 2410 9430 2420
rect 9440 2410 9460 2420
rect 9470 2410 9480 2420
rect 9570 2410 9640 2420
rect 9710 2410 9800 2420
rect 0 2400 930 2410
rect 1020 2400 1900 2410
rect 3280 2400 4530 2410
rect 4560 2400 4590 2410
rect 4650 2400 4660 2410
rect 4670 2400 4700 2410
rect 4790 2400 4800 2410
rect 6370 2400 6740 2410
rect 7360 2400 7400 2410
rect 9160 2400 9170 2410
rect 9300 2400 9320 2410
rect 9400 2400 9420 2410
rect 9440 2400 9480 2410
rect 9600 2400 9650 2410
rect 9680 2400 9810 2410
rect 0 2390 920 2400
rect 1020 2390 1890 2400
rect 3290 2390 4560 2400
rect 4570 2390 4600 2400
rect 4680 2390 4700 2400
rect 4710 2390 4720 2400
rect 6370 2390 6740 2400
rect 7380 2390 7410 2400
rect 9160 2390 9180 2400
rect 9290 2390 9320 2400
rect 9430 2390 9470 2400
rect 9600 2390 9650 2400
rect 9680 2390 9840 2400
rect 0 2380 920 2390
rect 1010 2380 1890 2390
rect 3290 2380 4590 2390
rect 6380 2380 6740 2390
rect 7400 2380 7430 2390
rect 9160 2380 9200 2390
rect 9280 2380 9310 2390
rect 9400 2380 9460 2390
rect 9590 2380 9610 2390
rect 9630 2380 9690 2390
rect 9720 2380 9820 2390
rect 0 2370 910 2380
rect 1010 2370 1880 2380
rect 3290 2370 4540 2380
rect 4710 2370 4720 2380
rect 6380 2370 6730 2380
rect 7410 2370 7440 2380
rect 8390 2370 8400 2380
rect 9160 2370 9200 2380
rect 9260 2370 9320 2380
rect 9380 2370 9410 2380
rect 9420 2370 9450 2380
rect 9600 2370 9620 2380
rect 9630 2370 9680 2380
rect 9710 2370 9800 2380
rect 9810 2370 9820 2380
rect 0 2360 910 2370
rect 1010 2360 1880 2370
rect 3290 2360 4480 2370
rect 4580 2360 4690 2370
rect 6390 2360 6730 2370
rect 7430 2360 7440 2370
rect 8390 2360 8400 2370
rect 9160 2360 9210 2370
rect 9260 2360 9270 2370
rect 9300 2360 9320 2370
rect 9390 2360 9400 2370
rect 9420 2360 9460 2370
rect 9680 2360 9800 2370
rect 9810 2360 9830 2370
rect 0 2350 900 2360
rect 1000 2350 1880 2360
rect 3300 2350 4590 2360
rect 4600 2350 4610 2360
rect 4640 2350 4650 2360
rect 6390 2350 6730 2360
rect 8390 2350 8400 2360
rect 9160 2350 9210 2360
rect 9330 2350 9350 2360
rect 9390 2350 9460 2360
rect 9670 2350 9800 2360
rect 9810 2350 9840 2360
rect 0 2340 900 2350
rect 1000 2340 1880 2350
rect 3300 2340 4500 2350
rect 6400 2340 6730 2350
rect 7460 2340 7470 2350
rect 8390 2340 8420 2350
rect 9160 2340 9210 2350
rect 9360 2340 9430 2350
rect 9550 2340 9620 2350
rect 9660 2340 9710 2350
rect 9730 2340 9770 2350
rect 9810 2340 9830 2350
rect 0 2330 890 2340
rect 1000 2330 1870 2340
rect 3310 2330 4510 2340
rect 4520 2330 4530 2340
rect 6400 2330 6730 2340
rect 8390 2330 8400 2340
rect 8410 2330 8440 2340
rect 9160 2330 9210 2340
rect 9260 2330 9270 2340
rect 9300 2330 9330 2340
rect 9450 2330 9490 2340
rect 9560 2330 9710 2340
rect 9730 2330 9770 2340
rect 0 2320 880 2330
rect 990 2320 1870 2330
rect 3310 2320 4510 2330
rect 6410 2320 6730 2330
rect 7480 2320 7500 2330
rect 8380 2320 8410 2330
rect 8420 2320 8490 2330
rect 9150 2320 9210 2330
rect 9250 2320 9360 2330
rect 9450 2320 9490 2330
rect 9540 2320 9550 2330
rect 9560 2320 9710 2330
rect 9730 2320 9790 2330
rect 9800 2320 9810 2330
rect 0 2310 880 2320
rect 990 2310 1870 2320
rect 3310 2310 4500 2320
rect 6420 2310 6730 2320
rect 7490 2310 7510 2320
rect 8370 2310 8520 2320
rect 9160 2310 9210 2320
rect 9230 2310 9360 2320
rect 9390 2310 9410 2320
rect 9440 2310 9470 2320
rect 9490 2310 9820 2320
rect 0 2300 870 2310
rect 990 2300 1870 2310
rect 3310 2300 4470 2310
rect 6420 2300 6730 2310
rect 7500 2300 7530 2310
rect 8360 2300 8540 2310
rect 9150 2300 9210 2310
rect 9230 2300 9360 2310
rect 9380 2300 9420 2310
rect 9440 2300 9470 2310
rect 9500 2300 9620 2310
rect 9640 2300 9830 2310
rect 0 2290 870 2300
rect 990 2290 1860 2300
rect 3320 2290 4440 2300
rect 6430 2290 6730 2300
rect 7500 2290 7540 2300
rect 8360 2290 8550 2300
rect 9160 2290 9200 2300
rect 9220 2290 9250 2300
rect 9260 2290 9480 2300
rect 9590 2290 9610 2300
rect 9640 2290 9720 2300
rect 9740 2290 9820 2300
rect 0 2280 860 2290
rect 980 2280 1860 2290
rect 3320 2280 4070 2290
rect 4180 2280 4330 2290
rect 6430 2280 6730 2290
rect 7510 2280 7560 2290
rect 8360 2280 8560 2290
rect 9150 2280 9190 2290
rect 9210 2280 9250 2290
rect 9260 2280 9490 2290
rect 9590 2280 9730 2290
rect 9740 2280 9790 2290
rect 0 2270 860 2280
rect 980 2270 1860 2280
rect 3320 2270 4070 2280
rect 6440 2270 6730 2280
rect 7510 2270 7570 2280
rect 8360 2270 8570 2280
rect 9150 2270 9180 2280
rect 9190 2270 9260 2280
rect 9270 2270 9350 2280
rect 9370 2270 9500 2280
rect 9560 2270 9790 2280
rect 0 2260 850 2270
rect 980 2260 1850 2270
rect 3320 2260 4130 2270
rect 6440 2260 6730 2270
rect 6890 2260 6900 2270
rect 7090 2260 7120 2270
rect 7520 2260 7580 2270
rect 8360 2260 8580 2270
rect 9150 2260 9340 2270
rect 9370 2260 9520 2270
rect 9530 2260 9540 2270
rect 9550 2260 9790 2270
rect 0 2250 850 2260
rect 980 2250 1850 2260
rect 3320 2250 4260 2260
rect 4270 2250 4290 2260
rect 4310 2250 4330 2260
rect 6450 2250 6740 2260
rect 6900 2250 6910 2260
rect 6920 2250 6940 2260
rect 7110 2250 7150 2260
rect 7170 2250 7180 2260
rect 7520 2250 7590 2260
rect 8360 2250 8600 2260
rect 9140 2250 9590 2260
rect 9600 2250 9800 2260
rect 0 2240 840 2250
rect 980 2240 1850 2250
rect 3330 2240 4340 2250
rect 6450 2240 6740 2250
rect 6940 2240 6950 2250
rect 7130 2240 7220 2250
rect 7520 2240 7600 2250
rect 8360 2240 8630 2250
rect 9110 2240 9250 2250
rect 9270 2240 9590 2250
rect 9600 2240 9800 2250
rect 0 2230 840 2240
rect 980 2230 1850 2240
rect 3330 2230 4350 2240
rect 6460 2230 6740 2240
rect 6930 2230 6980 2240
rect 6990 2230 7000 2240
rect 7140 2230 7240 2240
rect 7520 2230 7610 2240
rect 8360 2230 8660 2240
rect 8740 2230 8760 2240
rect 9090 2230 9250 2240
rect 9290 2230 9580 2240
rect 9590 2230 9800 2240
rect 0 2220 830 2230
rect 980 2220 1850 2230
rect 3340 2220 4360 2230
rect 6460 2220 6740 2230
rect 6960 2220 7040 2230
rect 7090 2220 7100 2230
rect 7140 2220 7260 2230
rect 7530 2220 7620 2230
rect 8360 2220 8690 2230
rect 8710 2220 8820 2230
rect 9060 2220 9250 2230
rect 9310 2220 9550 2230
rect 9590 2220 9810 2230
rect 0 2210 830 2220
rect 980 2210 1850 2220
rect 3340 2210 4340 2220
rect 6470 2210 6740 2220
rect 6970 2210 7290 2220
rect 7530 2210 7630 2220
rect 8360 2210 8830 2220
rect 9010 2210 9250 2220
rect 9340 2210 9550 2220
rect 9600 2210 9810 2220
rect 0 2200 820 2210
rect 980 2200 1850 2210
rect 3340 2200 4350 2210
rect 6470 2200 6740 2210
rect 6990 2200 7300 2210
rect 7530 2200 7640 2210
rect 8360 2200 8850 2210
rect 8940 2200 9250 2210
rect 9360 2200 9580 2210
rect 9590 2200 9670 2210
rect 9720 2200 9810 2210
rect 0 2190 820 2200
rect 980 2190 1850 2200
rect 3340 2190 4360 2200
rect 6470 2190 6740 2200
rect 7010 2190 7320 2200
rect 7530 2190 7650 2200
rect 8360 2190 9250 2200
rect 9380 2190 9680 2200
rect 9730 2190 9810 2200
rect 0 2180 810 2190
rect 980 2180 1840 2190
rect 2680 2180 2750 2190
rect 3340 2180 4350 2190
rect 6480 2180 6740 2190
rect 7030 2180 7330 2190
rect 7350 2180 7380 2190
rect 7520 2180 7650 2190
rect 8360 2180 9250 2190
rect 9400 2180 9720 2190
rect 9740 2180 9820 2190
rect 9970 2180 9980 2190
rect 0 2170 800 2180
rect 980 2170 1840 2180
rect 2450 2170 2510 2180
rect 2660 2170 2750 2180
rect 3330 2170 4360 2180
rect 6480 2170 6750 2180
rect 7050 2170 7380 2180
rect 7520 2170 7670 2180
rect 8370 2170 9240 2180
rect 9420 2170 9810 2180
rect 0 2160 800 2170
rect 980 2160 1840 2170
rect 2440 2160 2530 2170
rect 2650 2160 2740 2170
rect 3330 2160 4360 2170
rect 6490 2160 6750 2170
rect 7060 2160 7310 2170
rect 7320 2160 7380 2170
rect 7510 2160 7670 2170
rect 8370 2160 9240 2170
rect 9430 2160 9560 2170
rect 9570 2160 9790 2170
rect 0 2150 790 2160
rect 980 2150 1840 2160
rect 2440 2150 2540 2160
rect 2640 2150 2730 2160
rect 3330 2150 4360 2160
rect 6490 2150 6750 2160
rect 7080 2150 7290 2160
rect 7320 2150 7390 2160
rect 7520 2150 7670 2160
rect 8370 2150 9270 2160
rect 9460 2150 9560 2160
rect 9600 2150 9790 2160
rect 0 2140 790 2150
rect 970 2140 1840 2150
rect 2450 2140 2540 2150
rect 2640 2140 2710 2150
rect 3340 2140 4360 2150
rect 6500 2140 6750 2150
rect 7090 2140 7250 2150
rect 7320 2140 7400 2150
rect 7510 2140 7670 2150
rect 7680 2140 7700 2150
rect 8380 2140 9290 2150
rect 9470 2140 9560 2150
rect 9600 2140 9780 2150
rect 0 2130 780 2140
rect 970 2130 1840 2140
rect 2460 2130 2530 2140
rect 3340 2130 4360 2140
rect 6510 2130 6750 2140
rect 7070 2130 7240 2140
rect 7320 2130 7400 2140
rect 7510 2130 7710 2140
rect 8380 2130 9230 2140
rect 9250 2130 9310 2140
rect 9490 2130 9570 2140
rect 9590 2130 9670 2140
rect 9690 2130 9780 2140
rect 0 2120 780 2130
rect 970 2120 1840 2130
rect 3340 2120 4370 2130
rect 6510 2120 6750 2130
rect 7090 2120 7220 2130
rect 7320 2120 7410 2130
rect 7490 2120 7730 2130
rect 8390 2120 9230 2130
rect 9250 2120 9330 2130
rect 9510 2120 9570 2130
rect 9590 2120 9670 2130
rect 9710 2120 9770 2130
rect 0 2110 770 2120
rect 970 2110 1840 2120
rect 3340 2110 4360 2120
rect 6510 2110 6760 2120
rect 7320 2110 7420 2120
rect 7480 2110 7750 2120
rect 8400 2110 9340 2120
rect 9530 2110 9560 2120
rect 9720 2110 9740 2120
rect 0 2100 770 2110
rect 970 2100 1840 2110
rect 3340 2100 4350 2110
rect 6520 2100 6760 2110
rect 7320 2100 7830 2110
rect 8410 2100 9360 2110
rect 9630 2100 9700 2110
rect 0 2090 760 2100
rect 960 2090 1840 2100
rect 3340 2090 4340 2100
rect 6530 2090 6760 2100
rect 7240 2090 7250 2100
rect 7320 2090 7830 2100
rect 8420 2090 9250 2100
rect 9260 2090 9360 2100
rect 9560 2090 9710 2100
rect 0 2080 760 2090
rect 950 2080 1840 2090
rect 3340 2080 4340 2090
rect 6530 2080 6760 2090
rect 7320 2080 7830 2090
rect 8430 2080 9230 2090
rect 9270 2080 9330 2090
rect 9480 2080 9690 2090
rect 0 2070 750 2080
rect 950 2070 1840 2080
rect 3340 2070 4350 2080
rect 6530 2070 6760 2080
rect 7180 2070 7210 2080
rect 7320 2070 7830 2080
rect 8460 2070 9220 2080
rect 9400 2070 9670 2080
rect 0 2060 750 2070
rect 950 2060 1840 2070
rect 3350 2060 4350 2070
rect 6540 2060 6760 2070
rect 7330 2060 7730 2070
rect 7760 2060 7830 2070
rect 8480 2060 9170 2070
rect 9320 2060 9560 2070
rect 9590 2060 9640 2070
rect 0 2050 740 2060
rect 950 2050 1840 2060
rect 3350 2050 4370 2060
rect 6540 2050 6770 2060
rect 7330 2050 7730 2060
rect 7740 2050 7750 2060
rect 7760 2050 7830 2060
rect 8510 2050 9150 2060
rect 9250 2050 9490 2060
rect 0 2040 740 2050
rect 950 2040 1840 2050
rect 3350 2040 4370 2050
rect 6540 2040 6770 2050
rect 7330 2040 7730 2050
rect 7780 2040 7850 2050
rect 8530 2040 9140 2050
rect 9170 2040 9470 2050
rect 0 2030 730 2040
rect 960 2030 1840 2040
rect 3350 2030 4370 2040
rect 6540 2030 6770 2040
rect 7330 2030 7730 2040
rect 7790 2030 7850 2040
rect 8550 2030 9110 2040
rect 9150 2030 9320 2040
rect 9390 2030 9460 2040
rect 0 2020 730 2030
rect 950 2020 1840 2030
rect 3350 2020 4350 2030
rect 4360 2020 4370 2030
rect 6540 2020 6770 2030
rect 7330 2020 7740 2030
rect 7790 2020 7860 2030
rect 7870 2020 7890 2030
rect 8570 2020 9090 2030
rect 9150 2020 9220 2030
rect 9400 2020 9410 2030
rect 9420 2020 9460 2030
rect 0 2010 720 2020
rect 940 2010 1840 2020
rect 3350 2010 4370 2020
rect 6540 2010 6770 2020
rect 7330 2010 7760 2020
rect 7790 2010 7850 2020
rect 7860 2010 7940 2020
rect 8600 2010 9080 2020
rect 0 2000 720 2010
rect 930 2000 1840 2010
rect 3350 2000 4340 2010
rect 4350 2000 4360 2010
rect 6540 2000 6770 2010
rect 7330 2000 7850 2010
rect 7890 2000 7950 2010
rect 8620 2000 9070 2010
rect 0 1990 710 2000
rect 930 1990 1840 2000
rect 3350 1990 4340 2000
rect 6540 1990 6770 2000
rect 7330 1990 7720 2000
rect 7760 1990 7820 2000
rect 7830 1990 7860 2000
rect 8680 1990 9060 2000
rect 0 1980 710 1990
rect 930 1980 1840 1990
rect 3350 1980 4330 1990
rect 6550 1980 6770 1990
rect 7330 1980 7720 1990
rect 7850 1980 7870 1990
rect 8710 1980 9060 1990
rect 0 1970 700 1980
rect 930 1970 1840 1980
rect 3350 1970 4350 1980
rect 6550 1970 6780 1980
rect 7330 1970 7720 1980
rect 7860 1970 7880 1980
rect 8730 1970 9040 1980
rect 0 1960 700 1970
rect 940 1960 1840 1970
rect 3350 1960 4360 1970
rect 6550 1960 6780 1970
rect 7330 1960 7730 1970
rect 7870 1960 7890 1970
rect 8770 1960 8810 1970
rect 8950 1960 9010 1970
rect 0 1950 690 1960
rect 940 1950 1840 1960
rect 3350 1950 4360 1960
rect 6550 1950 6780 1960
rect 7330 1950 7730 1960
rect 7880 1950 7950 1960
rect 9890 1950 9900 1960
rect 0 1940 690 1950
rect 930 1940 1840 1950
rect 3350 1940 4360 1950
rect 6560 1940 6780 1950
rect 7340 1940 7730 1950
rect 9890 1940 9900 1950
rect 0 1930 680 1940
rect 930 1930 1840 1940
rect 3350 1930 4380 1940
rect 6560 1930 6780 1940
rect 7340 1930 7730 1940
rect 9660 1930 9680 1940
rect 9880 1930 9900 1940
rect 0 1920 680 1930
rect 920 1920 1840 1930
rect 3350 1920 4380 1930
rect 6570 1920 6780 1930
rect 7340 1920 7730 1930
rect 9880 1920 9910 1930
rect 0 1910 670 1920
rect 920 1910 1840 1920
rect 3350 1910 4410 1920
rect 4590 1910 4610 1920
rect 6570 1910 6780 1920
rect 7340 1910 7730 1920
rect 9890 1910 9900 1920
rect 9960 1910 9970 1920
rect 0 1900 670 1910
rect 920 1900 1840 1910
rect 3350 1900 4390 1910
rect 4420 1900 4430 1910
rect 4520 1900 4540 1910
rect 6580 1900 6780 1910
rect 7340 1900 7730 1910
rect 9690 1900 9720 1910
rect 9960 1900 9970 1910
rect 0 1890 660 1900
rect 920 1890 1840 1900
rect 3350 1890 4350 1900
rect 4380 1890 4400 1900
rect 4540 1890 4550 1900
rect 4560 1890 4570 1900
rect 6590 1890 6780 1900
rect 7340 1890 7740 1900
rect 9680 1890 9740 1900
rect 0 1880 660 1890
rect 910 1880 1840 1890
rect 3350 1880 4330 1890
rect 4370 1880 4400 1890
rect 6570 1880 6790 1890
rect 7340 1880 7740 1890
rect 9690 1880 9760 1890
rect 0 1870 650 1880
rect 920 1870 1840 1880
rect 2600 1870 2620 1880
rect 3340 1870 4310 1880
rect 4360 1870 4390 1880
rect 4570 1870 4590 1880
rect 4600 1870 4610 1880
rect 6580 1870 6790 1880
rect 7340 1870 7740 1880
rect 9160 1870 9190 1880
rect 9690 1870 9770 1880
rect 0 1860 650 1870
rect 920 1860 1850 1870
rect 3340 1860 4280 1870
rect 4340 1860 4380 1870
rect 4420 1860 4430 1870
rect 4500 1860 4510 1870
rect 4550 1860 4580 1870
rect 6590 1860 6790 1870
rect 7340 1860 7740 1870
rect 9120 1860 9190 1870
rect 9690 1860 9770 1870
rect 9990 1860 9990 1870
rect 0 1850 640 1860
rect 910 1850 1840 1860
rect 2780 1850 2790 1860
rect 3340 1850 4280 1860
rect 4320 1850 4350 1860
rect 4400 1850 4430 1860
rect 4500 1850 4510 1860
rect 5140 1850 5150 1860
rect 6600 1850 6790 1860
rect 7340 1850 7740 1860
rect 9120 1850 9190 1860
rect 9310 1850 9330 1860
rect 9690 1850 9730 1860
rect 9750 1850 9760 1860
rect 9980 1850 9990 1860
rect 0 1840 640 1850
rect 910 1840 1850 1850
rect 2760 1840 2820 1850
rect 3340 1840 4340 1850
rect 4370 1840 4420 1850
rect 4500 1840 4510 1850
rect 5080 1840 5140 1850
rect 6610 1840 6790 1850
rect 7340 1840 7740 1850
rect 9120 1840 9180 1850
rect 9320 1840 9330 1850
rect 9700 1840 9760 1850
rect 9980 1840 9990 1850
rect 0 1830 630 1840
rect 910 1830 1850 1840
rect 2710 1830 2850 1840
rect 3340 1830 4270 1840
rect 4290 1830 4330 1840
rect 4350 1830 4430 1840
rect 4500 1830 4510 1840
rect 5080 1830 5100 1840
rect 6560 1830 6590 1840
rect 6620 1830 6790 1840
rect 7340 1830 7750 1840
rect 9120 1830 9180 1840
rect 9210 1830 9220 1840
rect 9310 1830 9320 1840
rect 9400 1830 9410 1840
rect 9700 1830 9760 1840
rect 9970 1830 9990 1840
rect 0 1820 630 1830
rect 910 1820 1850 1830
rect 2430 1820 2440 1830
rect 2500 1820 2540 1830
rect 2560 1820 2860 1830
rect 3330 1820 4270 1830
rect 4290 1820 4330 1830
rect 4340 1820 4420 1830
rect 4500 1820 4510 1830
rect 5080 1820 5090 1830
rect 6570 1820 6610 1830
rect 6630 1820 6790 1830
rect 7350 1820 7740 1830
rect 9110 1820 9190 1830
rect 9390 1820 9420 1830
rect 9700 1820 9760 1830
rect 9960 1820 9980 1830
rect 0 1810 630 1820
rect 900 1810 1850 1820
rect 2360 1810 2410 1820
rect 2430 1810 2820 1820
rect 3330 1810 4270 1820
rect 4290 1810 4330 1820
rect 4350 1810 4420 1820
rect 4500 1810 4510 1820
rect 4600 1810 4610 1820
rect 5080 1810 5090 1820
rect 6560 1810 6790 1820
rect 7350 1810 7750 1820
rect 9110 1810 9200 1820
rect 9280 1810 9290 1820
rect 9390 1810 9430 1820
rect 9700 1810 9760 1820
rect 9960 1810 9980 1820
rect 0 1800 620 1810
rect 900 1800 1850 1810
rect 2330 1800 2460 1810
rect 2500 1800 2790 1810
rect 3330 1800 4270 1810
rect 4300 1800 4330 1810
rect 4340 1800 4420 1810
rect 4440 1800 4450 1810
rect 4500 1800 4510 1810
rect 4540 1800 4550 1810
rect 5240 1800 5250 1810
rect 6580 1800 6790 1810
rect 7350 1800 7750 1810
rect 9110 1800 9200 1810
rect 9410 1800 9450 1810
rect 9700 1800 9770 1810
rect 9960 1800 9970 1810
rect 0 1790 620 1800
rect 900 1790 1850 1800
rect 2330 1790 2390 1800
rect 2550 1790 2570 1800
rect 3320 1790 4110 1800
rect 4180 1790 4280 1800
rect 4300 1790 4330 1800
rect 4340 1790 4360 1800
rect 4400 1790 4420 1800
rect 4430 1790 4440 1800
rect 4500 1790 4510 1800
rect 4540 1790 4550 1800
rect 4640 1790 4650 1800
rect 5230 1790 5250 1800
rect 6590 1790 6790 1800
rect 7350 1790 7750 1800
rect 9110 1790 9220 1800
rect 9430 1790 9450 1800
rect 9700 1790 9760 1800
rect 9950 1790 9970 1800
rect 0 1780 610 1790
rect 890 1780 1850 1790
rect 3320 1780 4100 1790
rect 4200 1780 4280 1790
rect 4300 1780 4330 1790
rect 4410 1780 4420 1790
rect 4500 1780 4510 1790
rect 4630 1780 4650 1790
rect 4800 1780 4810 1790
rect 5230 1780 5240 1790
rect 6600 1780 6790 1790
rect 7350 1780 7750 1790
rect 9110 1780 9240 1790
rect 9700 1780 9740 1790
rect 9920 1780 9930 1790
rect 9940 1780 9960 1790
rect 0 1770 610 1780
rect 900 1770 1860 1780
rect 3320 1770 4090 1780
rect 4210 1770 4280 1780
rect 4300 1770 4330 1780
rect 4370 1770 4380 1780
rect 4410 1770 4430 1780
rect 4500 1770 4510 1780
rect 4630 1770 4650 1780
rect 4800 1770 4810 1780
rect 6620 1770 6800 1780
rect 7350 1770 7760 1780
rect 9110 1770 9220 1780
rect 9700 1770 9740 1780
rect 9920 1770 9930 1780
rect 9940 1770 9960 1780
rect 0 1760 610 1770
rect 890 1760 1860 1770
rect 3320 1760 4080 1770
rect 4220 1760 4280 1770
rect 4300 1760 4340 1770
rect 4360 1760 4390 1770
rect 4410 1760 4420 1770
rect 4450 1760 4460 1770
rect 5210 1760 5230 1770
rect 6620 1760 6800 1770
rect 7350 1760 7760 1770
rect 9110 1760 9210 1770
rect 9710 1760 9740 1770
rect 9930 1760 9950 1770
rect 0 1750 600 1760
rect 890 1750 1870 1760
rect 3310 1750 4070 1760
rect 4220 1750 4280 1760
rect 4300 1750 4380 1760
rect 4410 1750 4430 1760
rect 4450 1750 4460 1760
rect 4500 1750 4510 1760
rect 5210 1750 5220 1760
rect 5330 1750 5340 1760
rect 6620 1750 6800 1760
rect 7350 1750 7760 1760
rect 9110 1750 9200 1760
rect 9710 1750 9740 1760
rect 9760 1750 9780 1760
rect 9930 1750 9960 1760
rect 0 1740 600 1750
rect 890 1740 1870 1750
rect 3310 1740 4070 1750
rect 4230 1740 4280 1750
rect 4300 1740 4360 1750
rect 4410 1740 4430 1750
rect 5200 1740 5220 1750
rect 5330 1740 5340 1750
rect 6640 1740 6800 1750
rect 7350 1740 7770 1750
rect 9120 1740 9200 1750
rect 9710 1740 9740 1750
rect 9760 1740 9780 1750
rect 9930 1740 9940 1750
rect 0 1730 590 1740
rect 880 1730 1870 1740
rect 3310 1730 4070 1740
rect 4230 1730 4280 1740
rect 4310 1730 4350 1740
rect 4390 1730 4430 1740
rect 5200 1730 5210 1740
rect 5320 1730 5330 1740
rect 6660 1730 6800 1740
rect 7350 1730 7770 1740
rect 9120 1730 9200 1740
rect 9710 1730 9740 1740
rect 9760 1730 9780 1740
rect 9920 1730 9930 1740
rect 0 1720 590 1730
rect 880 1720 1880 1730
rect 3300 1720 4070 1730
rect 4230 1720 4280 1730
rect 4310 1720 4350 1730
rect 4360 1720 4430 1730
rect 4500 1720 4510 1730
rect 5190 1720 5210 1730
rect 5320 1720 5330 1730
rect 6670 1720 6800 1730
rect 7350 1720 7770 1730
rect 9120 1720 9190 1730
rect 9710 1720 9740 1730
rect 9760 1720 9780 1730
rect 9840 1720 9860 1730
rect 9910 1720 9920 1730
rect 0 1710 590 1720
rect 880 1710 1880 1720
rect 3300 1710 3480 1720
rect 3490 1710 4070 1720
rect 4240 1710 4290 1720
rect 4310 1710 4430 1720
rect 5190 1710 5200 1720
rect 5310 1710 5320 1720
rect 6200 1710 6230 1720
rect 6670 1710 6800 1720
rect 7360 1710 7760 1720
rect 9120 1710 9200 1720
rect 9710 1710 9740 1720
rect 9750 1710 9790 1720
rect 9840 1710 9860 1720
rect 9910 1710 9920 1720
rect 0 1700 580 1710
rect 870 1700 1880 1710
rect 3290 1700 4070 1710
rect 4240 1700 4290 1710
rect 4310 1700 4400 1710
rect 4780 1700 4810 1710
rect 5040 1700 5050 1710
rect 5180 1700 5190 1710
rect 6210 1700 6230 1710
rect 6670 1700 6800 1710
rect 7360 1700 7760 1710
rect 9120 1700 9200 1710
rect 9710 1700 9740 1710
rect 9760 1700 9780 1710
rect 9900 1700 9910 1710
rect 0 1690 580 1700
rect 870 1690 1880 1700
rect 3290 1690 4070 1700
rect 4250 1690 4290 1700
rect 4310 1690 4340 1700
rect 4350 1690 4400 1700
rect 4500 1690 4510 1700
rect 4780 1690 4790 1700
rect 5030 1690 5050 1700
rect 5180 1690 5190 1700
rect 5300 1690 5310 1700
rect 6210 1690 6240 1700
rect 6660 1690 6800 1700
rect 7360 1690 7770 1700
rect 9120 1690 9200 1700
rect 9710 1690 9740 1700
rect 9760 1690 9780 1700
rect 9900 1690 9910 1700
rect 0 1680 570 1690
rect 870 1680 1880 1690
rect 3280 1680 4070 1690
rect 4250 1680 4290 1690
rect 4310 1680 4340 1690
rect 4350 1680 4390 1690
rect 4500 1680 4510 1690
rect 5030 1680 5040 1690
rect 5170 1680 5180 1690
rect 5300 1680 5310 1690
rect 5450 1680 5460 1690
rect 6200 1680 6250 1690
rect 6660 1680 6800 1690
rect 7360 1680 7770 1690
rect 9120 1680 9200 1690
rect 9710 1680 9740 1690
rect 9760 1680 9780 1690
rect 9890 1680 9910 1690
rect 0 1670 570 1680
rect 870 1670 1890 1680
rect 3280 1670 4070 1680
rect 4260 1670 4290 1680
rect 4310 1670 4340 1680
rect 4360 1670 4380 1680
rect 4500 1670 4510 1680
rect 4530 1670 4560 1680
rect 5030 1670 5040 1680
rect 5160 1670 5180 1680
rect 5290 1670 5300 1680
rect 5440 1670 5450 1680
rect 6200 1670 6250 1680
rect 6650 1670 6800 1680
rect 7360 1670 7770 1680
rect 9120 1670 9200 1680
rect 9710 1670 9750 1680
rect 9770 1670 9790 1680
rect 9880 1670 9910 1680
rect 0 1660 570 1670
rect 870 1660 1890 1670
rect 3270 1660 4080 1670
rect 4260 1660 4290 1670
rect 4310 1660 4350 1670
rect 4500 1660 4550 1670
rect 5160 1660 5180 1670
rect 6200 1660 6260 1670
rect 6650 1660 6800 1670
rect 7360 1660 7770 1670
rect 9120 1660 9200 1670
rect 9720 1660 9740 1670
rect 9880 1660 9890 1670
rect 0 1650 560 1660
rect 870 1650 1890 1660
rect 3260 1650 4080 1660
rect 4270 1650 4290 1660
rect 4320 1650 4350 1660
rect 4400 1650 4430 1660
rect 4460 1650 4470 1660
rect 4540 1650 4550 1660
rect 4640 1650 4650 1660
rect 4710 1650 4730 1660
rect 4760 1650 4770 1660
rect 5160 1650 5170 1660
rect 5280 1650 5290 1660
rect 5420 1650 5430 1660
rect 6200 1650 6260 1660
rect 6650 1650 6800 1660
rect 7360 1650 7770 1660
rect 9120 1650 9200 1660
rect 0 1640 560 1650
rect 870 1640 1900 1650
rect 3260 1640 4080 1650
rect 4270 1640 4300 1650
rect 4320 1640 4430 1650
rect 4460 1640 4470 1650
rect 4540 1640 4550 1650
rect 4620 1640 4670 1650
rect 4710 1640 4760 1650
rect 4880 1640 4900 1650
rect 5280 1640 5290 1650
rect 6200 1640 6270 1650
rect 6650 1640 6800 1650
rect 7360 1640 7770 1650
rect 9120 1640 9220 1650
rect 9870 1640 9880 1650
rect 0 1630 560 1640
rect 870 1630 1910 1640
rect 3260 1630 4090 1640
rect 4280 1630 4300 1640
rect 4320 1630 4390 1640
rect 4450 1630 4470 1640
rect 4530 1630 4550 1640
rect 4620 1630 4660 1640
rect 4730 1630 4750 1640
rect 4850 1630 4880 1640
rect 5270 1630 5280 1640
rect 6200 1630 6270 1640
rect 6660 1630 6800 1640
rect 7360 1630 7770 1640
rect 9120 1630 9230 1640
rect 9860 1630 9880 1640
rect 0 1620 550 1630
rect 860 1620 1910 1630
rect 3250 1620 4090 1630
rect 4280 1620 4300 1630
rect 4320 1620 4360 1630
rect 4440 1620 4470 1630
rect 4500 1620 4540 1630
rect 5260 1620 5280 1630
rect 6200 1620 6280 1630
rect 6680 1620 6800 1630
rect 7360 1620 7770 1630
rect 9120 1620 9240 1630
rect 9860 1620 9870 1630
rect 0 1610 550 1620
rect 860 1610 1920 1620
rect 3250 1610 4090 1620
rect 4290 1610 4300 1620
rect 4320 1610 4350 1620
rect 4410 1610 4470 1620
rect 4990 1610 5020 1620
rect 5260 1610 5270 1620
rect 6210 1610 6280 1620
rect 6700 1610 6800 1620
rect 7360 1610 7780 1620
rect 9130 1610 9180 1620
rect 9850 1610 9870 1620
rect 0 1600 540 1610
rect 860 1600 1920 1610
rect 3240 1600 4100 1610
rect 4290 1600 4300 1610
rect 4320 1600 4350 1610
rect 4360 1600 4460 1610
rect 5250 1600 5270 1610
rect 6210 1600 6280 1610
rect 6710 1600 6800 1610
rect 7370 1600 7780 1610
rect 9130 1600 9150 1610
rect 9840 1600 9870 1610
rect 0 1590 540 1600
rect 860 1590 1920 1600
rect 3230 1590 4100 1600
rect 4330 1590 4450 1600
rect 4570 1590 4840 1600
rect 5250 1590 5260 1600
rect 6210 1590 6280 1600
rect 6720 1590 6800 1600
rect 7370 1590 7780 1600
rect 9840 1590 9860 1600
rect 0 1580 540 1590
rect 850 1580 1930 1590
rect 3220 1580 4100 1590
rect 4310 1580 4420 1590
rect 4500 1580 4610 1590
rect 4850 1580 4940 1590
rect 5230 1580 5250 1590
rect 5370 1580 5380 1590
rect 5500 1580 5510 1590
rect 6210 1580 6280 1590
rect 6730 1580 6800 1590
rect 7370 1580 7790 1590
rect 9830 1580 9860 1590
rect 0 1570 530 1580
rect 850 1570 1940 1580
rect 3220 1570 4110 1580
rect 4310 1570 4390 1580
rect 4440 1570 4520 1580
rect 4960 1570 4990 1580
rect 5200 1570 5230 1580
rect 5360 1570 5370 1580
rect 5420 1570 5430 1580
rect 6220 1570 6280 1580
rect 6730 1570 6800 1580
rect 7370 1570 7780 1580
rect 9830 1570 9840 1580
rect 9950 1570 9980 1580
rect 0 1560 530 1570
rect 850 1560 1940 1570
rect 3210 1560 4110 1570
rect 4320 1560 4490 1570
rect 4990 1560 5030 1570
rect 6220 1560 6290 1570
rect 6730 1560 6790 1570
rect 7370 1560 7780 1570
rect 9820 1560 9840 1570
rect 9930 1560 9990 1570
rect 0 1550 530 1560
rect 840 1550 1950 1560
rect 3210 1550 4120 1560
rect 4320 1550 4460 1560
rect 5050 1550 5080 1560
rect 5340 1550 5350 1560
rect 6220 1550 6290 1560
rect 6730 1550 6790 1560
rect 7370 1550 7790 1560
rect 9710 1550 9800 1560
rect 9820 1550 9830 1560
rect 9930 1550 9990 1560
rect 0 1540 520 1550
rect 840 1540 1960 1550
rect 3200 1540 4120 1550
rect 4330 1540 4430 1550
rect 4440 1540 4460 1550
rect 5100 1540 5110 1550
rect 5330 1540 5340 1550
rect 5630 1540 5650 1550
rect 6230 1540 6290 1550
rect 6730 1540 6790 1550
rect 7370 1540 7790 1550
rect 9710 1540 9790 1550
rect 9810 1540 9830 1550
rect 9930 1540 9990 1550
rect 0 1530 520 1540
rect 840 1530 1960 1540
rect 3190 1530 4130 1540
rect 4340 1530 4410 1540
rect 4440 1530 4470 1540
rect 5330 1530 5340 1540
rect 5630 1530 5640 1540
rect 6230 1530 6300 1540
rect 6730 1530 6790 1540
rect 7370 1530 7790 1540
rect 9710 1530 9790 1540
rect 9810 1530 9820 1540
rect 9940 1530 9950 1540
rect 9990 1530 9990 1540
rect 0 1520 520 1530
rect 830 1520 1970 1530
rect 3180 1520 4130 1530
rect 4340 1520 4400 1530
rect 4440 1520 4470 1530
rect 5320 1520 5330 1530
rect 6200 1520 6220 1530
rect 6230 1520 6300 1530
rect 6730 1520 6790 1530
rect 7380 1520 7790 1530
rect 9710 1520 9780 1530
rect 9800 1520 9830 1530
rect 9990 1520 9990 1530
rect 0 1510 510 1520
rect 840 1510 1980 1520
rect 3170 1510 4130 1520
rect 4350 1510 4390 1520
rect 4450 1510 4470 1520
rect 6200 1510 6220 1520
rect 6240 1510 6300 1520
rect 6760 1510 6790 1520
rect 7380 1510 7800 1520
rect 9710 1510 9780 1520
rect 9790 1510 9820 1520
rect 9980 1510 9990 1520
rect 0 1500 510 1510
rect 830 1500 1990 1510
rect 3160 1500 4130 1510
rect 4350 1500 4360 1510
rect 4380 1500 4390 1510
rect 4450 1500 4470 1510
rect 6200 1500 6300 1510
rect 6760 1500 6790 1510
rect 7380 1500 7800 1510
rect 9140 1500 9200 1510
rect 9720 1500 9770 1510
rect 9790 1500 9820 1510
rect 0 1490 510 1500
rect 830 1490 1990 1500
rect 3150 1490 4140 1500
rect 4350 1490 4370 1500
rect 4450 1490 4470 1500
rect 5230 1490 5240 1500
rect 6200 1490 6300 1500
rect 6770 1490 6790 1500
rect 7380 1490 7800 1500
rect 9130 1490 9190 1500
rect 9720 1490 9770 1500
rect 9780 1490 9810 1500
rect 9910 1490 9920 1500
rect 0 1480 500 1490
rect 830 1480 2000 1490
rect 3140 1480 4140 1490
rect 4360 1480 4380 1490
rect 4440 1480 4470 1490
rect 5250 1480 5260 1490
rect 6200 1480 6310 1490
rect 6770 1480 6790 1490
rect 7380 1480 7800 1490
rect 9130 1480 9180 1490
rect 9350 1480 9360 1490
rect 9720 1480 9760 1490
rect 9780 1480 9800 1490
rect 0 1470 500 1480
rect 840 1470 2010 1480
rect 3130 1470 4140 1480
rect 4360 1470 4380 1480
rect 4440 1470 4560 1480
rect 4980 1470 4990 1480
rect 6190 1470 6310 1480
rect 6760 1470 6790 1480
rect 7380 1470 7800 1480
rect 9130 1470 9180 1480
rect 9720 1470 9760 1480
rect 9770 1470 9800 1480
rect 0 1460 500 1470
rect 840 1460 900 1470
rect 990 1460 2020 1470
rect 3120 1460 4140 1470
rect 4370 1460 4380 1470
rect 4390 1460 4680 1470
rect 4980 1460 4990 1470
rect 6190 1460 6300 1470
rect 6760 1460 6790 1470
rect 7380 1460 7810 1470
rect 9130 1460 9170 1470
rect 9710 1460 9750 1470
rect 9760 1460 9790 1470
rect 0 1450 490 1460
rect 840 1450 880 1460
rect 1000 1450 2020 1460
rect 3110 1450 4150 1460
rect 4370 1450 4480 1460
rect 4500 1450 4520 1460
rect 4540 1450 4560 1460
rect 4580 1450 4600 1460
rect 4620 1450 4640 1460
rect 4650 1450 4680 1460
rect 4690 1450 4740 1460
rect 4850 1450 4880 1460
rect 5300 1450 5310 1460
rect 6200 1450 6310 1460
rect 6780 1450 6800 1460
rect 7380 1450 7810 1460
rect 9130 1450 9160 1460
rect 9590 1450 9630 1460
rect 9710 1450 9750 1460
rect 9760 1450 9780 1460
rect 0 1440 490 1450
rect 840 1440 860 1450
rect 1010 1440 2030 1450
rect 3100 1440 4150 1450
rect 4370 1440 4430 1450
rect 4450 1440 4480 1450
rect 4500 1440 4520 1450
rect 4540 1440 4560 1450
rect 4580 1440 4600 1450
rect 4620 1440 4640 1450
rect 4660 1440 4670 1450
rect 4690 1440 4710 1450
rect 4730 1440 4790 1450
rect 4850 1440 4880 1450
rect 4970 1440 4980 1450
rect 5310 1440 5320 1450
rect 6200 1440 6310 1450
rect 6780 1440 6800 1450
rect 7390 1440 7810 1450
rect 9140 1440 9150 1450
rect 9610 1440 9630 1450
rect 9710 1440 9740 1450
rect 9750 1440 9780 1450
rect 0 1430 490 1440
rect 840 1430 860 1440
rect 1020 1430 2040 1440
rect 3090 1430 4150 1440
rect 4370 1430 4430 1440
rect 4460 1430 4470 1440
rect 4500 1430 4520 1440
rect 4540 1430 4560 1440
rect 4580 1430 4600 1440
rect 4620 1430 4630 1440
rect 4650 1430 4670 1440
rect 4690 1430 4710 1440
rect 4730 1430 4740 1440
rect 4760 1430 4830 1440
rect 4850 1430 4860 1440
rect 4870 1430 4880 1440
rect 4970 1430 4980 1440
rect 5320 1430 5330 1440
rect 6200 1430 6310 1440
rect 6780 1430 6800 1440
rect 7390 1430 7820 1440
rect 9620 1430 9630 1440
rect 9700 1430 9730 1440
rect 9750 1430 9780 1440
rect 0 1420 480 1430
rect 840 1420 850 1430
rect 1020 1420 2050 1430
rect 3080 1420 4160 1430
rect 4380 1420 4400 1430
rect 4410 1420 4440 1430
rect 4460 1420 4470 1430
rect 4500 1420 4520 1430
rect 4540 1420 4560 1430
rect 4580 1420 4600 1430
rect 4620 1420 4630 1430
rect 4660 1420 4670 1430
rect 4690 1420 4710 1430
rect 4720 1420 4740 1430
rect 4760 1420 4780 1430
rect 4800 1420 4810 1430
rect 4820 1420 4860 1430
rect 4870 1420 4890 1430
rect 4970 1420 4980 1430
rect 5330 1420 5340 1430
rect 6200 1420 6310 1430
rect 6780 1420 6800 1430
rect 7390 1420 7820 1430
rect 9700 1420 9730 1430
rect 9740 1420 9760 1430
rect 0 1410 480 1420
rect 1030 1410 2060 1420
rect 3070 1410 4160 1420
rect 4380 1410 4440 1420
rect 4460 1410 4480 1420
rect 4500 1410 4520 1420
rect 4540 1410 4560 1420
rect 4580 1410 4640 1420
rect 4650 1410 4680 1420
rect 4690 1410 4710 1420
rect 4720 1410 4740 1420
rect 4760 1410 4770 1420
rect 4800 1410 4810 1420
rect 4840 1410 4850 1420
rect 4870 1410 4890 1420
rect 6200 1410 6310 1420
rect 6790 1410 6800 1420
rect 7390 1410 7820 1420
rect 9700 1410 9720 1420
rect 9740 1410 9760 1420
rect 0 1400 480 1410
rect 1030 1400 2060 1410
rect 3060 1400 4160 1410
rect 4390 1400 4440 1410
rect 4460 1400 4480 1410
rect 4500 1400 4520 1410
rect 4530 1400 4740 1410
rect 4760 1400 4770 1410
rect 4790 1400 4800 1410
rect 4870 1400 4890 1410
rect 5350 1400 5360 1410
rect 6200 1400 6310 1410
rect 6790 1400 6800 1410
rect 7390 1400 7820 1410
rect 9700 1400 9720 1410
rect 9730 1400 9760 1410
rect 0 1390 470 1400
rect 1030 1390 2070 1400
rect 3050 1390 4170 1400
rect 4390 1390 4440 1400
rect 4460 1390 4550 1400
rect 4740 1390 4780 1400
rect 4790 1390 4800 1400
rect 4830 1390 4840 1400
rect 4870 1390 4880 1400
rect 4890 1390 4900 1400
rect 6200 1390 6310 1400
rect 6790 1390 6800 1400
rect 7390 1390 7820 1400
rect 9230 1390 9250 1400
rect 9690 1390 9710 1400
rect 9730 1390 9750 1400
rect 0 1380 470 1390
rect 1020 1380 2080 1390
rect 3030 1380 4170 1390
rect 4400 1380 4500 1390
rect 4780 1380 4840 1390
rect 4860 1380 4870 1390
rect 4890 1380 4900 1390
rect 4920 1380 4940 1390
rect 4960 1380 4970 1390
rect 6200 1380 6310 1390
rect 6790 1380 6800 1390
rect 7390 1380 7820 1390
rect 9220 1380 9260 1390
rect 9690 1380 9710 1390
rect 9720 1380 9750 1390
rect 0 1370 470 1380
rect 1020 1370 2080 1380
rect 3020 1370 4170 1380
rect 4400 1370 4460 1380
rect 4480 1370 4500 1380
rect 4820 1370 4840 1380
rect 4860 1370 4870 1380
rect 4920 1370 4950 1380
rect 4960 1370 4970 1380
rect 5600 1370 5610 1380
rect 6200 1370 6310 1380
rect 6790 1370 6810 1380
rect 7400 1370 7830 1380
rect 9210 1370 9250 1380
rect 9680 1370 9700 1380
rect 9710 1370 9740 1380
rect 9970 1370 9990 1380
rect 0 1360 470 1370
rect 1020 1360 2080 1370
rect 3010 1360 4180 1370
rect 4400 1360 4430 1370
rect 4480 1360 4510 1370
rect 4830 1360 4840 1370
rect 4860 1360 4890 1370
rect 4930 1360 4940 1370
rect 4960 1360 4970 1370
rect 5400 1360 5410 1370
rect 5590 1360 5600 1370
rect 6200 1360 6310 1370
rect 6790 1360 6810 1370
rect 7400 1360 7830 1370
rect 9200 1360 9260 1370
rect 9680 1360 9690 1370
rect 9710 1360 9740 1370
rect 9970 1360 9990 1370
rect 0 1350 460 1360
rect 1020 1350 2080 1360
rect 2990 1350 3560 1360
rect 3610 1350 4180 1360
rect 4410 1350 4420 1360
rect 4480 1350 4510 1360
rect 4830 1350 4840 1360
rect 4860 1350 4870 1360
rect 4960 1350 4970 1360
rect 5410 1350 5420 1360
rect 6200 1350 6310 1360
rect 6790 1350 6810 1360
rect 7400 1350 7830 1360
rect 9190 1350 9260 1360
rect 9680 1350 9690 1360
rect 9700 1350 9740 1360
rect 9810 1350 9820 1360
rect 9970 1350 9990 1360
rect 0 1340 460 1350
rect 820 1340 830 1350
rect 1020 1340 2090 1350
rect 2980 1340 3540 1350
rect 3630 1340 4180 1350
rect 4490 1340 4510 1350
rect 4830 1340 4850 1350
rect 5420 1340 5430 1350
rect 6200 1340 6310 1350
rect 6790 1340 6810 1350
rect 7400 1340 7830 1350
rect 9180 1340 9260 1350
rect 9650 1340 9670 1350
rect 9700 1340 9730 1350
rect 9810 1340 9830 1350
rect 9970 1340 9990 1350
rect 0 1330 460 1340
rect 1020 1330 2080 1340
rect 2970 1330 3530 1340
rect 3650 1330 4190 1340
rect 4490 1330 4510 1340
rect 5430 1330 5440 1340
rect 6200 1330 6310 1340
rect 6800 1330 6810 1340
rect 7400 1330 7830 1340
rect 9170 1330 9260 1340
rect 9650 1330 9670 1340
rect 9690 1330 9720 1340
rect 9800 1330 9830 1340
rect 9990 1330 9990 1340
rect 0 1320 450 1330
rect 1020 1320 2080 1330
rect 2960 1320 3520 1330
rect 3660 1320 4190 1330
rect 4490 1320 4510 1330
rect 5440 1320 5450 1330
rect 6200 1320 6310 1330
rect 6800 1320 6820 1330
rect 7400 1320 7830 1330
rect 9160 1320 9260 1330
rect 9650 1320 9670 1330
rect 9690 1320 9710 1330
rect 9770 1320 9830 1330
rect 0 1310 450 1320
rect 810 1310 820 1320
rect 1020 1310 2080 1320
rect 2930 1310 3510 1320
rect 3670 1310 4190 1320
rect 4500 1310 4510 1320
rect 5450 1310 5460 1320
rect 6200 1310 6320 1320
rect 6810 1310 6820 1320
rect 7400 1310 7840 1320
rect 9150 1310 9260 1320
rect 9680 1310 9710 1320
rect 9770 1310 9830 1320
rect 0 1300 450 1310
rect 810 1300 820 1310
rect 1020 1300 2080 1310
rect 2920 1300 3510 1310
rect 3680 1300 4200 1310
rect 4500 1300 4520 1310
rect 5450 1300 5470 1310
rect 6200 1300 6320 1310
rect 6800 1300 6810 1310
rect 7400 1300 7830 1310
rect 9140 1300 9260 1310
rect 9680 1300 9700 1310
rect 9770 1300 9780 1310
rect 9800 1300 9810 1310
rect 0 1290 440 1300
rect 1010 1290 2070 1300
rect 2910 1290 3510 1300
rect 3700 1290 4200 1300
rect 4500 1290 4520 1300
rect 5450 1290 5480 1300
rect 5490 1290 5510 1300
rect 5550 1290 5560 1300
rect 5590 1290 5680 1300
rect 6210 1290 6320 1300
rect 6790 1290 6820 1300
rect 7410 1290 7840 1300
rect 9140 1290 9260 1300
rect 9670 1290 9700 1300
rect 9770 1290 9780 1300
rect 9800 1290 9820 1300
rect 0 1280 440 1290
rect 1010 1280 2040 1290
rect 2890 1280 3500 1290
rect 3710 1280 4200 1290
rect 4500 1280 4520 1290
rect 4950 1280 4960 1290
rect 5300 1280 5370 1290
rect 6210 1280 6310 1290
rect 6790 1280 6820 1290
rect 7410 1280 7840 1290
rect 9140 1280 9260 1290
rect 9670 1280 9690 1290
rect 9760 1280 9790 1290
rect 9800 1280 9820 1290
rect 9960 1280 9970 1290
rect 0 1270 440 1280
rect 1010 1270 2040 1280
rect 2880 1270 3500 1280
rect 3720 1270 4200 1280
rect 4500 1270 4520 1280
rect 4950 1270 4960 1280
rect 5160 1270 5200 1280
rect 5230 1270 5250 1280
rect 6210 1270 6310 1280
rect 6790 1270 6820 1280
rect 7410 1270 7850 1280
rect 9140 1270 9310 1280
rect 9660 1270 9690 1280
rect 9750 1270 9760 1280
rect 9770 1270 9820 1280
rect 9960 1270 9980 1280
rect 0 1260 430 1270
rect 1010 1260 2040 1270
rect 2860 1260 3500 1270
rect 3730 1260 4200 1270
rect 4510 1260 4530 1270
rect 5090 1260 5120 1270
rect 6210 1260 6310 1270
rect 6790 1260 6820 1270
rect 7410 1260 7850 1270
rect 9140 1260 9310 1270
rect 9660 1260 9680 1270
rect 9750 1260 9760 1270
rect 9770 1260 9830 1270
rect 0 1250 430 1260
rect 1010 1250 2040 1260
rect 2840 1250 3500 1260
rect 3740 1250 4200 1260
rect 4510 1250 4530 1260
rect 4940 1250 4950 1260
rect 5020 1250 5070 1260
rect 6220 1250 6310 1260
rect 6790 1250 6820 1260
rect 7410 1250 7850 1260
rect 9140 1250 9310 1260
rect 9650 1250 9670 1260
rect 9760 1250 9830 1260
rect 0 1240 430 1250
rect 1010 1240 2030 1250
rect 2820 1240 3510 1250
rect 3760 1240 4200 1250
rect 4510 1240 4530 1250
rect 4940 1240 5010 1250
rect 6230 1240 6310 1250
rect 6800 1240 6820 1250
rect 7410 1240 7850 1250
rect 9140 1240 9280 1250
rect 9600 1240 9610 1250
rect 9640 1240 9670 1250
rect 9770 1240 9820 1250
rect 9990 1240 9990 1250
rect 0 1230 420 1240
rect 1010 1230 2030 1240
rect 2800 1230 3510 1240
rect 3770 1230 4200 1240
rect 4520 1230 4530 1240
rect 4930 1230 4950 1240
rect 5680 1230 5690 1240
rect 6230 1230 6310 1240
rect 6800 1230 6820 1240
rect 7410 1230 7860 1240
rect 9140 1230 9280 1240
rect 9640 1230 9660 1240
rect 9730 1230 9750 1240
rect 9780 1230 9820 1240
rect 9970 1230 9990 1240
rect 0 1220 420 1230
rect 1000 1220 2030 1230
rect 2780 1220 3520 1230
rect 3790 1220 4210 1230
rect 4520 1220 4530 1230
rect 4790 1220 4870 1230
rect 5680 1220 5690 1230
rect 6240 1220 6310 1230
rect 6360 1220 6370 1230
rect 6800 1220 6820 1230
rect 7410 1220 7860 1230
rect 9140 1220 9280 1230
rect 9500 1220 9520 1230
rect 9630 1220 9660 1230
rect 9730 1220 9760 1230
rect 9800 1220 9820 1230
rect 9970 1220 9990 1230
rect 0 1210 420 1220
rect 790 1210 800 1220
rect 1000 1210 2020 1220
rect 2760 1210 3520 1220
rect 3810 1210 4210 1220
rect 4520 1210 4540 1220
rect 4680 1210 4790 1220
rect 6240 1210 6360 1220
rect 6800 1210 6820 1220
rect 7410 1210 7860 1220
rect 9140 1210 9280 1220
rect 9510 1210 9530 1220
rect 9630 1210 9650 1220
rect 9720 1210 9760 1220
rect 9970 1210 9990 1220
rect 0 1200 410 1210
rect 980 1200 990 1210
rect 1000 1200 2020 1210
rect 2750 1200 3530 1210
rect 3820 1200 4210 1210
rect 4520 1200 4540 1210
rect 4570 1200 4700 1210
rect 6250 1200 6380 1210
rect 6800 1200 6820 1210
rect 7420 1200 7860 1210
rect 9150 1200 9280 1210
rect 9510 1200 9530 1210
rect 9620 1200 9650 1210
rect 9710 1200 9770 1210
rect 9970 1200 9990 1210
rect 0 1190 410 1200
rect 980 1190 2010 1200
rect 2740 1190 3540 1200
rect 3840 1190 4210 1200
rect 4450 1190 4470 1200
rect 4480 1190 4610 1200
rect 5690 1190 5700 1200
rect 6250 1190 6390 1200
rect 6800 1190 6820 1200
rect 7420 1190 7870 1200
rect 9140 1190 9280 1200
rect 9310 1190 9320 1200
rect 9510 1190 9540 1200
rect 9620 1190 9640 1200
rect 9710 1190 9770 1200
rect 9780 1190 9810 1200
rect 0 1180 410 1190
rect 960 1180 2010 1190
rect 2730 1180 3550 1190
rect 3850 1180 4210 1190
rect 4450 1180 4540 1190
rect 5680 1180 5700 1190
rect 6250 1180 6390 1190
rect 6810 1180 6820 1190
rect 7420 1180 7870 1190
rect 9150 1180 9280 1190
rect 9320 1180 9350 1190
rect 9510 1180 9540 1190
rect 9610 1180 9640 1190
rect 9710 1180 9760 1190
rect 9780 1180 9810 1190
rect 0 1170 400 1180
rect 960 1170 980 1180
rect 990 1170 2010 1180
rect 2740 1170 2750 1180
rect 2830 1170 3550 1180
rect 3860 1170 4210 1180
rect 6250 1170 6370 1180
rect 6810 1170 6820 1180
rect 7420 1170 7870 1180
rect 9150 1170 9280 1180
rect 9320 1170 9360 1180
rect 9510 1170 9540 1180
rect 9600 1170 9630 1180
rect 9710 1170 9760 1180
rect 9770 1170 9810 1180
rect 0 1160 400 1170
rect 990 1160 2010 1170
rect 2850 1160 3560 1170
rect 3880 1160 4210 1170
rect 5690 1160 5700 1170
rect 6250 1160 6380 1170
rect 6810 1160 6820 1170
rect 7420 1160 7880 1170
rect 9150 1160 9280 1170
rect 9330 1160 9360 1170
rect 9520 1160 9550 1170
rect 9600 1160 9630 1170
rect 9710 1160 9800 1170
rect 0 1150 390 1160
rect 640 1150 660 1160
rect 670 1150 680 1160
rect 990 1150 2010 1160
rect 2850 1150 3570 1160
rect 3890 1150 4220 1160
rect 5690 1150 5700 1160
rect 6250 1150 6380 1160
rect 6810 1150 6820 1160
rect 7420 1150 7870 1160
rect 9160 1150 9290 1160
rect 9330 1150 9370 1160
rect 9520 1150 9550 1160
rect 9590 1150 9620 1160
rect 9720 1150 9820 1160
rect 0 1140 390 1150
rect 610 1140 680 1150
rect 760 1140 770 1150
rect 980 1140 2010 1150
rect 2870 1140 3580 1150
rect 3900 1140 4220 1150
rect 5690 1140 5700 1150
rect 6260 1140 6380 1150
rect 6810 1140 6820 1150
rect 7420 1140 7880 1150
rect 9160 1140 9290 1150
rect 9330 1140 9380 1150
rect 9590 1140 9610 1150
rect 9720 1140 9820 1150
rect 0 1130 390 1140
rect 620 1130 750 1140
rect 990 1130 2000 1140
rect 2880 1130 3590 1140
rect 3920 1130 4220 1140
rect 5690 1130 5700 1140
rect 6260 1130 6410 1140
rect 6810 1130 6830 1140
rect 7420 1130 7880 1140
rect 9160 1130 9290 1140
rect 9350 1130 9380 1140
rect 9580 1130 9610 1140
rect 9720 1130 9820 1140
rect 0 1120 380 1130
rect 630 1120 760 1130
rect 990 1120 2000 1130
rect 2890 1120 3600 1130
rect 3930 1120 4220 1130
rect 5690 1120 5700 1130
rect 6260 1120 6400 1130
rect 6810 1120 6830 1130
rect 7420 1120 7880 1130
rect 9150 1120 9290 1130
rect 9350 1120 9390 1130
rect 9570 1120 9600 1130
rect 9730 1120 9820 1130
rect 0 1110 380 1120
rect 610 1110 750 1120
rect 990 1110 1990 1120
rect 2890 1110 3610 1120
rect 3940 1110 4220 1120
rect 5690 1110 5700 1120
rect 6260 1110 6400 1120
rect 6810 1110 6830 1120
rect 7420 1110 7880 1120
rect 9150 1110 9290 1120
rect 9370 1110 9390 1120
rect 9570 1110 9600 1120
rect 9730 1110 9810 1120
rect 0 1100 380 1110
rect 610 1100 750 1110
rect 980 1100 1570 1110
rect 1610 1100 1990 1110
rect 2890 1100 3620 1110
rect 3960 1100 4110 1110
rect 4120 1100 4220 1110
rect 5690 1100 5700 1110
rect 6270 1100 6400 1110
rect 6820 1100 6830 1110
rect 7420 1100 7880 1110
rect 9150 1100 9290 1110
rect 9360 1100 9390 1110
rect 9560 1100 9590 1110
rect 9730 1100 9820 1110
rect 0 1090 370 1100
rect 620 1090 750 1100
rect 980 1090 1540 1100
rect 1630 1090 1990 1100
rect 2890 1090 3630 1100
rect 3980 1090 4100 1100
rect 4130 1090 4220 1100
rect 6270 1090 6420 1100
rect 6810 1090 6830 1100
rect 7420 1090 7880 1100
rect 9150 1090 9230 1100
rect 9280 1090 9290 1100
rect 9370 1090 9410 1100
rect 9560 1090 9580 1100
rect 9730 1090 9820 1100
rect 0 1080 370 1090
rect 620 1080 750 1090
rect 980 1080 1530 1090
rect 1640 1080 1990 1090
rect 2900 1080 3650 1090
rect 3990 1080 4090 1090
rect 4110 1080 4220 1090
rect 5690 1080 5700 1090
rect 6270 1080 6430 1090
rect 6820 1080 6830 1090
rect 7430 1080 7890 1090
rect 9160 1080 9180 1090
rect 9280 1080 9290 1090
rect 9370 1080 9410 1090
rect 9550 1080 9570 1090
rect 9730 1080 9830 1090
rect 9960 1080 9970 1090
rect 9980 1080 9990 1090
rect 0 1070 360 1080
rect 620 1070 750 1080
rect 980 1070 1510 1080
rect 1650 1070 1980 1080
rect 2910 1070 3660 1080
rect 4020 1070 4100 1080
rect 4110 1070 4220 1080
rect 5680 1070 5700 1080
rect 6270 1070 6460 1080
rect 6470 1070 6480 1080
rect 6820 1070 6830 1080
rect 7430 1070 7890 1080
rect 9270 1070 9300 1080
rect 9370 1070 9410 1080
rect 9550 1070 9560 1080
rect 9730 1070 9830 1080
rect 9950 1070 9990 1080
rect 0 1060 360 1070
rect 630 1060 740 1070
rect 980 1060 1500 1070
rect 1650 1060 1980 1070
rect 2900 1060 3670 1070
rect 4030 1060 4070 1070
rect 4080 1060 4100 1070
rect 4130 1060 4220 1070
rect 5690 1060 5700 1070
rect 6270 1060 6450 1070
rect 6820 1060 6830 1070
rect 7430 1060 7900 1070
rect 9260 1060 9300 1070
rect 9370 1060 9420 1070
rect 9540 1060 9560 1070
rect 9730 1060 9830 1070
rect 9950 1060 9990 1070
rect 0 1050 350 1060
rect 630 1050 740 1060
rect 970 1050 1490 1060
rect 1650 1050 1990 1060
rect 2900 1050 3670 1060
rect 4040 1050 4070 1060
rect 4080 1050 4090 1060
rect 4130 1050 4220 1060
rect 5690 1050 5700 1060
rect 6280 1050 6440 1060
rect 6820 1050 6830 1060
rect 7430 1050 7900 1060
rect 9260 1050 9300 1060
rect 9370 1050 9420 1060
rect 9540 1050 9550 1060
rect 9720 1050 9800 1060
rect 9820 1050 9840 1060
rect 9970 1050 9980 1060
rect 0 1040 350 1050
rect 630 1040 740 1050
rect 970 1040 1480 1050
rect 1660 1040 1980 1050
rect 2900 1040 3680 1050
rect 4080 1040 4110 1050
rect 4120 1040 4200 1050
rect 5690 1040 5700 1050
rect 6280 1040 6410 1050
rect 6820 1040 6830 1050
rect 7430 1040 7900 1050
rect 9130 1040 9140 1050
rect 9250 1040 9300 1050
rect 9380 1040 9420 1050
rect 9530 1040 9560 1050
rect 9730 1040 9820 1050
rect 0 1030 340 1040
rect 630 1030 730 1040
rect 970 1030 1470 1040
rect 1650 1030 1980 1040
rect 2900 1030 3690 1040
rect 4070 1030 4200 1040
rect 4210 1030 4220 1040
rect 5690 1030 5700 1040
rect 6290 1030 6400 1040
rect 6820 1030 6830 1040
rect 7430 1030 7900 1040
rect 9120 1030 9140 1040
rect 9250 1030 9290 1040
rect 9380 1030 9420 1040
rect 9530 1030 9560 1040
rect 9740 1030 9820 1040
rect 0 1020 340 1030
rect 650 1020 730 1030
rect 960 1020 1460 1030
rect 1650 1020 1980 1030
rect 2900 1020 3700 1030
rect 4090 1020 4200 1030
rect 4210 1020 4220 1030
rect 5690 1020 5700 1030
rect 6290 1020 6370 1030
rect 6820 1020 6830 1030
rect 7430 1020 7910 1030
rect 9120 1020 9140 1030
rect 9380 1020 9430 1030
rect 9520 1020 9530 1030
rect 9740 1020 9830 1030
rect 0 1010 330 1020
rect 670 1010 730 1020
rect 960 1010 1450 1020
rect 1650 1010 1980 1020
rect 2900 1010 3710 1020
rect 4110 1010 4210 1020
rect 5680 1010 5700 1020
rect 6290 1010 6360 1020
rect 6820 1010 6830 1020
rect 7430 1010 7900 1020
rect 9130 1010 9140 1020
rect 9390 1010 9430 1020
rect 9510 1010 9530 1020
rect 9740 1010 9790 1020
rect 9810 1010 9820 1020
rect 0 1000 330 1010
rect 670 1000 680 1010
rect 690 1000 720 1010
rect 960 1000 1440 1010
rect 1650 1000 1980 1010
rect 2890 1000 3720 1010
rect 4120 1000 4190 1010
rect 4200 1000 4210 1010
rect 5680 1000 5700 1010
rect 6300 1000 6360 1010
rect 6820 1000 6830 1010
rect 7430 1000 7900 1010
rect 9130 1000 9140 1010
rect 9410 1000 9420 1010
rect 9510 1000 9520 1010
rect 9740 1000 9780 1010
rect 9810 1000 9820 1010
rect 0 990 320 1000
rect 680 990 720 1000
rect 960 990 1430 1000
rect 1640 990 1980 1000
rect 2890 990 3730 1000
rect 4140 990 4170 1000
rect 4180 990 4200 1000
rect 5690 990 5700 1000
rect 6300 990 6350 1000
rect 7430 990 7910 1000
rect 9130 990 9140 1000
rect 9500 990 9520 1000
rect 9740 990 9770 1000
rect 9810 990 9820 1000
rect 0 980 320 990
rect 680 980 690 990
rect 700 980 720 990
rect 950 980 1420 990
rect 1630 980 1980 990
rect 2890 980 3740 990
rect 4170 980 4190 990
rect 5690 980 5700 990
rect 6300 980 6350 990
rect 7430 980 7920 990
rect 9130 980 9150 990
rect 9500 980 9510 990
rect 9770 980 9780 990
rect 0 970 310 980
rect 700 970 710 980
rect 950 970 1400 980
rect 1610 970 1980 980
rect 2880 970 3750 980
rect 5680 970 5700 980
rect 6300 970 6350 980
rect 7430 970 7920 980
rect 9130 970 9150 980
rect 9490 970 9500 980
rect 9770 970 9780 980
rect 0 960 310 970
rect 950 960 1390 970
rect 1600 960 1980 970
rect 2870 960 3760 970
rect 5030 960 5040 970
rect 5680 960 5690 970
rect 6300 960 6350 970
rect 7430 960 7920 970
rect 9130 960 9140 970
rect 9480 960 9510 970
rect 0 950 300 960
rect 940 950 1380 960
rect 1590 950 1980 960
rect 2850 950 3770 960
rect 4900 950 5090 960
rect 6300 950 6360 960
rect 7430 950 7920 960
rect 9120 950 9140 960
rect 9210 950 9250 960
rect 9480 950 9510 960
rect 0 940 300 950
rect 930 940 1360 950
rect 1590 940 1980 950
rect 2850 940 3780 950
rect 4850 940 5140 950
rect 6300 940 6360 950
rect 7430 940 7920 950
rect 9120 940 9160 950
rect 9220 940 9260 950
rect 9470 940 9510 950
rect 0 930 290 940
rect 940 930 1350 940
rect 1570 930 1980 940
rect 2840 930 3790 940
rect 4820 930 5010 940
rect 5020 930 5190 940
rect 6300 930 6370 940
rect 7430 930 7920 940
rect 9120 930 9160 940
rect 9220 930 9250 940
rect 9470 930 9490 940
rect 0 920 280 930
rect 940 920 1340 930
rect 1570 920 1990 930
rect 2820 920 3800 930
rect 4830 920 4910 930
rect 4920 920 4950 930
rect 5080 920 5210 930
rect 6300 920 6370 930
rect 7430 920 7920 930
rect 9120 920 9170 930
rect 9460 920 9490 930
rect 0 910 280 920
rect 940 910 1330 920
rect 1560 910 1990 920
rect 2800 910 3810 920
rect 4840 910 4870 920
rect 5130 910 5250 920
rect 6300 910 6380 920
rect 7430 910 7930 920
rect 9120 910 9170 920
rect 9460 910 9480 920
rect 0 900 270 910
rect 930 900 1310 910
rect 1550 900 1990 910
rect 2780 900 3820 910
rect 4840 900 4870 910
rect 4920 900 5000 910
rect 5170 900 5250 910
rect 5680 900 5700 910
rect 6290 900 6370 910
rect 6830 900 6840 910
rect 7430 900 7930 910
rect 9120 900 9170 910
rect 9450 900 9470 910
rect 0 890 260 900
rect 940 890 1300 900
rect 1540 890 1990 900
rect 2770 890 3830 900
rect 4880 890 5080 900
rect 5180 890 5280 900
rect 5690 890 5700 900
rect 6290 890 6370 900
rect 7430 890 7930 900
rect 9120 890 9170 900
rect 9450 890 9470 900
rect 0 880 260 890
rect 930 880 1290 890
rect 1530 880 2000 890
rect 2750 880 3840 890
rect 4860 880 5110 890
rect 5180 880 5290 890
rect 5690 880 5700 890
rect 6290 880 6380 890
rect 7430 880 7930 890
rect 9120 880 9170 890
rect 9440 880 9470 890
rect 0 870 250 880
rect 930 870 1280 880
rect 1520 870 2000 880
rect 2730 870 3840 880
rect 4860 870 5170 880
rect 5190 870 5300 880
rect 5690 870 5700 880
rect 6290 870 6380 880
rect 7430 870 7930 880
rect 9120 870 9180 880
rect 9430 870 9470 880
rect 0 860 240 870
rect 930 860 1260 870
rect 1500 860 2000 870
rect 2710 860 3850 870
rect 4870 860 5190 870
rect 5220 860 5240 870
rect 5260 860 5320 870
rect 5690 860 5700 870
rect 6290 860 6390 870
rect 7430 860 7930 870
rect 9120 860 9180 870
rect 9430 860 9460 870
rect 0 850 240 860
rect 930 850 1250 860
rect 1490 850 2010 860
rect 2690 850 3860 860
rect 4880 850 4960 860
rect 4990 850 5060 860
rect 5080 850 5210 860
rect 5270 850 5340 860
rect 5670 850 5700 860
rect 6290 850 6390 860
rect 7430 850 7930 860
rect 9120 850 9180 860
rect 9420 850 9450 860
rect 0 840 230 850
rect 930 840 1240 850
rect 1490 840 2010 850
rect 2670 840 3870 850
rect 4880 840 5010 850
rect 5030 840 5060 850
rect 5080 840 5220 850
rect 5280 840 5350 850
rect 5610 840 5700 850
rect 6290 840 6400 850
rect 7430 840 7940 850
rect 9120 840 9190 850
rect 9420 840 9450 850
rect 0 830 220 840
rect 920 830 1220 840
rect 1470 830 2020 840
rect 2650 830 3880 840
rect 4890 830 5010 840
rect 5040 830 5230 840
rect 5290 830 5360 840
rect 5610 830 5630 840
rect 5690 830 5700 840
rect 6290 830 6410 840
rect 7430 830 7940 840
rect 9120 830 9190 840
rect 9410 830 9430 840
rect 0 820 210 830
rect 920 820 1210 830
rect 1470 820 2020 830
rect 2630 820 3900 830
rect 4890 820 4920 830
rect 4930 820 5130 830
rect 5150 820 5170 830
rect 5180 820 5240 830
rect 5310 820 5370 830
rect 5690 820 5700 830
rect 6290 820 6410 830
rect 7430 820 7940 830
rect 9120 820 9190 830
rect 9400 820 9430 830
rect 0 810 200 820
rect 920 810 1200 820
rect 1470 810 2020 820
rect 2610 810 3910 820
rect 4900 810 5140 820
rect 5150 810 5160 820
rect 5200 810 5250 820
rect 5260 810 5270 820
rect 5320 810 5360 820
rect 5370 810 5380 820
rect 5690 810 5700 820
rect 6300 810 6410 820
rect 7430 810 7940 820
rect 9120 810 9200 820
rect 9400 810 9420 820
rect 0 800 190 810
rect 920 800 1180 810
rect 1480 800 2030 810
rect 2590 800 3920 810
rect 4900 800 5090 810
rect 5120 800 5170 810
rect 5240 800 5250 810
rect 5320 800 5390 810
rect 5690 800 5700 810
rect 6300 800 6410 810
rect 7430 800 7940 810
rect 9110 800 9200 810
rect 9390 800 9420 810
rect 0 790 180 800
rect 920 790 1170 800
rect 1480 790 2030 800
rect 2570 790 3930 800
rect 4910 790 5210 800
rect 5250 790 5270 800
rect 5350 790 5400 800
rect 5690 790 5700 800
rect 6300 790 6420 800
rect 7430 790 7950 800
rect 9110 790 9200 800
rect 9390 790 9420 800
rect 0 780 170 790
rect 910 780 1150 790
rect 1470 780 2040 790
rect 2550 780 3660 790
rect 3680 780 3950 790
rect 4910 780 5220 790
rect 5250 780 5310 790
rect 5350 780 5400 790
rect 5690 780 5700 790
rect 6310 780 6420 790
rect 7430 780 7950 790
rect 8150 780 8160 790
rect 9110 780 9200 790
rect 9380 780 9410 790
rect 0 770 160 780
rect 910 770 1140 780
rect 1460 770 2050 780
rect 2530 770 3660 780
rect 3740 770 3970 780
rect 4910 770 5230 780
rect 5250 770 5320 780
rect 5360 770 5410 780
rect 5690 770 5700 780
rect 6310 770 6410 780
rect 7430 770 7950 780
rect 8150 770 8160 780
rect 9110 770 9200 780
rect 9380 770 9410 780
rect 0 760 150 770
rect 900 760 1130 770
rect 1450 760 2050 770
rect 2510 760 3570 770
rect 3850 760 3990 770
rect 4920 760 5270 770
rect 5290 760 5330 770
rect 5350 760 5420 770
rect 5690 760 5700 770
rect 6310 760 6420 770
rect 7430 760 7950 770
rect 8150 760 8160 770
rect 9110 760 9210 770
rect 9370 760 9400 770
rect 0 750 140 760
rect 900 750 1110 760
rect 1440 750 2050 760
rect 2500 750 3530 760
rect 3880 750 3990 760
rect 4920 750 5170 760
rect 5190 750 5280 760
rect 5300 750 5340 760
rect 5360 750 5430 760
rect 5690 750 5700 760
rect 6320 750 6430 760
rect 7430 750 7960 760
rect 8150 750 8160 760
rect 9110 750 9210 760
rect 9360 750 9400 760
rect 0 740 130 750
rect 900 740 1100 750
rect 1420 740 2060 750
rect 2480 740 3450 750
rect 3900 740 4000 750
rect 4920 740 5290 750
rect 5320 740 5350 750
rect 5360 740 5440 750
rect 5690 740 5700 750
rect 6320 740 6430 750
rect 7430 740 7960 750
rect 8150 740 8160 750
rect 9110 740 9120 750
rect 9130 740 9220 750
rect 9360 740 9390 750
rect 0 730 120 740
rect 890 730 1090 740
rect 1410 730 2060 740
rect 2470 730 3420 740
rect 3910 730 4000 740
rect 4920 730 5360 740
rect 5380 730 5450 740
rect 5690 730 5700 740
rect 6320 730 6430 740
rect 7430 730 7970 740
rect 9110 730 9120 740
rect 9140 730 9210 740
rect 9350 730 9390 740
rect 0 720 110 730
rect 900 720 1080 730
rect 1410 720 2070 730
rect 2450 720 3400 730
rect 3920 720 4010 730
rect 4920 720 5150 730
rect 5170 720 5180 730
rect 5200 720 5370 730
rect 5380 720 5460 730
rect 5690 720 5700 730
rect 6330 720 6440 730
rect 7430 720 7970 730
rect 9110 720 9120 730
rect 9140 720 9210 730
rect 9350 720 9380 730
rect 0 710 90 720
rect 890 710 1060 720
rect 1400 710 2070 720
rect 2430 710 3380 720
rect 3930 710 4020 720
rect 4920 710 5050 720
rect 5060 710 5130 720
rect 5190 710 5370 720
rect 5390 710 5470 720
rect 5690 710 5700 720
rect 6330 710 6460 720
rect 7430 710 7970 720
rect 9120 710 9210 720
rect 9340 710 9380 720
rect 0 700 80 710
rect 910 700 1040 710
rect 1390 700 2080 710
rect 2420 700 3360 710
rect 3940 700 4010 710
rect 4930 700 5050 710
rect 5060 700 5140 710
rect 5200 700 5250 710
rect 5260 700 5350 710
rect 5360 700 5380 710
rect 5400 700 5480 710
rect 5690 700 5700 710
rect 6330 700 6460 710
rect 7430 700 7980 710
rect 9120 700 9210 710
rect 9340 700 9370 710
rect 0 690 60 700
rect 910 690 1030 700
rect 1380 690 2080 700
rect 2400 690 3350 700
rect 4930 690 5140 700
rect 5200 690 5390 700
rect 5410 690 5490 700
rect 5690 690 5700 700
rect 6330 690 6460 700
rect 7420 690 7980 700
rect 9120 690 9210 700
rect 9330 690 9360 700
rect 0 680 50 690
rect 920 680 1010 690
rect 1360 680 2090 690
rect 2380 680 3330 690
rect 4930 680 5140 690
rect 5210 680 5400 690
rect 5410 680 5490 690
rect 5690 680 5700 690
rect 6340 680 6460 690
rect 7420 680 7980 690
rect 9090 680 9100 690
rect 9110 680 9210 690
rect 9330 680 9350 690
rect 0 670 30 680
rect 920 670 1000 680
rect 1360 670 2090 680
rect 2370 670 3320 680
rect 4930 670 5110 680
rect 5120 670 5150 680
rect 5210 670 5400 680
rect 5420 670 5500 680
rect 5690 670 5700 680
rect 6340 670 6470 680
rect 7420 670 7990 680
rect 9090 670 9210 680
rect 9320 670 9330 680
rect 0 660 10 670
rect 950 660 970 670
rect 1350 660 2090 670
rect 2350 660 3300 670
rect 4720 660 4740 670
rect 4930 660 5140 670
rect 5150 660 5160 670
rect 5180 660 5190 670
rect 5210 660 5330 670
rect 5340 660 5400 670
rect 5430 660 5510 670
rect 5690 660 5700 670
rect 6340 660 6470 670
rect 7420 660 7990 670
rect 9090 660 9210 670
rect 9320 660 9330 670
rect 1340 650 2100 660
rect 2330 650 3270 660
rect 4720 650 4750 660
rect 4930 650 5140 660
rect 5190 650 5200 660
rect 5210 650 5290 660
rect 5330 650 5410 660
rect 5430 650 5520 660
rect 5690 650 5700 660
rect 6340 650 6480 660
rect 7420 650 7990 660
rect 9090 650 9110 660
rect 9310 650 9320 660
rect 1330 640 2100 650
rect 2310 640 3250 650
rect 4720 640 4760 650
rect 4930 640 5160 650
rect 5180 640 5210 650
rect 5220 640 5290 650
rect 5320 640 5360 650
rect 5370 640 5420 650
rect 5440 640 5500 650
rect 5510 640 5530 650
rect 5690 640 5700 650
rect 6340 640 6480 650
rect 7420 640 8000 650
rect 9090 640 9110 650
rect 9310 640 9320 650
rect 1330 630 2110 640
rect 2300 630 3230 640
rect 4720 630 4760 640
rect 4930 630 5280 640
rect 5290 630 5300 640
rect 5320 630 5360 640
rect 5370 630 5400 640
rect 5440 630 5510 640
rect 5520 630 5530 640
rect 5690 630 5700 640
rect 6340 630 6490 640
rect 7420 630 8000 640
rect 9080 630 9110 640
rect 9300 630 9330 640
rect 1330 620 1360 630
rect 1390 620 2110 630
rect 2280 620 3160 630
rect 4720 620 4780 630
rect 4940 620 5280 630
rect 5290 620 5310 630
rect 5320 620 5360 630
rect 5370 620 5400 630
rect 5440 620 5510 630
rect 5520 620 5540 630
rect 5690 620 5700 630
rect 6340 620 6500 630
rect 7420 620 8010 630
rect 9080 620 9100 630
rect 1410 610 2110 620
rect 2270 610 3140 620
rect 4720 610 4770 620
rect 4940 610 5280 620
rect 5290 610 5360 620
rect 5370 610 5420 620
rect 5430 610 5440 620
rect 5450 610 5550 620
rect 5690 610 5700 620
rect 6340 610 6510 620
rect 7420 610 8010 620
rect 9070 610 9100 620
rect 9290 610 9300 620
rect 1420 600 2110 610
rect 2250 600 3140 610
rect 4720 600 4760 610
rect 4940 600 5560 610
rect 5690 600 5700 610
rect 6340 600 6510 610
rect 7420 600 8010 610
rect 9070 600 9100 610
rect 9280 600 9300 610
rect 1430 590 2120 600
rect 2230 590 3120 600
rect 4720 590 4740 600
rect 4940 590 5450 600
rect 5460 590 5570 600
rect 5690 590 5700 600
rect 6340 590 6510 600
rect 7420 590 8020 600
rect 9280 590 9290 600
rect 1430 580 2120 590
rect 2220 580 3050 590
rect 3090 580 3110 590
rect 4720 580 4730 590
rect 4950 580 5240 590
rect 5250 580 5450 590
rect 5460 580 5540 590
rect 5550 580 5580 590
rect 5690 580 5700 590
rect 6340 580 6520 590
rect 7420 580 8030 590
rect 9270 580 9290 590
rect 1440 570 2130 580
rect 2200 570 3040 580
rect 4710 570 4740 580
rect 4950 570 5230 580
rect 5240 570 5250 580
rect 5260 570 5280 580
rect 5290 570 5540 580
rect 5550 570 5580 580
rect 5690 570 5700 580
rect 6340 570 6520 580
rect 7420 570 8040 580
rect 9140 570 9150 580
rect 9260 570 9280 580
rect 1450 560 2130 570
rect 2180 560 3020 570
rect 4540 560 4550 570
rect 4710 560 4730 570
rect 4950 560 5250 570
rect 5270 560 5460 570
rect 5470 560 5590 570
rect 5690 560 5700 570
rect 6340 560 6520 570
rect 7420 560 8050 570
rect 9140 560 9160 570
rect 9260 560 9280 570
rect 1460 550 2140 560
rect 2170 550 3010 560
rect 4530 550 4540 560
rect 4710 550 4730 560
rect 4950 550 5470 560
rect 5480 550 5570 560
rect 5580 550 5600 560
rect 5690 550 5700 560
rect 6340 550 6530 560
rect 7420 550 8060 560
rect 9140 550 9170 560
rect 9250 550 9280 560
rect 1480 540 2990 550
rect 4510 540 4540 550
rect 4690 540 4730 550
rect 4950 540 5470 550
rect 5480 540 5620 550
rect 5690 540 5700 550
rect 6340 540 6540 550
rect 7420 540 8070 550
rect 9070 540 9080 550
rect 9120 540 9170 550
rect 9250 540 9270 550
rect 1490 530 2970 540
rect 4500 530 4530 540
rect 4690 530 4720 540
rect 4950 530 5430 540
rect 5470 530 5480 540
rect 5490 530 5570 540
rect 5580 530 5620 540
rect 5690 530 5700 540
rect 6340 530 6540 540
rect 7420 530 8080 540
rect 9070 530 9080 540
rect 9100 530 9160 540
rect 9240 530 9260 540
rect 1500 520 2950 530
rect 4480 520 4530 530
rect 4690 520 4720 530
rect 4960 520 5390 530
rect 5400 520 5430 530
rect 5500 520 5590 530
rect 5610 520 5630 530
rect 5680 520 5700 530
rect 6340 520 6550 530
rect 7420 520 8080 530
rect 9090 520 9160 530
rect 9230 520 9250 530
rect 9950 520 9970 530
rect 1500 510 2900 520
rect 4470 510 4530 520
rect 4690 510 4720 520
rect 4960 510 5370 520
rect 5400 510 5420 520
rect 5480 510 5640 520
rect 5680 510 5700 520
rect 6330 510 6560 520
rect 7420 510 8100 520
rect 9090 510 9180 520
rect 9230 510 9250 520
rect 9940 510 9980 520
rect 1520 500 2870 510
rect 4460 500 4530 510
rect 4690 500 4720 510
rect 4960 500 5360 510
rect 5400 500 5420 510
rect 5470 500 5490 510
rect 5500 500 5650 510
rect 5680 500 5700 510
rect 6330 500 6560 510
rect 7420 500 8100 510
rect 9100 500 9130 510
rect 9160 500 9170 510
rect 9220 500 9250 510
rect 9930 500 9990 510
rect 1530 490 2850 500
rect 4430 490 4530 500
rect 4690 490 4720 500
rect 4960 490 5360 500
rect 5400 490 5420 500
rect 5470 490 5490 500
rect 5510 490 5630 500
rect 5640 490 5660 500
rect 5670 490 5700 500
rect 6330 490 6570 500
rect 7420 490 8110 500
rect 9030 490 9050 500
rect 9080 490 9130 500
rect 9220 490 9250 500
rect 9930 490 9940 500
rect 810 480 830 490
rect 1530 480 2820 490
rect 4400 480 4530 490
rect 4690 480 4720 490
rect 4970 480 5360 490
rect 5390 480 5420 490
rect 5460 480 5630 490
rect 5640 480 5700 490
rect 6330 480 6570 490
rect 7410 480 8120 490
rect 9030 480 9060 490
rect 9080 480 9120 490
rect 9210 480 9240 490
rect 690 470 770 480
rect 790 470 820 480
rect 1540 470 2780 480
rect 4380 470 4450 480
rect 4490 470 4530 480
rect 4690 470 4720 480
rect 4960 470 5360 480
rect 5380 470 5430 480
rect 5450 470 5700 480
rect 6320 470 6570 480
rect 7420 470 8160 480
rect 9210 470 9230 480
rect 9860 470 9870 480
rect 680 460 820 470
rect 1540 460 2110 470
rect 2160 460 2750 470
rect 4280 460 4290 470
rect 4330 460 4440 470
rect 4490 460 4530 470
rect 4690 460 4710 470
rect 4970 460 5610 470
rect 5620 460 5700 470
rect 6320 460 6580 470
rect 7420 460 8170 470
rect 9200 460 9230 470
rect 680 450 810 460
rect 1550 450 2070 460
rect 2200 450 2700 460
rect 4290 450 4440 460
rect 4500 450 4530 460
rect 4690 450 4700 460
rect 4970 450 5260 460
rect 5270 450 5700 460
rect 6330 450 6590 460
rect 7410 450 8180 460
rect 9010 450 9040 460
rect 9200 450 9230 460
rect 680 440 800 450
rect 1550 440 2010 450
rect 2260 440 2660 450
rect 4310 440 4430 450
rect 4510 440 4540 450
rect 4690 440 4700 450
rect 4970 440 5230 450
rect 5240 440 5250 450
rect 5270 440 5710 450
rect 6330 440 6600 450
rect 7410 440 8210 450
rect 9030 440 9040 450
rect 9190 440 9220 450
rect 390 430 400 440
rect 680 430 790 440
rect 1550 430 1850 440
rect 1870 430 1970 440
rect 2290 430 2630 440
rect 4320 430 4430 440
rect 4510 430 4540 440
rect 4690 430 4700 440
rect 4970 430 5230 440
rect 5240 430 5260 440
rect 5270 430 5710 440
rect 6340 430 6600 440
rect 7410 430 8230 440
rect 9190 430 9210 440
rect 400 420 410 430
rect 680 420 780 430
rect 1720 420 1810 430
rect 2320 420 2580 430
rect 4320 420 4430 430
rect 4510 420 4550 430
rect 4690 420 4700 430
rect 4970 420 5230 430
rect 5240 420 5260 430
rect 5270 420 5300 430
rect 5310 420 5710 430
rect 6340 420 6610 430
rect 7420 420 8250 430
rect 9180 420 9210 430
rect 400 410 420 420
rect 680 410 770 420
rect 2370 410 2520 420
rect 4310 410 4340 420
rect 4370 410 4430 420
rect 4510 410 4550 420
rect 4690 410 4710 420
rect 4970 410 5150 420
rect 5160 410 5230 420
rect 5240 410 5250 420
rect 5270 410 5340 420
rect 5360 410 5710 420
rect 6340 410 6620 420
rect 7420 410 8260 420
rect 9100 410 9120 420
rect 9170 410 9200 420
rect 410 400 420 410
rect 680 400 770 410
rect 4310 400 4320 410
rect 4380 400 4420 410
rect 4510 400 4550 410
rect 4680 400 4700 410
rect 4970 400 5150 410
rect 5160 400 5220 410
rect 5240 400 5250 410
rect 5270 400 5340 410
rect 5360 400 5720 410
rect 6340 400 6620 410
rect 7420 400 8270 410
rect 9170 400 9200 410
rect 410 390 420 400
rect 680 390 770 400
rect 4300 390 4310 400
rect 4380 390 4430 400
rect 4500 390 4550 400
rect 4680 390 4710 400
rect 4970 390 5150 400
rect 5160 390 5220 400
rect 5270 390 5340 400
rect 5360 390 5730 400
rect 6340 390 6620 400
rect 7420 390 8290 400
rect 9070 390 9080 400
rect 9160 390 9190 400
rect 420 380 430 390
rect 680 380 770 390
rect 4290 380 4300 390
rect 4390 380 4430 390
rect 4490 380 4550 390
rect 4680 380 4710 390
rect 4980 380 5210 390
rect 5270 380 5330 390
rect 5360 380 5750 390
rect 6340 380 6640 390
rect 7420 380 8280 390
rect 9070 380 9090 390
rect 9160 380 9180 390
rect 420 370 430 380
rect 680 370 780 380
rect 4280 370 4290 380
rect 4400 370 4550 380
rect 4670 370 4710 380
rect 4980 370 5210 380
rect 5240 370 5250 380
rect 5260 370 5330 380
rect 5380 370 5760 380
rect 6350 370 6650 380
rect 7420 370 8290 380
rect 9070 370 9090 380
rect 9150 370 9180 380
rect 420 360 440 370
rect 680 360 800 370
rect 810 360 920 370
rect 4270 360 4280 370
rect 4420 360 4550 370
rect 4690 360 4700 370
rect 4980 360 5210 370
rect 5250 360 5320 370
rect 5380 360 5660 370
rect 5670 360 5770 370
rect 6340 360 6650 370
rect 7420 360 8300 370
rect 9150 360 9170 370
rect 420 350 440 360
rect 680 350 950 360
rect 4470 350 4500 360
rect 4540 350 4550 360
rect 4980 350 5210 360
rect 5250 350 5330 360
rect 5370 350 5780 360
rect 6340 350 6670 360
rect 7420 350 8310 360
rect 9140 350 9160 360
rect 420 340 440 350
rect 680 340 1010 350
rect 4480 340 4490 350
rect 4980 340 5120 350
rect 5130 340 5210 350
rect 5250 340 5330 350
rect 5370 340 5670 350
rect 5680 340 5740 350
rect 5760 340 5790 350
rect 6340 340 6680 350
rect 7420 340 8320 350
rect 9030 340 9040 350
rect 9140 340 9160 350
rect 9240 340 9260 350
rect 9380 340 9420 350
rect 430 330 440 340
rect 720 330 1030 340
rect 4980 330 5110 340
rect 5140 330 5210 340
rect 5220 330 5230 340
rect 5240 330 5340 340
rect 5360 330 5670 340
rect 5680 330 5730 340
rect 5770 330 5810 340
rect 6340 330 6680 340
rect 7420 330 8320 340
rect 9040 330 9090 340
rect 9130 330 9150 340
rect 9240 330 9250 340
rect 9320 330 9350 340
rect 9380 330 9410 340
rect 430 320 440 330
rect 780 320 1040 330
rect 4980 320 5110 330
rect 5130 320 5200 330
rect 5220 320 5670 330
rect 5690 320 5720 330
rect 5790 320 5820 330
rect 6340 320 6690 330
rect 7420 320 8330 330
rect 9040 320 9090 330
rect 9120 320 9140 330
rect 9320 320 9360 330
rect 9390 320 9410 330
rect 430 310 450 320
rect 810 310 1030 320
rect 4620 310 4650 320
rect 4980 310 5200 320
rect 5210 310 5680 320
rect 5690 310 5720 320
rect 5810 310 5840 320
rect 6340 310 6690 320
rect 7410 310 8350 320
rect 9040 310 9080 320
rect 9120 310 9140 320
rect 9300 310 9400 320
rect 440 300 450 310
rect 870 300 880 310
rect 1000 300 1030 310
rect 4570 300 4590 310
rect 4620 300 4650 310
rect 4980 300 5720 310
rect 5830 300 5850 310
rect 6350 300 6700 310
rect 7410 300 8350 310
rect 9110 300 9130 310
rect 9220 300 9250 310
rect 9300 300 9390 310
rect 440 290 450 300
rect 1270 290 1280 300
rect 4580 290 4590 300
rect 4630 290 4650 300
rect 4980 290 5720 300
rect 5840 290 5860 300
rect 6350 290 6700 300
rect 7420 290 8370 300
rect 9100 290 9130 300
rect 9220 290 9270 300
rect 9310 290 9400 300
rect 440 280 450 290
rect 4990 280 5070 290
rect 5080 280 5720 290
rect 5830 280 5880 290
rect 6350 280 6710 290
rect 7420 280 8360 290
rect 8950 280 8970 290
rect 8990 280 9020 290
rect 9100 280 9120 290
rect 9220 280 9280 290
rect 9310 280 9410 290
rect 4990 270 5730 280
rect 5830 270 5900 280
rect 6060 270 6110 280
rect 6360 270 6710 280
rect 7410 270 8370 280
rect 8940 270 9020 280
rect 9090 270 9110 280
rect 9240 270 9290 280
rect 9330 270 9420 280
rect 4990 260 5740 270
rect 5830 260 5920 270
rect 6030 260 6110 270
rect 6360 260 6720 270
rect 7410 260 8380 270
rect 8950 260 9030 270
rect 9090 260 9110 270
rect 9200 260 9230 270
rect 9240 260 9260 270
rect 9340 260 9390 270
rect 9410 260 9420 270
rect 4990 250 5740 260
rect 5810 250 5940 260
rect 6010 250 6100 260
rect 6360 250 6730 260
rect 7410 250 8390 260
rect 8960 250 9040 260
rect 9080 250 9110 260
rect 9200 250 9230 260
rect 4990 240 5710 250
rect 5780 240 6040 250
rect 6070 240 6090 250
rect 6360 240 6740 250
rect 7410 240 8400 250
rect 8970 240 9030 250
rect 9080 240 9100 250
rect 9210 240 9240 250
rect 5000 230 5670 240
rect 5680 230 6010 240
rect 6080 230 6090 240
rect 6360 230 6750 240
rect 7410 230 8400 240
rect 8970 230 9030 240
rect 9070 230 9100 240
rect 5000 220 5940 230
rect 5950 220 5970 230
rect 6040 220 6060 230
rect 6360 220 6750 230
rect 7410 220 8420 230
rect 8970 220 9020 230
rect 9070 220 9090 230
rect 9170 220 9190 230
rect 5000 210 5610 220
rect 5620 210 5720 220
rect 5730 210 5990 220
rect 6030 210 6060 220
rect 6360 210 6760 220
rect 7410 210 8430 220
rect 8970 210 9020 220
rect 9060 210 9080 220
rect 5000 200 5720 210
rect 5740 200 6000 210
rect 6010 200 6020 210
rect 6030 200 6060 210
rect 6370 200 6780 210
rect 7410 200 8440 210
rect 8970 200 9010 210
rect 9050 200 9080 210
rect 9830 200 9840 210
rect 180 190 200 200
rect 5000 190 5720 200
rect 5750 190 6020 200
rect 6030 190 6040 200
rect 6370 190 6790 200
rect 7400 190 8450 200
rect 8950 190 9010 200
rect 9050 190 9070 200
rect 9150 190 9160 200
rect 9810 190 9820 200
rect 160 180 210 190
rect 400 180 420 190
rect 5010 180 5450 190
rect 5490 180 5610 190
rect 5620 180 5720 190
rect 5740 180 5970 190
rect 5980 180 6000 190
rect 6010 180 6020 190
rect 6030 180 6040 190
rect 6370 180 6790 190
rect 7410 180 8460 190
rect 8930 180 9000 190
rect 9040 180 9070 190
rect 9140 180 9170 190
rect 9250 180 9260 190
rect 9270 180 9290 190
rect 9800 180 9820 190
rect 9920 180 9940 190
rect 9980 180 9990 190
rect 180 170 210 180
rect 400 170 420 180
rect 5010 170 5370 180
rect 5420 170 5450 180
rect 5540 170 5580 180
rect 5590 170 5690 180
rect 5700 170 5970 180
rect 5980 170 6000 180
rect 6010 170 6020 180
rect 6380 170 6800 180
rect 7400 170 8460 180
rect 8910 170 9000 180
rect 9040 170 9070 180
rect 9140 170 9160 180
rect 9220 170 9320 180
rect 9790 170 9830 180
rect 9860 170 9890 180
rect 9980 170 9990 180
rect 400 160 430 170
rect 5010 160 5350 170
rect 5660 160 5930 170
rect 5980 160 6000 170
rect 6390 160 6800 170
rect 7400 160 8480 170
rect 8910 160 9000 170
rect 9030 160 9070 170
rect 9140 160 9150 170
rect 9200 160 9320 170
rect 9750 160 9760 170
rect 9780 160 9830 170
rect 9850 160 9890 170
rect 9900 160 9920 170
rect 400 150 430 160
rect 5010 150 5360 160
rect 5700 150 5950 160
rect 5980 150 6000 160
rect 6390 150 6810 160
rect 7400 150 8490 160
rect 8900 150 9010 160
rect 9020 150 9070 160
rect 9210 150 9330 160
rect 9720 150 9740 160
rect 9750 150 9760 160
rect 9790 150 9880 160
rect 9890 150 9930 160
rect 390 140 450 150
rect 5020 140 5340 150
rect 5720 140 5970 150
rect 5980 140 5990 150
rect 6400 140 6810 150
rect 7400 140 8500 150
rect 8910 140 9080 150
rect 9170 140 9180 150
rect 9220 140 9310 150
rect 9320 140 9340 150
rect 9720 140 9740 150
rect 9770 140 9820 150
rect 9830 140 9880 150
rect 9890 140 9930 150
rect 390 130 460 140
rect 5020 130 5340 140
rect 5740 130 5970 140
rect 6400 130 6820 140
rect 7390 130 8500 140
rect 8920 130 9080 140
rect 9170 130 9180 140
rect 9220 130 9340 140
rect 9720 130 9750 140
rect 9770 130 9820 140
rect 9830 130 9920 140
rect 390 120 480 130
rect 5020 120 5340 130
rect 5750 120 5770 130
rect 5790 120 5870 130
rect 5880 120 5930 130
rect 6410 120 6820 130
rect 7390 120 8510 130
rect 8940 120 9050 130
rect 9060 120 9100 130
rect 9220 120 9340 130
rect 9730 120 9740 130
rect 9760 120 9860 130
rect 9870 120 9910 130
rect 9940 120 9960 130
rect 220 110 240 120
rect 390 110 500 120
rect 5030 110 5350 120
rect 5750 110 5770 120
rect 6410 110 6820 120
rect 7390 110 8520 120
rect 8960 110 9040 120
rect 9060 110 9090 120
rect 9220 110 9360 120
rect 9750 110 9850 120
rect 9890 110 9920 120
rect 9990 110 9990 120
rect 220 100 250 110
rect 380 100 520 110
rect 5030 100 5350 110
rect 5750 100 5770 110
rect 6420 100 6830 110
rect 7390 100 8540 110
rect 8970 100 9030 110
rect 9070 100 9090 110
rect 9230 100 9370 110
rect 9750 100 9840 110
rect 9890 100 9910 110
rect 9980 100 9990 110
rect 220 90 240 100
rect 380 90 520 100
rect 5030 90 5360 100
rect 5750 90 5770 100
rect 6420 90 6830 100
rect 7390 90 8550 100
rect 8970 90 9050 100
rect 9070 90 9080 100
rect 9250 90 9430 100
rect 9750 90 9850 100
rect 9980 90 9990 100
rect 230 80 250 90
rect 370 80 540 90
rect 5040 80 5290 90
rect 5300 80 5360 90
rect 5750 80 5770 90
rect 6420 80 6840 90
rect 7380 80 8550 90
rect 8980 80 9060 90
rect 9150 80 9170 90
rect 9250 80 9430 90
rect 9570 80 9580 90
rect 9740 80 9870 90
rect 220 70 250 80
rect 360 70 560 80
rect 5040 70 5360 80
rect 5720 70 5790 80
rect 6440 70 6840 80
rect 7380 70 8570 80
rect 8940 70 8950 80
rect 8970 70 9010 80
rect 9030 70 9060 80
rect 9160 70 9170 80
rect 9240 70 9450 80
rect 9580 70 9600 80
rect 9740 70 9870 80
rect 220 60 260 70
rect 360 60 590 70
rect 5050 60 5250 70
rect 5260 60 5370 70
rect 5700 60 5800 70
rect 6430 60 6840 70
rect 7380 60 8580 70
rect 8970 60 9010 70
rect 9160 60 9180 70
rect 9230 60 9470 70
rect 9680 60 9690 70
rect 9750 60 9830 70
rect 9840 60 9880 70
rect 9910 60 9920 70
rect 9970 60 9990 70
rect 220 50 260 60
rect 360 50 620 60
rect 5050 50 5250 60
rect 5260 50 5370 60
rect 5680 50 5810 60
rect 6430 50 6850 60
rect 7370 50 8590 60
rect 8960 50 9010 60
rect 9170 50 9210 60
rect 9230 50 9270 60
rect 9310 50 9480 60
rect 9680 50 9710 60
rect 9750 50 9890 60
rect 9980 50 9990 60
rect 220 40 270 50
rect 350 40 640 50
rect 5050 40 5160 50
rect 5170 40 5320 50
rect 5330 40 5380 50
rect 5670 40 5820 50
rect 6460 40 6850 50
rect 7360 40 8600 50
rect 8960 40 9010 50
rect 9170 40 9260 50
rect 9300 40 9510 50
rect 9540 40 9560 50
rect 9690 40 9700 50
rect 9770 40 9900 50
rect 220 30 270 40
rect 350 30 640 40
rect 5050 30 5380 40
rect 5660 30 5830 40
rect 6460 30 6860 40
rect 7360 30 8610 40
rect 8930 30 9020 40
rect 9170 30 9530 40
rect 9790 30 9920 40
rect 220 20 270 30
rect 350 20 620 30
rect 5060 20 5310 30
rect 5320 20 5390 30
rect 5650 20 5840 30
rect 6470 20 6870 30
rect 7350 20 8580 30
rect 8600 20 8640 30
rect 8660 20 8700 30
rect 8930 20 8990 30
rect 9170 20 9480 30
rect 9790 20 9920 30
rect 220 10 280 20
rect 350 10 620 20
rect 5060 10 5340 20
rect 5350 10 5390 20
rect 5640 10 5850 20
rect 6470 10 6880 20
rect 7350 10 8580 20
rect 8660 10 8700 20
rect 8920 10 9000 20
rect 9190 10 9490 20
rect 9790 10 9940 20
rect 220 0 270 10
rect 350 0 600 10
rect 5060 0 5340 10
rect 5360 0 5400 10
rect 5640 0 5860 10
rect 6490 0 6900 10
rect 7350 0 8580 10
rect 8690 0 8710 10
rect 8910 0 9010 10
rect 9100 0 9110 10
rect 9190 0 9480 10
rect 9790 0 9940 10
<< metal1 >>
rect 2190 7490 2270 7500
rect 3680 7490 3740 7500
rect 9810 7490 9990 7500
rect 2180 7480 2250 7490
rect 2260 7480 2270 7490
rect 3330 7480 3340 7490
rect 3560 7480 3570 7490
rect 3680 7480 3750 7490
rect 9810 7480 9920 7490
rect 9960 7480 9990 7490
rect 2170 7470 2220 7480
rect 3560 7470 3570 7480
rect 9800 7470 9840 7480
rect 9940 7470 9990 7480
rect 2170 7460 2220 7470
rect 3560 7460 3570 7470
rect 3660 7460 3670 7470
rect 9800 7460 9820 7470
rect 9850 7460 9860 7470
rect 9930 7460 9990 7470
rect 2160 7450 2210 7460
rect 3560 7450 3580 7460
rect 9800 7450 9820 7460
rect 9860 7450 9870 7460
rect 9920 7450 9990 7460
rect 2160 7440 2190 7450
rect 3570 7440 3580 7450
rect 9780 7440 9810 7450
rect 9920 7440 9970 7450
rect 2150 7430 2190 7440
rect 3570 7430 3600 7440
rect 9770 7430 9790 7440
rect 9910 7430 9970 7440
rect 2140 7420 2170 7430
rect 3640 7420 3660 7430
rect 9750 7420 9770 7430
rect 9910 7420 9950 7430
rect 2120 7410 2150 7420
rect 3580 7410 3590 7420
rect 9690 7410 9750 7420
rect 9890 7410 9940 7420
rect 2110 7400 2140 7410
rect 3620 7400 3630 7410
rect 9670 7400 9710 7410
rect 9890 7400 9930 7410
rect 2110 7390 2140 7400
rect 3610 7390 3640 7400
rect 9650 7390 9690 7400
rect 9860 7390 9930 7400
rect 2100 7380 2130 7390
rect 2140 7380 2150 7390
rect 3330 7380 3340 7390
rect 3630 7380 3640 7390
rect 9640 7380 9670 7390
rect 9710 7380 9750 7390
rect 9800 7380 9940 7390
rect 9970 7380 9990 7390
rect 2080 7370 2130 7380
rect 9640 7370 9650 7380
rect 9690 7370 9990 7380
rect 2080 7360 2110 7370
rect 9640 7360 9650 7370
rect 9680 7360 9990 7370
rect 2060 7350 2110 7360
rect 3340 7350 3350 7360
rect 9640 7350 9650 7360
rect 9670 7350 9990 7360
rect 2070 7340 2090 7350
rect 3350 7340 3360 7350
rect 9640 7340 9650 7350
rect 9670 7340 9990 7350
rect 2060 7330 2080 7340
rect 3340 7330 3360 7340
rect 9640 7330 9650 7340
rect 9670 7330 9790 7340
rect 9800 7330 9850 7340
rect 9870 7330 9880 7340
rect 9890 7330 9980 7340
rect 2060 7320 2080 7330
rect 3340 7320 3360 7330
rect 9640 7320 9770 7330
rect 9780 7320 9790 7330
rect 9800 7320 9850 7330
rect 9880 7320 9980 7330
rect 2050 7310 2080 7320
rect 3340 7310 3360 7320
rect 9650 7310 9770 7320
rect 9800 7310 9850 7320
rect 9880 7310 9960 7320
rect 2040 7300 2070 7310
rect 2080 7300 2090 7310
rect 3330 7300 3360 7310
rect 9660 7300 9700 7310
rect 9730 7300 9850 7310
rect 9880 7300 9940 7310
rect 2040 7290 2070 7300
rect 2530 7290 2540 7300
rect 3350 7290 3360 7300
rect 3400 7290 3410 7300
rect 9670 7290 9690 7300
rect 9740 7290 9780 7300
rect 9840 7290 9850 7300
rect 9880 7290 9980 7300
rect 2020 7280 2060 7290
rect 2530 7280 2550 7290
rect 3330 7280 3360 7290
rect 3400 7280 3420 7290
rect 3830 7280 3860 7290
rect 9670 7280 9690 7290
rect 9880 7280 9980 7290
rect 2020 7270 2050 7280
rect 2380 7270 2390 7280
rect 2520 7270 2590 7280
rect 3340 7270 3370 7280
rect 3400 7270 3430 7280
rect 3830 7270 3860 7280
rect 9880 7270 9970 7280
rect 2020 7260 2050 7270
rect 2520 7260 2570 7270
rect 3320 7260 3360 7270
rect 3410 7260 3430 7270
rect 3830 7260 3840 7270
rect 3850 7260 3860 7270
rect 9880 7260 9970 7270
rect 2010 7250 2050 7260
rect 2510 7250 2560 7260
rect 3320 7250 3330 7260
rect 3340 7250 3370 7260
rect 3410 7250 3440 7260
rect 3830 7250 3860 7260
rect 9880 7250 9960 7260
rect 2000 7240 2030 7250
rect 2340 7240 2350 7250
rect 2440 7240 2460 7250
rect 2500 7240 2570 7250
rect 3330 7240 3370 7250
rect 3410 7240 3440 7250
rect 3830 7240 3870 7250
rect 9880 7240 9950 7250
rect 2000 7230 2020 7240
rect 2320 7230 2330 7240
rect 2430 7230 2460 7240
rect 2500 7230 2540 7240
rect 3350 7230 3380 7240
rect 3420 7230 3440 7240
rect 3830 7230 3860 7240
rect 9850 7230 9860 7240
rect 9880 7230 9950 7240
rect 1990 7220 2030 7230
rect 2320 7220 2330 7230
rect 2410 7220 2460 7230
rect 2490 7220 2500 7230
rect 2510 7220 2530 7230
rect 3350 7220 3370 7230
rect 3420 7220 3440 7230
rect 3830 7220 3850 7230
rect 9850 7220 9950 7230
rect 1980 7210 2020 7220
rect 2410 7210 2450 7220
rect 2490 7210 2500 7220
rect 3350 7210 3360 7220
rect 3420 7210 3440 7220
rect 3830 7210 3880 7220
rect 9840 7210 9950 7220
rect 1980 7200 2020 7210
rect 2190 7200 2200 7210
rect 2210 7200 2220 7210
rect 2260 7200 2270 7210
rect 2400 7200 2440 7210
rect 3340 7200 3360 7210
rect 3370 7200 3400 7210
rect 3440 7200 3450 7210
rect 3830 7200 3870 7210
rect 9830 7200 9860 7210
rect 9880 7200 9960 7210
rect 1980 7190 2010 7200
rect 2140 7190 2170 7200
rect 2190 7190 2200 7200
rect 2220 7190 2230 7200
rect 2240 7190 2250 7200
rect 2260 7190 2270 7200
rect 2290 7190 2300 7200
rect 2330 7190 2420 7200
rect 3310 7190 3400 7200
rect 3430 7190 3440 7200
rect 3830 7190 3870 7200
rect 9830 7190 9850 7200
rect 9890 7190 9970 7200
rect 1960 7180 1970 7190
rect 1980 7180 2000 7190
rect 2130 7180 2210 7190
rect 2220 7180 2300 7190
rect 2310 7180 2340 7190
rect 2370 7180 2390 7190
rect 3340 7180 3400 7190
rect 3830 7180 3860 7190
rect 9830 7180 9850 7190
rect 9890 7180 9970 7190
rect 1970 7170 2000 7180
rect 2110 7170 2120 7180
rect 2130 7170 2330 7180
rect 3350 7170 3410 7180
rect 3830 7170 3880 7180
rect 9830 7170 9850 7180
rect 9900 7170 9970 7180
rect 9990 7170 9990 7180
rect 1960 7160 2000 7170
rect 2110 7160 2280 7170
rect 2290 7160 2320 7170
rect 3830 7160 3880 7170
rect 9700 7160 9710 7170
rect 9830 7160 9970 7170
rect 9980 7160 9990 7170
rect 1950 7150 1990 7160
rect 2100 7150 2260 7160
rect 2270 7150 2280 7160
rect 3850 7150 3880 7160
rect 9690 7150 9710 7160
rect 9820 7150 9860 7160
rect 9870 7150 9970 7160
rect 9980 7150 9990 7160
rect 1950 7140 1980 7150
rect 2090 7140 2260 7150
rect 3500 7140 3530 7150
rect 3690 7140 3700 7150
rect 3830 7140 3880 7150
rect 9700 7140 9720 7150
rect 9820 7140 9880 7150
rect 9900 7140 9970 7150
rect 9990 7140 9990 7150
rect 1950 7130 1990 7140
rect 2080 7130 2150 7140
rect 2160 7130 2230 7140
rect 3370 7130 3400 7140
rect 3510 7130 3540 7140
rect 3670 7130 3700 7140
rect 3840 7130 3880 7140
rect 9700 7130 9720 7140
rect 9820 7130 9860 7140
rect 9920 7130 9970 7140
rect 9990 7130 9990 7140
rect 1940 7120 1980 7130
rect 2060 7120 2140 7130
rect 2150 7120 2210 7130
rect 3510 7120 3550 7130
rect 3660 7120 3700 7130
rect 3780 7120 3790 7130
rect 3840 7120 3870 7130
rect 9680 7120 9730 7130
rect 9820 7120 9860 7130
rect 9920 7120 9970 7130
rect 9990 7120 9990 7130
rect 1930 7110 1980 7120
rect 2040 7110 2140 7120
rect 2160 7110 2200 7120
rect 3520 7110 3550 7120
rect 3660 7110 3710 7120
rect 3830 7110 3870 7120
rect 9660 7110 9730 7120
rect 9820 7110 9850 7120
rect 9930 7110 9970 7120
rect 9990 7110 9990 7120
rect 1930 7100 1990 7110
rect 2030 7100 2120 7110
rect 2150 7100 2160 7110
rect 3420 7100 3470 7110
rect 3530 7100 3560 7110
rect 3630 7100 3730 7110
rect 3830 7100 3870 7110
rect 9670 7100 9730 7110
rect 9810 7100 9850 7110
rect 9940 7100 9990 7110
rect 1930 7090 2000 7100
rect 2020 7090 2040 7100
rect 2060 7090 2080 7100
rect 2090 7090 2110 7100
rect 2130 7090 2140 7100
rect 2260 7090 2280 7100
rect 3420 7090 3480 7100
rect 3530 7090 3560 7100
rect 3630 7090 3700 7100
rect 3830 7090 3870 7100
rect 9670 7090 9740 7100
rect 9800 7090 9840 7100
rect 9950 7090 9990 7100
rect 1930 7080 1990 7090
rect 2020 7080 2060 7090
rect 2120 7080 2140 7090
rect 3410 7080 3490 7090
rect 3540 7080 3550 7090
rect 3630 7080 3700 7090
rect 3730 7080 3750 7090
rect 3840 7080 3860 7090
rect 9590 7080 9620 7090
rect 9670 7080 9740 7090
rect 9800 7080 9840 7090
rect 9960 7080 9980 7090
rect 1930 7070 2050 7080
rect 2110 7070 2130 7080
rect 2170 7070 2180 7080
rect 3440 7070 3500 7080
rect 3550 7070 3560 7080
rect 3630 7070 3690 7080
rect 3740 7070 3770 7080
rect 3830 7070 3870 7080
rect 9580 7070 9620 7080
rect 9680 7070 9740 7080
rect 9780 7070 9830 7080
rect 1930 7060 2010 7070
rect 2020 7060 2030 7070
rect 2170 7060 2190 7070
rect 3390 7060 3400 7070
rect 3430 7060 3510 7070
rect 3560 7060 3580 7070
rect 3630 7060 3690 7070
rect 3750 7060 3780 7070
rect 3850 7060 3860 7070
rect 9570 7060 9610 7070
rect 9680 7060 9750 7070
rect 9770 7060 9830 7070
rect 1930 7050 2010 7060
rect 2090 7050 2100 7060
rect 2290 7050 2360 7060
rect 3440 7050 3520 7060
rect 3630 7050 3690 7060
rect 3750 7050 3770 7060
rect 3850 7050 3860 7060
rect 9580 7050 9600 7060
rect 9680 7050 9810 7060
rect 9980 7050 9990 7060
rect 1930 7040 1950 7050
rect 1980 7040 2010 7050
rect 2070 7040 2090 7050
rect 2240 7040 2260 7050
rect 2290 7040 2380 7050
rect 2520 7040 2540 7050
rect 2560 7040 2810 7050
rect 2840 7040 2850 7050
rect 3440 7040 3470 7050
rect 3480 7040 3510 7050
rect 3520 7040 3530 7050
rect 3630 7040 3690 7050
rect 9680 7040 9800 7050
rect 9950 7040 9990 7050
rect 1930 7030 1940 7040
rect 1980 7030 2020 7040
rect 2220 7030 2260 7040
rect 2300 7030 2340 7040
rect 2350 7030 2360 7040
rect 2370 7030 2410 7040
rect 2450 7030 2480 7040
rect 2490 7030 3030 7040
rect 3170 7030 3180 7040
rect 3470 7030 3490 7040
rect 3500 7030 3550 7040
rect 3650 7030 3700 7040
rect 9670 7030 9790 7040
rect 9930 7030 9990 7040
rect 1960 7020 2000 7030
rect 2060 7020 2070 7030
rect 2200 7020 2240 7030
rect 2410 7020 2420 7030
rect 2450 7020 3010 7030
rect 3070 7020 3090 7030
rect 3480 7020 3570 7030
rect 3640 7020 3700 7030
rect 9670 7020 9780 7030
rect 9920 7020 9990 7030
rect 1950 7010 2000 7020
rect 2200 7010 2260 7020
rect 2420 7010 2880 7020
rect 2900 7010 2980 7020
rect 3120 7010 3130 7020
rect 3470 7010 3580 7020
rect 3650 7010 3700 7020
rect 9670 7010 9770 7020
rect 9910 7010 9990 7020
rect 1950 7000 1970 7010
rect 2020 7000 2050 7010
rect 2180 7000 2260 7010
rect 2440 7000 2560 7010
rect 2580 7000 2720 7010
rect 2730 7000 2780 7010
rect 2800 7000 2820 7010
rect 2930 7000 2980 7010
rect 3170 7000 3180 7010
rect 3470 7000 3600 7010
rect 3660 7000 3710 7010
rect 9670 7000 9720 7010
rect 9840 7000 9860 7010
rect 9890 7000 9980 7010
rect 2030 6990 2040 7000
rect 2170 6990 2260 7000
rect 2450 6990 2500 7000
rect 2510 6990 2560 7000
rect 2590 6990 2640 7000
rect 2660 6990 2720 7000
rect 2750 6990 2780 7000
rect 3200 6990 3210 7000
rect 3480 6990 3610 7000
rect 3680 6990 3720 7000
rect 9670 6990 9690 7000
rect 9810 6990 9920 7000
rect 9960 6990 9970 7000
rect 2000 6980 2010 6990
rect 2180 6980 2270 6990
rect 2470 6980 2510 6990
rect 2520 6980 2580 6990
rect 2610 6980 2640 6990
rect 2690 6980 2720 6990
rect 2970 6980 2980 6990
rect 3490 6980 3630 6990
rect 9780 6980 9880 6990
rect 2180 6970 2280 6980
rect 2490 6970 2520 6980
rect 2540 6970 2580 6980
rect 2630 6970 2660 6980
rect 3270 6970 3280 6980
rect 3500 6970 3640 6980
rect 9760 6970 9770 6980
rect 9780 6970 9870 6980
rect 1980 6960 1990 6970
rect 2180 6960 2270 6970
rect 2490 6960 2530 6970
rect 2560 6960 2600 6970
rect 2640 6960 2660 6970
rect 3510 6960 3660 6970
rect 9660 6960 9670 6970
rect 9740 6960 9750 6970
rect 9780 6960 9790 6970
rect 9800 6960 9810 6970
rect 9820 6960 9860 6970
rect 1950 6950 1990 6960
rect 2190 6950 2300 6960
rect 2500 6950 2540 6960
rect 2580 6950 2610 6960
rect 3320 6950 3330 6960
rect 3520 6950 3680 6960
rect 9650 6950 9660 6960
rect 9720 6950 9740 6960
rect 9790 6950 9850 6960
rect 2190 6940 2310 6950
rect 2520 6940 2560 6950
rect 2600 6940 2610 6950
rect 3350 6940 3360 6950
rect 3530 6940 3720 6950
rect 9650 6940 9660 6950
rect 9710 6940 9720 6950
rect 9770 6940 9840 6950
rect 1940 6930 1950 6940
rect 2200 6930 2310 6940
rect 2540 6930 2580 6940
rect 2700 6930 2710 6940
rect 3550 6930 3730 6940
rect 9650 6930 9660 6940
rect 9680 6930 9710 6940
rect 9750 6930 9840 6940
rect 1930 6920 1940 6930
rect 2210 6920 2330 6930
rect 2550 6920 2580 6930
rect 2720 6920 2730 6930
rect 3400 6920 3410 6930
rect 3560 6920 3740 6930
rect 9650 6920 9660 6930
rect 9680 6920 9690 6930
rect 9700 6920 9840 6930
rect 1920 6910 1930 6920
rect 2220 6910 2360 6920
rect 2580 6910 2590 6920
rect 3590 6910 3740 6920
rect 9650 6910 9680 6920
rect 9700 6910 9840 6920
rect 1900 6900 1910 6910
rect 2230 6900 2360 6910
rect 2680 6900 2690 6910
rect 3520 6900 3530 6910
rect 3600 6900 3760 6910
rect 9680 6900 9850 6910
rect 1890 6890 1900 6900
rect 2250 6890 2380 6900
rect 2700 6890 2710 6900
rect 3470 6890 3480 6900
rect 3530 6890 3540 6900
rect 3620 6890 3770 6900
rect 9680 6890 9850 6900
rect 1890 6880 1900 6890
rect 2260 6880 2410 6890
rect 3490 6880 3500 6890
rect 3630 6880 3780 6890
rect 9680 6880 9850 6890
rect 2260 6870 2420 6880
rect 3510 6870 3520 6880
rect 3570 6870 3580 6880
rect 3650 6870 3780 6880
rect 9680 6870 9860 6880
rect 1920 6860 1940 6870
rect 2280 6860 2440 6870
rect 3530 6860 3540 6870
rect 3580 6860 3600 6870
rect 3670 6860 3790 6870
rect 9680 6860 9860 6870
rect 9950 6860 9980 6870
rect 2290 6850 2470 6860
rect 2720 6850 2730 6860
rect 3550 6850 3560 6860
rect 3680 6850 3810 6860
rect 9680 6850 9860 6860
rect 9940 6850 9990 6860
rect 1890 6840 1900 6850
rect 2300 6840 2490 6850
rect 3610 6840 3630 6850
rect 3690 6840 3820 6850
rect 9680 6840 9870 6850
rect 9920 6840 9990 6850
rect 2330 6830 2500 6840
rect 3700 6830 3820 6840
rect 9680 6830 9870 6840
rect 9930 6830 9990 6840
rect 1890 6820 1900 6830
rect 2350 6820 2510 6830
rect 3650 6820 3660 6830
rect 3710 6820 3830 6830
rect 9680 6820 9860 6830
rect 9910 6820 9990 6830
rect 1890 6810 1900 6820
rect 2370 6810 2550 6820
rect 3620 6810 3630 6820
rect 3670 6810 3680 6820
rect 3730 6810 3830 6820
rect 9630 6810 9640 6820
rect 9680 6810 9860 6820
rect 9920 6810 9990 6820
rect 1860 6800 1890 6810
rect 1950 6800 1970 6810
rect 2390 6800 2560 6810
rect 2570 6800 2580 6810
rect 3740 6800 3830 6810
rect 9680 6800 9870 6810
rect 9920 6800 9990 6810
rect 1880 6790 1900 6800
rect 1940 6790 1960 6800
rect 1980 6790 2020 6800
rect 2290 6790 2360 6800
rect 2410 6790 2680 6800
rect 3650 6790 3660 6800
rect 3680 6790 3710 6800
rect 3760 6790 3840 6800
rect 9620 6790 9640 6800
rect 9680 6790 9860 6800
rect 9920 6790 9990 6800
rect 1890 6780 1900 6790
rect 1920 6780 1940 6790
rect 1960 6780 1970 6790
rect 2010 6780 2030 6790
rect 2270 6780 2370 6790
rect 2460 6780 2710 6790
rect 3770 6780 3850 6790
rect 9610 6780 9650 6790
rect 9680 6780 9860 6790
rect 9930 6780 9990 6790
rect 1890 6770 1910 6780
rect 1960 6770 1970 6780
rect 2000 6770 2040 6780
rect 2260 6770 2300 6780
rect 2380 6770 2390 6780
rect 2500 6770 2730 6780
rect 2750 6770 2800 6780
rect 3680 6770 3690 6780
rect 3710 6770 3720 6780
rect 3780 6770 3850 6780
rect 9600 6770 9650 6780
rect 9680 6770 9860 6780
rect 9940 6770 9990 6780
rect 1890 6760 1910 6770
rect 1990 6760 2040 6770
rect 2250 6760 2290 6770
rect 2400 6760 2410 6770
rect 2530 6760 2570 6770
rect 2650 6760 2860 6770
rect 3720 6760 3740 6770
rect 3790 6760 3850 6770
rect 9600 6760 9640 6770
rect 9690 6760 9850 6770
rect 9950 6760 9990 6770
rect 1880 6750 1900 6760
rect 2030 6750 2060 6760
rect 2260 6750 2280 6760
rect 2420 6750 2430 6760
rect 2730 6750 2920 6760
rect 3710 6750 3720 6760
rect 3740 6750 3750 6760
rect 3800 6750 3850 6760
rect 9560 6750 9570 6760
rect 9600 6750 9640 6760
rect 9690 6750 9840 6760
rect 9960 6750 9990 6760
rect 1880 6740 1910 6750
rect 1940 6740 1950 6750
rect 1980 6740 1990 6750
rect 2250 6740 2260 6750
rect 2440 6740 2450 6750
rect 2820 6740 3030 6750
rect 3750 6740 3770 6750
rect 3810 6740 3870 6750
rect 9600 6740 9640 6750
rect 9690 6740 9840 6750
rect 1860 6730 1930 6740
rect 2240 6730 2260 6740
rect 2900 6730 3080 6740
rect 3110 6730 3120 6740
rect 3770 6730 3780 6740
rect 3830 6730 3870 6740
rect 9550 6730 9560 6740
rect 9600 6730 9640 6740
rect 9690 6730 9840 6740
rect 1890 6720 1980 6730
rect 2230 6720 2240 6730
rect 3030 6720 3150 6730
rect 3190 6720 3200 6730
rect 3840 6720 3880 6730
rect 9540 6720 9550 6730
rect 9560 6720 9570 6730
rect 9600 6720 9640 6730
rect 9690 6720 9850 6730
rect 1850 6710 1860 6720
rect 1890 6710 1980 6720
rect 2230 6710 2240 6720
rect 2510 6710 2520 6720
rect 3100 6710 3240 6720
rect 3780 6710 3800 6720
rect 3850 6710 3890 6720
rect 9560 6710 9570 6720
rect 9600 6710 9640 6720
rect 9690 6710 9850 6720
rect 1880 6700 1950 6710
rect 1960 6700 1980 6710
rect 2220 6700 2240 6710
rect 2540 6700 2550 6710
rect 3200 6700 3290 6710
rect 3800 6700 3810 6710
rect 3860 6700 3900 6710
rect 9540 6700 9550 6710
rect 9560 6700 9570 6710
rect 9600 6700 9640 6710
rect 9690 6700 9840 6710
rect 9990 6700 9990 6710
rect 1870 6690 1960 6700
rect 2220 6690 2250 6700
rect 2570 6690 2580 6700
rect 3230 6690 3350 6700
rect 3820 6690 3830 6700
rect 3870 6690 3910 6700
rect 9530 6690 9560 6700
rect 9600 6690 9640 6700
rect 9690 6690 9840 6700
rect 9980 6690 9990 6700
rect 1860 6680 1890 6690
rect 1910 6680 1970 6690
rect 2220 6680 2250 6690
rect 2580 6680 2630 6690
rect 3320 6680 3410 6690
rect 3800 6680 3810 6690
rect 3880 6680 3910 6690
rect 9520 6680 9550 6690
rect 9610 6680 9640 6690
rect 9690 6680 9710 6690
rect 9720 6680 9830 6690
rect 9950 6680 9970 6690
rect 1910 6670 1930 6680
rect 1950 6670 1960 6680
rect 2230 6670 2240 6680
rect 2580 6670 2670 6680
rect 3370 6670 3430 6680
rect 3820 6670 3830 6680
rect 3840 6670 3850 6680
rect 3890 6670 3910 6680
rect 9520 6670 9540 6680
rect 9610 6670 9650 6680
rect 9690 6670 9820 6680
rect 9920 6670 9940 6680
rect 1880 6660 1930 6670
rect 2220 6660 2240 6670
rect 2580 6660 2660 6670
rect 3420 6660 3480 6670
rect 3830 6660 3850 6670
rect 3900 6660 3920 6670
rect 9510 6660 9530 6670
rect 9610 6660 9650 6670
rect 9690 6660 9810 6670
rect 9890 6660 9910 6670
rect 1880 6650 1900 6660
rect 1930 6650 1940 6660
rect 2210 6650 2230 6660
rect 2590 6650 2650 6660
rect 3470 6650 3500 6660
rect 3850 6650 3860 6660
rect 3910 6650 3930 6660
rect 9500 6650 9510 6660
rect 9610 6650 9640 6660
rect 9690 6650 9710 6660
rect 9720 6650 9780 6660
rect 9850 6650 9870 6660
rect 1850 6640 1860 6650
rect 2200 6640 2220 6650
rect 2600 6640 2660 6650
rect 3500 6640 3530 6650
rect 3850 6640 3860 6650
rect 3910 6640 3940 6650
rect 9500 6640 9520 6650
rect 9620 6640 9650 6650
rect 9690 6640 9710 6650
rect 9820 6640 9840 6650
rect 1820 6630 1850 6640
rect 1860 6630 1890 6640
rect 2190 6630 2210 6640
rect 2600 6630 2650 6640
rect 3530 6630 3550 6640
rect 3920 6630 3940 6640
rect 9490 6630 9520 6640
rect 9620 6630 9650 6640
rect 9700 6630 9710 6640
rect 9760 6630 9770 6640
rect 9800 6630 9810 6640
rect 1750 6620 1780 6630
rect 1810 6620 1840 6630
rect 2180 6620 2210 6630
rect 2610 6620 2650 6630
rect 3560 6620 3600 6630
rect 3870 6620 3880 6630
rect 3930 6620 3950 6630
rect 9480 6620 9500 6630
rect 9620 6620 9630 6630
rect 9640 6620 9650 6630
rect 9690 6620 9700 6630
rect 9750 6620 9780 6630
rect 1620 6610 1670 6620
rect 1760 6610 1800 6620
rect 2170 6610 2190 6620
rect 2620 6610 2660 6620
rect 3590 6610 3620 6620
rect 3880 6610 3890 6620
rect 3930 6610 3950 6620
rect 9490 6610 9500 6620
rect 9630 6610 9640 6620
rect 9690 6610 9700 6620
rect 9730 6610 9750 6620
rect 1610 6600 1620 6610
rect 1630 6600 1640 6610
rect 1760 6600 1770 6610
rect 2160 6600 2180 6610
rect 2610 6600 2660 6610
rect 3620 6600 3640 6610
rect 3890 6600 3900 6610
rect 3940 6600 3960 6610
rect 9490 6600 9510 6610
rect 9630 6600 9640 6610
rect 9710 6600 9720 6610
rect 1600 6590 1610 6600
rect 1620 6590 1630 6600
rect 1760 6590 1770 6600
rect 2130 6590 2180 6600
rect 2620 6590 2660 6600
rect 3640 6590 3680 6600
rect 3900 6590 3910 6600
rect 3940 6590 3960 6600
rect 9490 6590 9510 6600
rect 1780 6580 1790 6590
rect 2090 6580 2100 6590
rect 2130 6580 2170 6590
rect 2620 6580 2670 6590
rect 3670 6580 3700 6590
rect 3950 6580 3960 6590
rect 9490 6580 9500 6590
rect 1560 6570 1570 6580
rect 1600 6570 1610 6580
rect 1790 6570 1800 6580
rect 2070 6570 2080 6580
rect 2130 6570 2170 6580
rect 2620 6570 2660 6580
rect 3710 6570 3720 6580
rect 3960 6570 3970 6580
rect 1800 6560 1810 6570
rect 1990 6560 2000 6570
rect 2020 6560 2040 6570
rect 2050 6560 2080 6570
rect 2620 6560 2680 6570
rect 3720 6560 3740 6570
rect 3960 6560 3980 6570
rect 1520 6550 1530 6560
rect 1580 6550 1590 6560
rect 1810 6550 1820 6560
rect 2000 6550 2010 6560
rect 2620 6550 2670 6560
rect 3750 6550 3760 6560
rect 3930 6550 3940 6560
rect 3970 6550 3990 6560
rect 1500 6540 1510 6550
rect 1580 6540 1590 6550
rect 1630 6540 1690 6550
rect 1710 6540 1730 6550
rect 1820 6540 1830 6550
rect 2630 6540 2680 6550
rect 3760 6540 3770 6550
rect 3980 6540 4000 6550
rect 1470 6530 1480 6540
rect 1500 6530 1510 6540
rect 1570 6530 1620 6540
rect 1740 6530 1750 6540
rect 1830 6530 1840 6540
rect 2030 6530 2050 6540
rect 2630 6530 2690 6540
rect 3780 6530 3800 6540
rect 3980 6530 4000 6540
rect 1440 6520 1490 6530
rect 1570 6520 1610 6530
rect 1730 6520 1770 6530
rect 1840 6520 1850 6530
rect 2040 6520 2050 6530
rect 2580 6520 2610 6530
rect 3810 6520 3820 6530
rect 3980 6520 4000 6530
rect 9990 6520 9990 6530
rect 1370 6510 1390 6520
rect 1420 6510 1430 6520
rect 1480 6510 1490 6520
rect 1570 6510 1600 6520
rect 1730 6510 1780 6520
rect 1840 6510 1850 6520
rect 2060 6510 2070 6520
rect 2550 6510 2570 6520
rect 3830 6510 3840 6520
rect 3960 6510 3970 6520
rect 3990 6510 4000 6520
rect 6380 6510 6390 6520
rect 6520 6510 6530 6520
rect 9970 6510 9990 6520
rect 1330 6500 1380 6510
rect 1450 6500 1470 6510
rect 1550 6500 1590 6510
rect 1720 6500 1790 6510
rect 1850 6500 1860 6510
rect 2080 6500 2090 6510
rect 2520 6500 2550 6510
rect 3850 6500 3860 6510
rect 3990 6500 4000 6510
rect 6380 6500 6430 6510
rect 6480 6500 6540 6510
rect 9940 6500 9980 6510
rect 1300 6490 1310 6500
rect 1330 6490 1370 6500
rect 1540 6490 1590 6500
rect 1690 6490 1800 6500
rect 1850 6490 1890 6500
rect 2100 6490 2110 6500
rect 2410 6490 2440 6500
rect 2480 6490 2550 6500
rect 3870 6490 3880 6500
rect 4000 6490 4010 6500
rect 6380 6490 6430 6500
rect 6450 6490 6540 6500
rect 9890 6490 9980 6500
rect 1280 6480 1290 6490
rect 1300 6480 1310 6490
rect 1330 6480 1380 6490
rect 1430 6480 1440 6490
rect 1550 6480 1580 6490
rect 1680 6480 1710 6490
rect 1760 6480 1800 6490
rect 1840 6480 1890 6490
rect 2100 6480 2120 6490
rect 2430 6480 2470 6490
rect 2480 6480 2550 6490
rect 3880 6480 3900 6490
rect 4000 6480 4010 6490
rect 6390 6480 6540 6490
rect 9870 6480 9890 6490
rect 9910 6480 9970 6490
rect 1270 6470 1280 6480
rect 1370 6470 1420 6480
rect 1440 6470 1450 6480
rect 1560 6470 1590 6480
rect 1660 6470 1690 6480
rect 1770 6470 1810 6480
rect 1850 6470 1900 6480
rect 1920 6470 1950 6480
rect 2120 6470 2130 6480
rect 2400 6470 2410 6480
rect 2430 6470 2510 6480
rect 2530 6470 2540 6480
rect 2560 6470 2570 6480
rect 3900 6470 3910 6480
rect 3990 6470 4000 6480
rect 4010 6470 4020 6480
rect 6400 6470 6530 6480
rect 9850 6470 9880 6480
rect 9930 6470 9960 6480
rect 1250 6460 1260 6470
rect 1310 6460 1330 6470
rect 1380 6460 1390 6470
rect 1400 6460 1410 6470
rect 1550 6460 1580 6470
rect 1620 6460 1680 6470
rect 1770 6460 1810 6470
rect 1860 6460 1910 6470
rect 1920 6460 1960 6470
rect 2100 6460 2150 6470
rect 2430 6460 2500 6470
rect 2520 6460 2530 6470
rect 3920 6460 3930 6470
rect 4010 6460 4020 6470
rect 6140 6460 6150 6470
rect 6160 6460 6170 6470
rect 6400 6460 6520 6470
rect 9780 6460 9880 6470
rect 9930 6460 9970 6470
rect 1240 6450 1250 6460
rect 1360 6450 1380 6460
rect 1550 6450 1580 6460
rect 1620 6450 1660 6460
rect 1770 6450 1810 6460
rect 1890 6450 1900 6460
rect 1940 6450 2100 6460
rect 2120 6450 2150 6460
rect 2390 6450 2400 6460
rect 2430 6450 2440 6460
rect 2470 6450 2490 6460
rect 2510 6450 2520 6460
rect 4020 6450 4030 6460
rect 6120 6450 6190 6460
rect 6410 6450 6530 6460
rect 6540 6450 6570 6460
rect 9750 6450 9870 6460
rect 9930 6450 9980 6460
rect 1250 6440 1260 6450
rect 1440 6440 1460 6450
rect 1550 6440 1580 6450
rect 1590 6440 1650 6450
rect 1770 6440 1820 6450
rect 1940 6440 2080 6450
rect 2120 6440 2140 6450
rect 2270 6440 2280 6450
rect 2490 6440 2520 6450
rect 2540 6440 2550 6450
rect 3950 6440 3960 6450
rect 6120 6440 6210 6450
rect 6310 6440 6330 6450
rect 6420 6440 6570 6450
rect 9700 6440 9800 6450
rect 9930 6440 9980 6450
rect 1280 6430 1290 6440
rect 1370 6430 1380 6440
rect 1420 6430 1470 6440
rect 1550 6430 1650 6440
rect 1770 6430 1810 6440
rect 1960 6430 2100 6440
rect 2290 6430 2310 6440
rect 2380 6430 2390 6440
rect 2410 6430 2430 6440
rect 2500 6430 2530 6440
rect 6120 6430 6210 6440
rect 6220 6430 6230 6440
rect 6280 6430 6290 6440
rect 6320 6430 6340 6440
rect 6420 6430 6470 6440
rect 6480 6430 6590 6440
rect 9680 6430 9800 6440
rect 9930 6430 9950 6440
rect 9970 6430 9990 6440
rect 1370 6420 1400 6430
rect 1420 6420 1470 6430
rect 1550 6420 1640 6430
rect 1790 6420 1820 6430
rect 1960 6420 2070 6430
rect 2080 6420 2090 6430
rect 2330 6420 2350 6430
rect 2370 6420 2380 6430
rect 2410 6420 2430 6430
rect 2490 6420 2500 6430
rect 2510 6420 2520 6430
rect 3980 6420 3990 6430
rect 5840 6420 5870 6430
rect 6110 6420 6220 6430
rect 6230 6420 6240 6430
rect 6260 6420 6290 6430
rect 6340 6420 6350 6430
rect 6370 6420 6450 6430
rect 6490 6420 6570 6430
rect 9660 6420 9760 6430
rect 9770 6420 9780 6430
rect 9930 6420 9940 6430
rect 9980 6420 9990 6430
rect 1370 6410 1400 6420
rect 1420 6410 1440 6420
rect 1470 6410 1490 6420
rect 1550 6410 1640 6420
rect 1970 6410 2040 6420
rect 2370 6410 2380 6420
rect 2510 6410 2520 6420
rect 4000 6410 4010 6420
rect 6120 6410 6180 6420
rect 6360 6410 6450 6420
rect 6490 6410 6550 6420
rect 6560 6410 6580 6420
rect 9650 6410 9770 6420
rect 9930 6410 9940 6420
rect 9990 6410 9990 6420
rect 1260 6400 1270 6410
rect 1370 6400 1400 6410
rect 1410 6400 1420 6410
rect 1460 6400 1480 6410
rect 1550 6400 1630 6410
rect 2400 6400 2410 6410
rect 2490 6400 2510 6410
rect 6360 6400 6460 6410
rect 6500 6400 6590 6410
rect 9650 6400 9720 6410
rect 9730 6400 9750 6410
rect 9930 6400 9940 6410
rect 1370 6390 1380 6400
rect 1460 6390 1470 6400
rect 1550 6390 1630 6400
rect 2390 6390 2400 6400
rect 2410 6390 2420 6400
rect 4030 6390 4040 6400
rect 6380 6390 6470 6400
rect 6490 6390 6590 6400
rect 9640 6390 9690 6400
rect 9720 6390 9750 6400
rect 9760 6390 9810 6400
rect 9920 6390 9940 6400
rect 1460 6380 1470 6390
rect 1550 6380 1620 6390
rect 2400 6380 2410 6390
rect 2470 6380 2480 6390
rect 4040 6380 4050 6390
rect 6390 6380 6600 6390
rect 9640 6380 9700 6390
rect 9710 6380 9830 6390
rect 9930 6380 9940 6390
rect 9990 6380 9990 6390
rect 1460 6370 1470 6380
rect 1550 6370 1610 6380
rect 1750 6370 1780 6380
rect 1820 6370 1830 6380
rect 2400 6370 2410 6380
rect 2460 6370 2470 6380
rect 6380 6370 6390 6380
rect 6400 6370 6600 6380
rect 9630 6370 9850 6380
rect 9930 6370 9950 6380
rect 9970 6370 9990 6380
rect 1240 6360 1260 6370
rect 1460 6360 1480 6370
rect 1550 6360 1610 6370
rect 1740 6360 1760 6370
rect 2410 6360 2420 6370
rect 2460 6360 2480 6370
rect 4070 6360 4080 6370
rect 6410 6360 6600 6370
rect 9630 6360 9710 6370
rect 9740 6360 9780 6370
rect 9790 6360 9860 6370
rect 9940 6360 9990 6370
rect 1250 6350 1260 6360
rect 1460 6350 1480 6360
rect 1550 6350 1600 6360
rect 1720 6350 1750 6360
rect 1830 6350 1840 6360
rect 2410 6350 2420 6360
rect 4080 6350 4090 6360
rect 6430 6350 6610 6360
rect 9630 6350 9690 6360
rect 9740 6350 9780 6360
rect 9800 6350 9860 6360
rect 9960 6350 9990 6360
rect 1430 6340 1470 6350
rect 1560 6340 1600 6350
rect 1710 6340 1740 6350
rect 1830 6340 1840 6350
rect 2450 6340 2470 6350
rect 5740 6340 5780 6350
rect 6450 6340 6670 6350
rect 9640 6340 9680 6350
rect 9740 6340 9780 6350
rect 9810 6340 9850 6350
rect 9960 6340 9990 6350
rect 1430 6330 1460 6340
rect 1560 6330 1590 6340
rect 1710 6330 1740 6340
rect 1830 6330 1840 6340
rect 2420 6330 2430 6340
rect 5750 6330 5790 6340
rect 6480 6330 6500 6340
rect 6510 6330 6680 6340
rect 6710 6330 6720 6340
rect 9480 6330 9500 6340
rect 9640 6330 9710 6340
rect 9740 6330 9770 6340
rect 9820 6330 9840 6340
rect 9940 6330 9990 6340
rect 1420 6320 1450 6330
rect 1560 6320 1590 6330
rect 1700 6320 1730 6330
rect 1830 6320 1840 6330
rect 2420 6320 2430 6330
rect 2470 6320 2480 6330
rect 5500 6320 5510 6330
rect 5710 6320 5720 6330
rect 5740 6320 5790 6330
rect 6520 6320 6700 6330
rect 6720 6320 6730 6330
rect 9470 6320 9500 6330
rect 9640 6320 9690 6330
rect 9740 6320 9790 6330
rect 9800 6320 9830 6330
rect 9940 6320 9990 6330
rect 1420 6310 1450 6320
rect 1560 6310 1590 6320
rect 1680 6310 1730 6320
rect 1800 6310 1830 6320
rect 2420 6310 2430 6320
rect 2440 6310 2450 6320
rect 4120 6310 4130 6320
rect 5700 6310 5720 6320
rect 5760 6310 5770 6320
rect 6540 6310 6750 6320
rect 9470 6310 9490 6320
rect 9640 6310 9690 6320
rect 9790 6310 9800 6320
rect 9950 6310 9990 6320
rect 1260 6300 1270 6310
rect 1420 6300 1430 6310
rect 1560 6300 1580 6310
rect 1660 6300 1720 6310
rect 1780 6300 1830 6310
rect 2420 6300 2430 6310
rect 2440 6300 2450 6310
rect 5410 6300 5430 6310
rect 5470 6300 5500 6310
rect 5520 6300 5570 6310
rect 5660 6300 5670 6310
rect 6560 6300 6610 6310
rect 6620 6300 6750 6310
rect 9400 6300 9410 6310
rect 9640 6300 9700 6310
rect 9940 6300 9980 6310
rect 1410 6290 1420 6300
rect 1570 6290 1580 6300
rect 1640 6290 1720 6300
rect 1760 6290 1830 6300
rect 2420 6290 2430 6300
rect 2440 6290 2450 6300
rect 4150 6290 4160 6300
rect 5410 6290 5450 6300
rect 5500 6290 5510 6300
rect 5640 6290 5670 6300
rect 6570 6290 6770 6300
rect 9640 6290 9700 6300
rect 9820 6290 9890 6300
rect 9930 6290 9960 6300
rect 1540 6280 1550 6290
rect 1570 6280 1580 6290
rect 1630 6280 1710 6290
rect 1760 6280 1820 6290
rect 2420 6280 2430 6290
rect 2460 6280 2470 6290
rect 4160 6280 4170 6290
rect 5400 6280 5410 6290
rect 5520 6280 5550 6290
rect 5600 6280 5620 6290
rect 6570 6280 6610 6290
rect 6620 6280 6770 6290
rect 9410 6280 9420 6290
rect 9640 6280 9680 6290
rect 9810 6280 9910 6290
rect 9930 6280 9950 6290
rect 1260 6270 1280 6280
rect 1410 6270 1420 6280
rect 1530 6270 1560 6280
rect 1570 6270 1580 6280
rect 1620 6270 1700 6280
rect 1750 6270 1820 6280
rect 2420 6270 2430 6280
rect 4170 6270 4180 6280
rect 5370 6270 5390 6280
rect 5520 6270 5540 6280
rect 6580 6270 6660 6280
rect 6680 6270 6710 6280
rect 6740 6270 6770 6280
rect 9410 6270 9430 6280
rect 9640 6270 9680 6280
rect 9810 6270 9870 6280
rect 9940 6270 9960 6280
rect 1410 6260 1420 6270
rect 1520 6260 1540 6270
rect 1550 6260 1570 6270
rect 1610 6260 1690 6270
rect 1740 6260 1810 6270
rect 2420 6260 2430 6270
rect 4180 6260 4190 6270
rect 5360 6260 5390 6270
rect 5400 6260 5420 6270
rect 5510 6260 5530 6270
rect 6590 6260 6650 6270
rect 6680 6260 6710 6270
rect 6740 6260 6770 6270
rect 9410 6260 9420 6270
rect 9590 6260 9610 6270
rect 9640 6260 9680 6270
rect 9810 6260 9850 6270
rect 1410 6250 1420 6260
rect 1560 6250 1580 6260
rect 1610 6250 1680 6260
rect 1740 6250 1810 6260
rect 2420 6250 2430 6260
rect 4190 6250 4200 6260
rect 5330 6250 5390 6260
rect 5410 6250 5420 6260
rect 5500 6250 5520 6260
rect 6590 6250 6650 6260
rect 6660 6250 6720 6260
rect 6740 6250 6770 6260
rect 9560 6250 9620 6260
rect 9660 6250 9680 6260
rect 9810 6250 9820 6260
rect 1410 6240 1420 6250
rect 1600 6240 1660 6250
rect 1730 6240 1800 6250
rect 2420 6240 2430 6250
rect 2440 6240 2450 6250
rect 4200 6240 4210 6250
rect 5330 6240 5340 6250
rect 5360 6240 5370 6250
rect 5490 6240 5520 6250
rect 6610 6240 6650 6250
rect 6660 6240 6770 6250
rect 9520 6240 9530 6250
rect 9600 6240 9620 6250
rect 9650 6240 9690 6250
rect 9800 6240 9810 6250
rect 1410 6230 1420 6240
rect 1560 6230 1570 6240
rect 1600 6230 1660 6240
rect 1710 6230 1790 6240
rect 2420 6230 2430 6240
rect 2440 6230 2450 6240
rect 4210 6230 4220 6240
rect 5320 6230 5330 6240
rect 5340 6230 5350 6240
rect 5370 6230 5380 6240
rect 5480 6230 5510 6240
rect 6620 6230 6630 6240
rect 6650 6230 6750 6240
rect 9420 6230 9440 6240
rect 9490 6230 9510 6240
rect 9520 6230 9530 6240
rect 9600 6230 9610 6240
rect 9660 6230 9680 6240
rect 9800 6230 9810 6240
rect 1600 6220 1660 6230
rect 1700 6220 1790 6230
rect 2420 6220 2430 6230
rect 2440 6220 2450 6230
rect 4220 6220 4230 6230
rect 5310 6220 5320 6230
rect 5360 6220 5370 6230
rect 5470 6220 5500 6230
rect 6650 6220 6750 6230
rect 9420 6220 9490 6230
rect 9500 6220 9520 6230
rect 9540 6220 9550 6230
rect 9600 6220 9610 6230
rect 9660 6220 9680 6230
rect 9790 6220 9810 6230
rect 1340 6210 1350 6220
rect 1420 6210 1430 6220
rect 1570 6210 1580 6220
rect 1610 6210 1670 6220
rect 1690 6210 1780 6220
rect 2420 6210 2430 6220
rect 2440 6210 2450 6220
rect 5300 6210 5320 6220
rect 5350 6210 5360 6220
rect 5390 6210 5400 6220
rect 5460 6210 5480 6220
rect 6670 6210 6760 6220
rect 9420 6210 9450 6220
rect 9480 6210 9500 6220
rect 9520 6210 9530 6220
rect 9600 6210 9610 6220
rect 9670 6210 9700 6220
rect 9790 6210 9800 6220
rect 1340 6200 1360 6210
rect 1570 6200 1580 6210
rect 1620 6200 1660 6210
rect 1700 6200 1730 6210
rect 1740 6200 1760 6210
rect 2420 6200 2430 6210
rect 2450 6200 2460 6210
rect 5380 6200 5390 6210
rect 5440 6200 5470 6210
rect 6670 6200 6760 6210
rect 9380 6200 9410 6210
rect 9600 6200 9610 6210
rect 9670 6200 9690 6210
rect 9780 6200 9800 6210
rect 1340 6190 1360 6200
rect 1570 6190 1580 6200
rect 1630 6190 1670 6200
rect 1690 6190 1720 6200
rect 2420 6190 2430 6200
rect 2450 6190 2460 6200
rect 5320 6190 5340 6200
rect 5440 6190 5460 6200
rect 6670 6190 6750 6200
rect 9360 6190 9430 6200
rect 9600 6190 9610 6200
rect 9680 6190 9690 6200
rect 9780 6190 9800 6200
rect 1350 6180 1370 6190
rect 1420 6180 1430 6190
rect 1580 6180 1590 6190
rect 1630 6180 1680 6190
rect 1690 6180 1720 6190
rect 4250 6180 4260 6190
rect 5310 6180 5330 6190
rect 5430 6180 5450 6190
rect 6680 6180 6740 6190
rect 9320 6180 9400 6190
rect 9420 6180 9430 6190
rect 9600 6180 9610 6190
rect 9680 6180 9700 6190
rect 9780 6180 9810 6190
rect 1300 6170 1310 6180
rect 1350 6170 1370 6180
rect 1580 6170 1590 6180
rect 1640 6170 1720 6180
rect 5420 6170 5440 6180
rect 6680 6170 6740 6180
rect 9300 6170 9430 6180
rect 9600 6170 9610 6180
rect 9680 6170 9700 6180
rect 9790 6170 9820 6180
rect 1270 6160 1290 6170
rect 1350 6160 1380 6170
rect 1650 6160 1720 6170
rect 4260 6160 4270 6170
rect 5420 6160 5430 6170
rect 6690 6160 6740 6170
rect 9270 6160 9340 6170
rect 9350 6160 9440 6170
rect 9450 6160 9460 6170
rect 9600 6160 9620 6170
rect 9670 6160 9690 6170
rect 9790 6160 9820 6170
rect 1270 6150 1290 6160
rect 1360 6150 1380 6160
rect 1600 6150 1610 6160
rect 1680 6150 1720 6160
rect 2450 6150 2460 6160
rect 4270 6150 4280 6160
rect 5300 6150 5310 6160
rect 5410 6150 5420 6160
rect 6690 6150 6750 6160
rect 6780 6150 6800 6160
rect 9240 6150 9470 6160
rect 9610 6150 9630 6160
rect 9640 6150 9690 6160
rect 9790 6150 9820 6160
rect 1280 6140 1300 6150
rect 1360 6140 1390 6150
rect 1430 6140 1440 6150
rect 1610 6140 1630 6150
rect 4280 6140 4290 6150
rect 5400 6140 5420 6150
rect 6710 6140 6750 6150
rect 6780 6140 6810 6150
rect 9220 6140 9480 6150
rect 9610 6140 9690 6150
rect 9800 6140 9830 6150
rect 1280 6130 1310 6140
rect 1360 6130 1390 6140
rect 1620 6130 1640 6140
rect 2430 6130 2440 6140
rect 4280 6130 4290 6140
rect 5290 6130 5300 6140
rect 5400 6130 5410 6140
rect 6720 6130 6760 6140
rect 6780 6130 6810 6140
rect 6830 6130 6840 6140
rect 9200 6130 9280 6140
rect 9300 6130 9480 6140
rect 9490 6130 9500 6140
rect 9630 6130 9690 6140
rect 9820 6130 9840 6140
rect 1290 6120 1320 6130
rect 1380 6120 1390 6130
rect 1440 6120 1450 6130
rect 1630 6120 1640 6130
rect 4290 6120 4300 6130
rect 5280 6120 5290 6130
rect 5390 6120 5400 6130
rect 6730 6120 6760 6130
rect 6780 6120 6840 6130
rect 9180 6120 9270 6130
rect 9350 6120 9470 6130
rect 9640 6120 9690 6130
rect 9820 6120 9840 6130
rect 1290 6110 1330 6120
rect 1380 6110 1400 6120
rect 1440 6110 1450 6120
rect 1630 6110 1650 6120
rect 3790 6110 3800 6120
rect 5280 6110 5290 6120
rect 5380 6110 5390 6120
rect 6730 6110 6830 6120
rect 9180 6110 9270 6120
rect 9360 6110 9480 6120
rect 9640 6110 9700 6120
rect 9830 6110 9850 6120
rect 1300 6100 1320 6110
rect 1330 6100 1340 6110
rect 1390 6100 1400 6110
rect 1590 6100 1650 6110
rect 2440 6100 2450 6110
rect 3790 6100 3800 6110
rect 4300 6100 4310 6110
rect 5270 6100 5280 6110
rect 5380 6100 5390 6110
rect 6730 6100 6830 6110
rect 9160 6100 9240 6110
rect 9390 6100 9410 6110
rect 9460 6100 9490 6110
rect 9600 6100 9610 6110
rect 9640 6100 9700 6110
rect 9830 6100 9850 6110
rect 1300 6090 1320 6100
rect 1340 6090 1360 6100
rect 1370 6090 1380 6100
rect 1390 6090 1410 6100
rect 1590 6090 1640 6100
rect 1770 6090 1780 6100
rect 2440 6090 2450 6100
rect 3790 6090 3800 6100
rect 3950 6090 3960 6100
rect 5370 6090 5380 6100
rect 6750 6090 6840 6100
rect 9120 6090 9250 6100
rect 9360 6090 9380 6100
rect 9480 6090 9520 6100
rect 9640 6090 9700 6100
rect 1340 6080 1390 6090
rect 1400 6080 1420 6090
rect 1590 6080 1630 6090
rect 1770 6080 1790 6090
rect 3780 6080 3800 6090
rect 3960 6080 3970 6090
rect 4310 6080 4320 6090
rect 5260 6080 5270 6090
rect 5360 6080 5380 6090
rect 6760 6080 6840 6090
rect 9120 6080 9260 6090
rect 9340 6080 9350 6090
rect 9490 6080 9520 6090
rect 9640 6080 9710 6090
rect 9850 6080 9860 6090
rect 1320 6070 1330 6080
rect 1350 6070 1380 6080
rect 1410 6070 1420 6080
rect 1590 6070 1610 6080
rect 1780 6070 1790 6080
rect 2450 6070 2460 6080
rect 3780 6070 3800 6080
rect 3860 6070 3870 6080
rect 5360 6070 5370 6080
rect 6760 6070 6770 6080
rect 6780 6070 6850 6080
rect 9090 6070 9220 6080
rect 9240 6070 9250 6080
rect 9330 6070 9340 6080
rect 9490 6070 9530 6080
rect 9640 6070 9710 6080
rect 9850 6070 9860 6080
rect 1310 6060 1340 6070
rect 1350 6060 1390 6070
rect 1410 6060 1420 6070
rect 1600 6060 1610 6070
rect 2450 6060 2460 6070
rect 2480 6060 2490 6070
rect 3240 6060 3260 6070
rect 3790 6060 3800 6070
rect 3820 6060 3840 6070
rect 5250 6060 5260 6070
rect 5360 6060 5370 6070
rect 6790 6060 6850 6070
rect 9080 6060 9230 6070
rect 9270 6060 9340 6070
rect 9430 6060 9440 6070
rect 9490 6060 9530 6070
rect 9630 6060 9710 6070
rect 9850 6060 9860 6070
rect 1330 6050 1340 6060
rect 1360 6050 1380 6060
rect 1410 6050 1430 6060
rect 1600 6050 1610 6060
rect 3230 6050 3280 6060
rect 5240 6050 5250 6060
rect 5360 6050 5370 6060
rect 6770 6050 6830 6060
rect 9080 6050 9240 6060
rect 9300 6050 9340 6060
rect 9390 6050 9440 6060
rect 9490 6050 9530 6060
rect 9640 6050 9720 6060
rect 1320 6040 1340 6050
rect 1360 6040 1370 6050
rect 1420 6040 1430 6050
rect 2490 6040 2500 6050
rect 3220 6040 3290 6050
rect 4330 6040 4340 6050
rect 5360 6040 5370 6050
rect 6780 6040 6810 6050
rect 9050 6040 9060 6050
rect 9070 6040 9210 6050
rect 9300 6040 9340 6050
rect 9390 6040 9440 6050
rect 9490 6040 9520 6050
rect 9640 6040 9720 6050
rect 1210 6030 1230 6040
rect 1320 6030 1330 6040
rect 1420 6030 1430 6040
rect 1610 6030 1620 6040
rect 3210 6030 3290 6040
rect 3780 6030 3790 6040
rect 5360 6030 5370 6040
rect 6770 6030 6810 6040
rect 6840 6030 6850 6040
rect 9020 6030 9190 6040
rect 9300 6030 9340 6040
rect 9400 6030 9430 6040
rect 9490 6030 9520 6040
rect 9650 6030 9720 6040
rect 9850 6030 9860 6040
rect 1170 6020 1190 6030
rect 1220 6020 1230 6030
rect 1300 6020 1310 6030
rect 1320 6020 1330 6030
rect 1420 6020 1430 6030
rect 1610 6020 1620 6030
rect 1680 6020 1700 6030
rect 3200 6020 3230 6030
rect 3240 6020 3290 6030
rect 5220 6020 5240 6030
rect 5360 6020 5370 6030
rect 6770 6020 6820 6030
rect 8850 6020 8900 6030
rect 8910 6020 9180 6030
rect 9280 6020 9290 6030
rect 9320 6020 9350 6030
rect 9400 6020 9410 6030
rect 9480 6020 9520 6030
rect 9650 6020 9720 6030
rect 9850 6020 9860 6030
rect 850 6010 890 6020
rect 1150 6010 1170 6020
rect 1200 6010 1220 6020
rect 1230 6010 1250 6020
rect 1280 6010 1310 6020
rect 1320 6010 1340 6020
rect 1420 6010 1430 6020
rect 1620 6010 1640 6020
rect 1660 6010 1670 6020
rect 1680 6010 1710 6020
rect 3190 6010 3290 6020
rect 3790 6010 3800 6020
rect 4340 6010 4350 6020
rect 5220 6010 5230 6020
rect 5350 6010 5360 6020
rect 6790 6010 6810 6020
rect 8830 6010 9100 6020
rect 9140 6010 9180 6020
rect 9250 6010 9280 6020
rect 9310 6010 9350 6020
rect 9470 6010 9500 6020
rect 9600 6010 9610 6020
rect 9650 6010 9720 6020
rect 9850 6010 9870 6020
rect 850 6000 910 6010
rect 1200 6000 1220 6010
rect 1240 6000 1250 6010
rect 1280 6000 1340 6010
rect 1420 6000 1430 6010
rect 1620 6000 1640 6010
rect 1660 6000 1670 6010
rect 1680 6000 1700 6010
rect 3180 6000 3200 6010
rect 3230 6000 3290 6010
rect 3800 6000 3810 6010
rect 4340 6000 4350 6010
rect 5340 6000 5350 6010
rect 6800 6000 6810 6010
rect 6820 6000 6850 6010
rect 6920 6000 6930 6010
rect 8820 6000 9090 6010
rect 9150 6000 9170 6010
rect 9230 6000 9300 6010
rect 9310 6000 9350 6010
rect 9460 6000 9480 6010
rect 9660 6000 9720 6010
rect 9870 6000 9880 6010
rect 850 5990 860 6000
rect 880 5990 920 6000
rect 1170 5990 1190 6000
rect 1210 5990 1230 6000
rect 1270 5990 1300 6000
rect 1310 5990 1340 6000
rect 1420 5990 1430 6000
rect 1630 5990 1650 6000
rect 1660 5990 1700 6000
rect 3170 5990 3180 6000
rect 3240 5990 3290 6000
rect 3790 5990 3800 6000
rect 4340 5990 4350 6000
rect 5200 5990 5210 6000
rect 5340 5990 5360 6000
rect 6800 5990 6860 6000
rect 6910 5990 6940 6000
rect 8800 5990 9040 6000
rect 9070 5990 9080 6000
rect 9150 5990 9170 6000
rect 9230 5990 9350 6000
rect 9460 5990 9470 6000
rect 9670 5990 9730 6000
rect 9880 5990 9900 6000
rect 850 5980 880 5990
rect 910 5980 920 5990
rect 1140 5980 1170 5990
rect 1200 5980 1220 5990
rect 1250 5980 1300 5990
rect 1630 5980 1650 5990
rect 1660 5980 1690 5990
rect 3160 5980 3180 5990
rect 3250 5980 3290 5990
rect 3830 5980 3840 5990
rect 4340 5980 4350 5990
rect 5190 5980 5200 5990
rect 5340 5980 5360 5990
rect 6810 5980 6950 5990
rect 8770 5980 9020 5990
rect 9150 5980 9160 5990
rect 9240 5980 9280 5990
rect 9300 5980 9310 5990
rect 9320 5980 9350 5990
rect 9470 5980 9480 5990
rect 9660 5980 9730 5990
rect 850 5970 870 5980
rect 910 5970 930 5980
rect 1130 5970 1160 5980
rect 1190 5970 1200 5980
rect 1260 5970 1290 5980
rect 1640 5970 1670 5980
rect 1680 5970 1690 5980
rect 3160 5970 3170 5980
rect 3250 5970 3290 5980
rect 4340 5970 4350 5980
rect 5340 5970 5350 5980
rect 6820 5970 6950 5980
rect 8760 5970 8970 5980
rect 9000 5970 9010 5980
rect 9310 5970 9360 5980
rect 9480 5970 9490 5980
rect 9680 5970 9740 5980
rect 850 5960 860 5970
rect 920 5960 950 5970
rect 1120 5960 1160 5970
rect 1180 5960 1190 5970
rect 1260 5960 1280 5970
rect 1670 5960 1680 5970
rect 3150 5960 3170 5970
rect 3250 5960 3290 5970
rect 3850 5960 3860 5970
rect 4100 5960 4110 5970
rect 4340 5960 4350 5970
rect 5340 5960 5350 5970
rect 6820 5960 6960 5970
rect 8650 5960 8670 5970
rect 8680 5960 8960 5970
rect 9150 5960 9160 5970
rect 9310 5960 9360 5970
rect 9420 5960 9430 5970
rect 9680 5960 9740 5970
rect 9880 5960 9890 5970
rect 850 5950 860 5960
rect 980 5950 1000 5960
rect 1070 5950 1090 5960
rect 1100 5950 1160 5960
rect 1180 5950 1190 5960
rect 1200 5950 1210 5960
rect 1260 5950 1280 5960
rect 1670 5950 1680 5960
rect 3140 5950 3160 5960
rect 3250 5950 3280 5960
rect 5330 5950 5340 5960
rect 6820 5950 6950 5960
rect 6960 5950 6970 5960
rect 8620 5950 8630 5960
rect 8640 5950 8960 5960
rect 9320 5950 9360 5960
rect 9420 5950 9440 5960
rect 9670 5950 9740 5960
rect 9890 5950 9900 5960
rect 9920 5950 9940 5960
rect 980 5940 990 5950
rect 1000 5940 1040 5950
rect 1060 5940 1140 5950
rect 1150 5940 1170 5950
rect 1180 5940 1190 5950
rect 1260 5940 1280 5950
rect 1670 5940 1680 5950
rect 3130 5940 3150 5950
rect 3250 5940 3280 5950
rect 3880 5940 3890 5950
rect 4330 5940 4340 5950
rect 5330 5940 5340 5950
rect 6830 5940 6940 5950
rect 8590 5940 8950 5950
rect 9170 5940 9180 5950
rect 9290 5940 9300 5950
rect 9320 5940 9330 5950
rect 9340 5940 9370 5950
rect 9420 5940 9450 5950
rect 9510 5940 9520 5950
rect 9690 5940 9750 5950
rect 9890 5940 9900 5950
rect 730 5930 750 5940
rect 970 5930 980 5940
rect 1000 5930 1130 5940
rect 1160 5930 1190 5940
rect 1270 5930 1280 5940
rect 1670 5930 1690 5940
rect 3120 5930 3140 5940
rect 3250 5930 3280 5940
rect 3760 5930 3770 5940
rect 3890 5930 3900 5940
rect 4160 5930 4170 5940
rect 4330 5930 4340 5940
rect 5150 5930 5160 5940
rect 5330 5930 5340 5940
rect 6820 5930 6950 5940
rect 8570 5930 8850 5940
rect 8920 5930 8950 5940
rect 9260 5930 9320 5940
rect 9350 5930 9370 5940
rect 9420 5930 9460 5940
rect 9510 5930 9520 5940
rect 9690 5930 9750 5940
rect 9890 5930 9900 5940
rect 730 5920 740 5930
rect 950 5920 970 5930
rect 1010 5920 1020 5930
rect 1030 5920 1040 5930
rect 1050 5920 1070 5930
rect 1210 5920 1220 5930
rect 1230 5920 1240 5930
rect 1680 5920 1700 5930
rect 2570 5920 2580 5930
rect 3100 5920 3120 5930
rect 3260 5920 3280 5930
rect 3900 5920 3910 5930
rect 4180 5920 4190 5930
rect 5140 5920 5150 5930
rect 5330 5920 5340 5930
rect 6830 5920 6870 5930
rect 6900 5920 6950 5930
rect 8540 5920 8830 5930
rect 8930 5920 8940 5930
rect 9250 5920 9310 5930
rect 9320 5920 9340 5930
rect 9350 5920 9370 5930
rect 9430 5920 9480 5930
rect 9500 5920 9510 5930
rect 9700 5920 9760 5930
rect 9890 5920 9900 5930
rect 720 5910 740 5920
rect 1010 5910 1060 5920
rect 1210 5910 1230 5920
rect 1680 5910 1710 5920
rect 3090 5910 3120 5920
rect 3260 5910 3290 5920
rect 3900 5910 3910 5920
rect 4200 5910 4210 5920
rect 4320 5910 4330 5920
rect 5170 5910 5180 5920
rect 6830 5910 6860 5920
rect 6910 5910 6960 5920
rect 8100 5910 8120 5920
rect 8530 5910 8730 5920
rect 8750 5910 8810 5920
rect 9160 5910 9170 5920
rect 9260 5910 9310 5920
rect 9320 5910 9350 5920
rect 9360 5910 9370 5920
rect 9430 5910 9440 5920
rect 9450 5910 9470 5920
rect 9710 5910 9760 5920
rect 9890 5910 9910 5920
rect 720 5900 740 5910
rect 960 5900 970 5910
rect 1050 5900 1070 5910
rect 1130 5900 1140 5910
rect 1160 5900 1180 5910
rect 1190 5900 1210 5910
rect 1700 5900 1720 5910
rect 2600 5900 2610 5910
rect 3070 5900 3100 5910
rect 3260 5900 3300 5910
rect 3910 5900 3920 5910
rect 4220 5900 4230 5910
rect 4280 5900 4300 5910
rect 5130 5900 5160 5910
rect 5320 5900 5330 5910
rect 6820 5900 6860 5910
rect 6910 5900 6960 5910
rect 8100 5900 8120 5910
rect 8460 5900 8500 5910
rect 8510 5900 8730 5910
rect 8750 5900 8800 5910
rect 9160 5900 9180 5910
rect 9260 5900 9300 5910
rect 9340 5900 9350 5910
rect 9360 5900 9380 5910
rect 9420 5900 9430 5910
rect 9440 5900 9460 5910
rect 9720 5900 9750 5910
rect 9890 5900 9900 5910
rect 710 5890 730 5900
rect 970 5890 980 5900
rect 1020 5890 1070 5900
rect 1100 5890 1160 5900
rect 1170 5890 1200 5900
rect 1710 5890 1730 5900
rect 2610 5890 2620 5900
rect 3060 5890 3100 5900
rect 3250 5890 3290 5900
rect 3920 5890 3930 5900
rect 4240 5890 4260 5900
rect 5130 5890 5170 5900
rect 5310 5890 5330 5900
rect 6830 5890 6850 5900
rect 6910 5890 6960 5900
rect 8100 5890 8130 5900
rect 8440 5890 8700 5900
rect 8760 5890 8800 5900
rect 8860 5890 8870 5900
rect 9160 5890 9170 5900
rect 9190 5890 9200 5900
rect 9340 5890 9350 5900
rect 9380 5890 9390 5900
rect 9410 5890 9420 5900
rect 9720 5890 9750 5900
rect 9890 5890 9900 5900
rect 980 5880 990 5890
rect 1020 5880 1130 5890
rect 1720 5880 1740 5890
rect 2610 5880 2640 5890
rect 3040 5880 3080 5890
rect 3250 5880 3290 5890
rect 3740 5880 3750 5890
rect 5150 5880 5160 5890
rect 5320 5880 5330 5890
rect 6830 5880 6850 5890
rect 6910 5880 6960 5890
rect 8100 5880 8150 5890
rect 8400 5880 8680 5890
rect 8760 5880 8790 5890
rect 8850 5880 8870 5890
rect 8950 5880 8960 5890
rect 9340 5880 9350 5890
rect 9730 5880 9750 5890
rect 9900 5880 9920 5890
rect 710 5870 720 5880
rect 770 5870 780 5880
rect 1040 5870 1050 5880
rect 1130 5870 1140 5880
rect 1740 5870 1780 5880
rect 1810 5870 1840 5880
rect 2620 5870 2660 5880
rect 2990 5870 3060 5880
rect 3250 5870 3290 5880
rect 3930 5870 3940 5880
rect 5140 5870 5150 5880
rect 5320 5870 5330 5880
rect 6830 5870 6850 5880
rect 6910 5870 6960 5880
rect 8090 5870 8150 5880
rect 8360 5870 8650 5880
rect 8760 5870 8790 5880
rect 8840 5870 8880 5880
rect 9340 5870 9360 5880
rect 9730 5870 9740 5880
rect 9910 5870 9920 5880
rect 710 5860 720 5870
rect 1040 5860 1050 5870
rect 1750 5860 1830 5870
rect 2630 5860 2690 5870
rect 2980 5860 3040 5870
rect 3260 5860 3290 5870
rect 3740 5860 3760 5870
rect 3940 5860 3950 5870
rect 5310 5860 5320 5870
rect 6830 5860 6850 5870
rect 6920 5860 6970 5870
rect 7920 5860 7940 5870
rect 8090 5860 8140 5870
rect 8330 5860 8620 5870
rect 8740 5860 8790 5870
rect 8840 5860 8890 5870
rect 8960 5860 8970 5870
rect 9170 5860 9190 5870
rect 9320 5860 9360 5870
rect 9910 5860 9920 5870
rect 670 5850 690 5860
rect 700 5850 720 5860
rect 800 5850 820 5860
rect 830 5850 870 5860
rect 970 5850 990 5860
rect 1840 5850 1850 5860
rect 2650 5850 2700 5860
rect 2930 5850 3000 5860
rect 3270 5850 3290 5860
rect 3730 5850 3740 5860
rect 3750 5850 3760 5860
rect 3940 5850 3950 5860
rect 5110 5850 5120 5860
rect 5130 5850 5140 5860
rect 5310 5850 5320 5860
rect 6830 5850 6850 5860
rect 6930 5850 6990 5860
rect 7910 5850 7950 5860
rect 8100 5850 8140 5860
rect 8300 5850 8620 5860
rect 8720 5850 8790 5860
rect 8840 5850 8900 5860
rect 8960 5850 8980 5860
rect 9070 5850 9080 5860
rect 9170 5850 9200 5860
rect 9280 5850 9320 5860
rect 9900 5850 9920 5860
rect 660 5840 720 5850
rect 730 5840 740 5850
rect 790 5840 810 5850
rect 830 5840 860 5850
rect 870 5840 880 5850
rect 970 5840 990 5850
rect 2660 5840 2710 5850
rect 2890 5840 2980 5850
rect 3260 5840 3290 5850
rect 3750 5840 3760 5850
rect 3800 5840 3830 5850
rect 5110 5840 5130 5850
rect 5310 5840 5320 5850
rect 6830 5840 6850 5850
rect 6920 5840 6990 5850
rect 7890 5840 7950 5850
rect 8100 5840 8130 5850
rect 8260 5840 8620 5850
rect 8720 5840 8790 5850
rect 8850 5840 8900 5850
rect 8960 5840 8980 5850
rect 9070 5840 9090 5850
rect 9170 5840 9210 5850
rect 9220 5840 9240 5850
rect 9250 5840 9340 5850
rect 9900 5840 9910 5850
rect 660 5830 740 5840
rect 780 5830 820 5840
rect 880 5830 890 5840
rect 910 5830 950 5840
rect 2670 5830 2710 5840
rect 2860 5830 2980 5840
rect 3260 5830 3290 5840
rect 3860 5830 3870 5840
rect 3950 5830 3960 5840
rect 5110 5830 5130 5840
rect 5300 5830 5320 5840
rect 6830 5830 6840 5840
rect 6920 5830 6980 5840
rect 7900 5830 7960 5840
rect 8100 5830 8110 5840
rect 8240 5830 8620 5840
rect 8720 5830 8800 5840
rect 8850 5830 8900 5840
rect 8960 5830 8990 5840
rect 9070 5830 9100 5840
rect 9170 5830 9330 5840
rect 9910 5830 9920 5840
rect 660 5820 740 5830
rect 790 5820 820 5830
rect 2670 5820 2740 5830
rect 2840 5820 2880 5830
rect 2930 5820 2950 5830
rect 3260 5820 3290 5830
rect 3720 5820 3730 5830
rect 3950 5820 3960 5830
rect 5110 5820 5120 5830
rect 5300 5820 5320 5830
rect 6830 5820 6850 5830
rect 6920 5820 6980 5830
rect 7900 5820 7970 5830
rect 8210 5820 8660 5830
rect 8720 5820 8800 5830
rect 8850 5820 8910 5830
rect 8970 5820 8990 5830
rect 9070 5820 9110 5830
rect 9160 5820 9310 5830
rect 9920 5820 9940 5830
rect 660 5810 730 5820
rect 810 5810 820 5820
rect 840 5810 880 5820
rect 1010 5810 1020 5820
rect 2690 5810 2870 5820
rect 3260 5810 3290 5820
rect 5110 5810 5120 5820
rect 5300 5810 5320 5820
rect 6830 5810 6850 5820
rect 6910 5810 6970 5820
rect 7900 5810 7970 5820
rect 8180 5810 8670 5820
rect 8730 5810 8790 5820
rect 8850 5810 8910 5820
rect 8970 5810 8990 5820
rect 9070 5810 9300 5820
rect 9930 5810 9940 5820
rect 580 5800 590 5810
rect 660 5800 730 5810
rect 810 5800 820 5810
rect 890 5800 900 5810
rect 2700 5800 2850 5810
rect 3260 5800 3290 5810
rect 3740 5800 3750 5810
rect 3800 5800 3810 5810
rect 5100 5800 5110 5810
rect 5300 5800 5320 5810
rect 6830 5800 6850 5810
rect 6910 5800 6970 5810
rect 7950 5800 7990 5810
rect 8150 5800 8670 5810
rect 8730 5800 8750 5810
rect 8760 5800 8800 5810
rect 8860 5800 8900 5810
rect 8970 5800 9000 5810
rect 9070 5800 9260 5810
rect 9930 5800 9940 5810
rect 580 5790 600 5800
rect 660 5790 700 5800
rect 800 5790 810 5800
rect 900 5790 910 5800
rect 2690 5790 2830 5800
rect 3260 5790 3300 5800
rect 3770 5790 3800 5800
rect 3810 5790 3820 5800
rect 3830 5790 3840 5800
rect 3860 5790 3880 5800
rect 3960 5790 3970 5800
rect 5300 5790 5310 5800
rect 6830 5790 6850 5800
rect 6910 5790 6920 5800
rect 6940 5790 6980 5800
rect 8120 5790 8390 5800
rect 8410 5790 8670 5800
rect 8730 5790 8740 5800
rect 8750 5790 8810 5800
rect 8860 5790 8900 5800
rect 8970 5790 9010 5800
rect 9060 5790 9250 5800
rect 9930 5790 9940 5800
rect 570 5780 590 5790
rect 790 5780 800 5790
rect 2300 5780 2320 5790
rect 2670 5780 2830 5790
rect 3260 5780 3290 5790
rect 3800 5780 3840 5790
rect 3860 5780 3880 5790
rect 5300 5780 5310 5790
rect 6830 5780 6850 5790
rect 6900 5780 6920 5790
rect 6940 5780 6980 5790
rect 8080 5780 8380 5790
rect 8420 5780 8680 5790
rect 8730 5780 8810 5790
rect 8870 5780 8890 5790
rect 8960 5780 9220 5790
rect 9240 5780 9250 5790
rect 9930 5780 9940 5790
rect 800 5770 810 5780
rect 900 5770 910 5780
rect 1850 5770 1870 5780
rect 2280 5770 2310 5780
rect 2670 5770 2810 5780
rect 3260 5770 3300 5780
rect 3780 5770 3800 5780
rect 3830 5770 3850 5780
rect 3970 5770 3980 5780
rect 5300 5770 5310 5780
rect 6840 5770 6860 5780
rect 6910 5770 6920 5780
rect 6930 5770 6980 5780
rect 8050 5770 8380 5780
rect 8420 5770 8680 5780
rect 8730 5770 8810 5780
rect 8950 5770 9090 5780
rect 9160 5770 9230 5780
rect 9930 5770 9940 5780
rect 790 5760 820 5770
rect 880 5760 890 5770
rect 1850 5760 1870 5770
rect 2270 5760 2310 5770
rect 2650 5760 2800 5770
rect 3260 5760 3300 5770
rect 3770 5760 3790 5770
rect 3850 5760 3890 5770
rect 3970 5760 3980 5770
rect 5100 5760 5110 5770
rect 5290 5760 5300 5770
rect 6840 5760 6870 5770
rect 6930 5760 6980 5770
rect 8020 5760 8380 5770
rect 8430 5760 8690 5770
rect 8740 5760 8760 5770
rect 8770 5760 8820 5770
rect 8940 5760 9070 5770
rect 9180 5760 9200 5770
rect 9930 5760 9940 5770
rect 800 5750 810 5760
rect 1850 5750 1870 5760
rect 2260 5750 2300 5760
rect 2640 5750 2710 5760
rect 2740 5750 2790 5760
rect 3260 5750 3300 5760
rect 3720 5750 3740 5760
rect 3760 5750 3820 5760
rect 3830 5750 3840 5760
rect 3860 5750 3890 5760
rect 3910 5750 3930 5760
rect 3980 5750 3990 5760
rect 5090 5750 5110 5760
rect 5290 5750 5300 5760
rect 6840 5750 6900 5760
rect 6930 5750 6970 5760
rect 7990 5750 8380 5760
rect 8430 5750 8690 5760
rect 8740 5750 8760 5760
rect 8780 5750 8830 5760
rect 8930 5750 9070 5760
rect 9930 5750 9940 5760
rect 1850 5740 1870 5750
rect 2250 5740 2290 5750
rect 2620 5740 2690 5750
rect 2740 5740 2780 5750
rect 3260 5740 3300 5750
rect 3720 5740 3730 5750
rect 3790 5740 3800 5750
rect 3840 5740 3920 5750
rect 6840 5740 6930 5750
rect 6950 5740 6970 5750
rect 7960 5740 8250 5750
rect 8280 5740 8380 5750
rect 8430 5740 8690 5750
rect 8740 5740 8760 5750
rect 8800 5740 8840 5750
rect 8910 5740 9040 5750
rect 9930 5740 9950 5750
rect 660 5730 680 5740
rect 720 5730 820 5740
rect 850 5730 870 5740
rect 1850 5730 1860 5740
rect 2250 5730 2290 5740
rect 2610 5730 2680 5740
rect 2720 5730 2760 5740
rect 3260 5730 3310 5740
rect 3710 5730 3720 5740
rect 3810 5730 3840 5740
rect 3880 5730 3890 5740
rect 3930 5730 3940 5740
rect 3970 5730 3990 5740
rect 5080 5730 5100 5740
rect 5280 5730 5290 5740
rect 6840 5730 6930 5740
rect 6950 5730 6970 5740
rect 7920 5730 8240 5740
rect 8280 5730 8380 5740
rect 8430 5730 8690 5740
rect 8760 5730 8770 5740
rect 8800 5730 9050 5740
rect 9930 5730 9950 5740
rect 1230 5720 1250 5730
rect 2240 5720 2280 5730
rect 2580 5720 2660 5730
rect 2710 5720 2770 5730
rect 3260 5720 3320 5730
rect 3700 5720 3710 5730
rect 3750 5720 3760 5730
rect 3830 5720 3850 5730
rect 3960 5720 3980 5730
rect 5080 5720 5100 5730
rect 5130 5720 5140 5730
rect 5280 5720 5290 5730
rect 6840 5720 6910 5730
rect 6930 5720 6970 5730
rect 7910 5720 8180 5730
rect 8220 5720 8230 5730
rect 8290 5720 8390 5730
rect 8440 5720 8700 5730
rect 8810 5720 9030 5730
rect 9930 5720 9950 5730
rect 780 5710 790 5720
rect 1200 5710 1210 5720
rect 1230 5710 1240 5720
rect 2240 5710 2280 5720
rect 2570 5710 2630 5720
rect 2690 5710 2760 5720
rect 3260 5710 3310 5720
rect 3720 5710 3750 5720
rect 3770 5710 3780 5720
rect 3850 5710 3870 5720
rect 5080 5710 5100 5720
rect 5110 5710 5130 5720
rect 6850 5710 6900 5720
rect 6950 5710 6960 5720
rect 7910 5710 8170 5720
rect 8220 5710 8240 5720
rect 8290 5710 8390 5720
rect 8440 5710 8600 5720
rect 8610 5710 8640 5720
rect 8650 5710 8700 5720
rect 8830 5710 8840 5720
rect 8920 5710 8930 5720
rect 8940 5710 8960 5720
rect 8970 5710 9040 5720
rect 9930 5710 9950 5720
rect 800 5700 810 5710
rect 1160 5700 1170 5710
rect 1220 5700 1230 5710
rect 1610 5700 1620 5710
rect 2230 5700 2280 5710
rect 2560 5700 2620 5710
rect 2680 5700 2720 5710
rect 2750 5700 2760 5710
rect 3260 5700 3320 5710
rect 3670 5700 3680 5710
rect 3720 5700 3750 5710
rect 3770 5700 3780 5710
rect 3800 5700 3820 5710
rect 3870 5700 3880 5710
rect 5080 5700 5110 5710
rect 5120 5700 5130 5710
rect 5280 5700 5290 5710
rect 6850 5700 6930 5710
rect 7920 5700 8120 5710
rect 8290 5700 8390 5710
rect 8440 5700 8620 5710
rect 8650 5700 8700 5710
rect 8750 5700 8760 5710
rect 8950 5700 9050 5710
rect 9950 5700 9960 5710
rect 1050 5690 1060 5700
rect 1120 5690 1130 5700
rect 1200 5690 1220 5700
rect 1610 5690 1620 5700
rect 1860 5690 1870 5700
rect 2220 5690 2270 5700
rect 2550 5690 2590 5700
rect 2660 5690 2710 5700
rect 2750 5690 2760 5700
rect 3260 5690 3310 5700
rect 3670 5690 3680 5700
rect 3710 5690 3750 5700
rect 3760 5690 3770 5700
rect 3810 5690 3820 5700
rect 3840 5690 3860 5700
rect 3910 5690 3920 5700
rect 5080 5690 5100 5700
rect 5120 5690 5150 5700
rect 6860 5690 6910 5700
rect 6930 5690 6940 5700
rect 7800 5690 7810 5700
rect 7920 5690 8110 5700
rect 8290 5690 8390 5700
rect 8440 5690 8630 5700
rect 8650 5690 8720 5700
rect 8740 5690 8760 5700
rect 8950 5690 9040 5700
rect 9950 5690 9990 5700
rect 820 5680 840 5690
rect 1040 5680 1070 5690
rect 1180 5680 1190 5690
rect 2220 5680 2260 5690
rect 2540 5680 2590 5690
rect 2650 5680 2690 5690
rect 2750 5680 2770 5690
rect 3270 5680 3310 5690
rect 3720 5680 3770 5690
rect 3780 5680 3790 5690
rect 3810 5680 3820 5690
rect 3880 5680 3910 5690
rect 3930 5680 3940 5690
rect 5080 5680 5090 5690
rect 5120 5680 5150 5690
rect 6860 5680 6910 5690
rect 7750 5680 7810 5690
rect 7920 5680 8030 5690
rect 8060 5680 8100 5690
rect 8290 5680 8390 5690
rect 8450 5680 8570 5690
rect 8600 5680 8750 5690
rect 8860 5680 8870 5690
rect 8880 5680 8890 5690
rect 8940 5680 8990 5690
rect 830 5670 840 5680
rect 1150 5670 1190 5680
rect 1860 5670 1870 5680
rect 2220 5670 2260 5680
rect 2530 5670 2590 5680
rect 2630 5670 2680 5680
rect 3270 5670 3310 5680
rect 3700 5670 3710 5680
rect 3720 5670 3790 5680
rect 3800 5670 3810 5680
rect 3830 5670 3840 5680
rect 3850 5670 3860 5680
rect 3870 5670 3890 5680
rect 3920 5670 3950 5680
rect 3990 5670 4000 5680
rect 5130 5670 5150 5680
rect 5270 5670 5280 5680
rect 6860 5670 6910 5680
rect 6950 5670 6960 5680
rect 7730 5670 7820 5680
rect 7920 5670 8020 5680
rect 8070 5670 8090 5680
rect 8300 5670 8400 5680
rect 8450 5670 8520 5680
rect 8530 5670 8580 5680
rect 8620 5670 8640 5680
rect 8670 5670 8740 5680
rect 8880 5670 8900 5680
rect 8940 5670 8990 5680
rect 9990 5670 9990 5680
rect 810 5660 830 5670
rect 1860 5660 1870 5670
rect 2210 5660 2250 5670
rect 2530 5660 2580 5670
rect 2590 5660 2650 5670
rect 3260 5660 3310 5670
rect 3660 5660 3670 5670
rect 3690 5660 3730 5670
rect 3760 5660 3770 5670
rect 3780 5660 3790 5670
rect 3800 5660 3840 5670
rect 3870 5660 3890 5670
rect 3910 5660 3950 5670
rect 5270 5660 5280 5670
rect 6860 5660 6890 5670
rect 6920 5660 6930 5670
rect 7720 5660 7820 5670
rect 7920 5660 8010 5670
rect 8080 5660 8090 5670
rect 8300 5660 8400 5670
rect 8450 5660 8500 5670
rect 8520 5660 8560 5670
rect 8650 5660 8680 5670
rect 8700 5660 8710 5670
rect 8720 5660 8730 5670
rect 8970 5660 8980 5670
rect 9990 5660 9990 5670
rect 810 5650 820 5660
rect 1870 5650 1880 5660
rect 2210 5650 2250 5660
rect 2520 5650 2570 5660
rect 2580 5650 2660 5660
rect 3260 5650 3310 5660
rect 3660 5650 3670 5660
rect 3680 5650 3690 5660
rect 3720 5650 3730 5660
rect 3760 5650 3770 5660
rect 3820 5650 3850 5660
rect 5130 5650 5140 5660
rect 5270 5650 5280 5660
rect 6870 5650 6880 5660
rect 6930 5650 6940 5660
rect 7710 5650 7820 5660
rect 7920 5650 8010 5660
rect 8070 5650 8090 5660
rect 8300 5650 8400 5660
rect 8450 5650 8470 5660
rect 8530 5650 8550 5660
rect 8610 5650 8620 5660
rect 8670 5650 8680 5660
rect 9980 5650 9990 5660
rect 800 5640 810 5650
rect 1870 5640 1880 5650
rect 2210 5640 2250 5650
rect 2500 5640 2640 5650
rect 3260 5640 3300 5650
rect 3700 5640 3720 5650
rect 3750 5640 3760 5650
rect 3780 5640 3790 5650
rect 3810 5640 3830 5650
rect 3850 5640 3860 5650
rect 3910 5640 3920 5650
rect 3930 5640 3940 5650
rect 5270 5640 5280 5650
rect 6870 5640 6880 5650
rect 6940 5640 6950 5650
rect 7690 5640 7820 5650
rect 7920 5640 8010 5650
rect 8080 5640 8090 5650
rect 8300 5640 8390 5650
rect 8530 5640 8560 5650
rect 8630 5640 8640 5650
rect 9980 5640 9990 5650
rect 770 5630 790 5640
rect 1860 5630 1890 5640
rect 2200 5630 2240 5640
rect 2500 5630 2640 5640
rect 3270 5630 3300 5640
rect 3700 5630 3710 5640
rect 3740 5630 3750 5640
rect 3770 5630 3790 5640
rect 3800 5630 3810 5640
rect 3860 5630 3870 5640
rect 5120 5630 5130 5640
rect 5270 5630 5280 5640
rect 6870 5630 6890 5640
rect 6940 5630 6960 5640
rect 7700 5630 7830 5640
rect 7920 5630 8000 5640
rect 8310 5630 8400 5640
rect 8530 5630 8550 5640
rect 8700 5630 8710 5640
rect 8720 5630 8730 5640
rect 8920 5630 8940 5640
rect 9960 5630 9980 5640
rect 750 5620 760 5630
rect 1860 5620 1890 5630
rect 1900 5620 1930 5630
rect 2190 5620 2240 5630
rect 2480 5620 2640 5630
rect 3260 5620 3300 5630
rect 3700 5620 3740 5630
rect 3790 5620 3800 5630
rect 6880 5620 6890 5630
rect 6940 5620 6960 5630
rect 7690 5620 7820 5630
rect 7930 5620 8010 5630
rect 8310 5620 8400 5630
rect 8510 5620 8540 5630
rect 8920 5620 8950 5630
rect 9960 5620 9980 5630
rect 730 5610 740 5620
rect 1860 5610 1930 5620
rect 2190 5610 2240 5620
rect 2470 5610 2630 5620
rect 3270 5610 3300 5620
rect 3670 5610 3700 5620
rect 5640 5610 5740 5620
rect 6880 5610 6890 5620
rect 6940 5610 6950 5620
rect 7680 5610 7800 5620
rect 7930 5610 8010 5620
rect 8310 5610 8340 5620
rect 8390 5610 8400 5620
rect 8470 5610 8500 5620
rect 8920 5610 8950 5620
rect 9960 5610 9970 5620
rect 1860 5600 1940 5610
rect 2190 5600 2240 5610
rect 2470 5600 2640 5610
rect 3270 5600 3310 5610
rect 3420 5600 3430 5610
rect 3650 5600 3660 5610
rect 3690 5600 3710 5610
rect 5110 5600 5120 5610
rect 5590 5600 5670 5610
rect 5700 5600 5770 5610
rect 6880 5600 6890 5610
rect 6930 5600 6950 5610
rect 7500 5600 7510 5610
rect 7520 5600 7530 5610
rect 7570 5600 7590 5610
rect 7680 5600 7790 5610
rect 7930 5600 8010 5610
rect 8400 5600 8460 5610
rect 8950 5600 8960 5610
rect 8980 5600 9010 5610
rect 9060 5600 9070 5610
rect 9960 5600 9980 5610
rect 700 5590 720 5600
rect 1870 5590 1940 5600
rect 2190 5590 2240 5600
rect 2470 5590 2610 5600
rect 2860 5590 2880 5600
rect 3270 5590 3310 5600
rect 3650 5590 3660 5600
rect 3700 5590 3710 5600
rect 3740 5590 3760 5600
rect 3770 5590 3780 5600
rect 5260 5590 5270 5600
rect 5580 5590 5640 5600
rect 5780 5590 5840 5600
rect 6890 5590 6900 5600
rect 6930 5590 6950 5600
rect 7460 5590 7540 5600
rect 7570 5590 7600 5600
rect 7680 5590 7780 5600
rect 7940 5590 8010 5600
rect 8390 5590 8430 5600
rect 8940 5590 8960 5600
rect 8970 5590 8980 5600
rect 9970 5590 9980 5600
rect 680 5580 690 5590
rect 1860 5580 1940 5590
rect 2190 5580 2230 5590
rect 2450 5580 2620 5590
rect 2870 5580 2890 5590
rect 3270 5580 3310 5590
rect 3650 5580 3670 5590
rect 4190 5580 4200 5590
rect 5110 5580 5120 5590
rect 5260 5580 5270 5590
rect 5580 5580 5640 5590
rect 5810 5580 5850 5590
rect 6890 5580 6900 5590
rect 6930 5580 6950 5590
rect 7430 5580 7610 5590
rect 7690 5580 7700 5590
rect 7760 5580 7780 5590
rect 7940 5580 8010 5590
rect 8380 5580 8410 5590
rect 8930 5580 8970 5590
rect 9980 5580 9990 5590
rect 670 5570 690 5580
rect 1870 5570 1940 5580
rect 2190 5570 2230 5580
rect 2450 5570 2620 5580
rect 2880 5570 2910 5580
rect 3270 5570 3310 5580
rect 3640 5570 3660 5580
rect 3700 5570 3710 5580
rect 4190 5570 4210 5580
rect 5590 5570 5640 5580
rect 5830 5570 5870 5580
rect 6330 5570 6420 5580
rect 6890 5570 6900 5580
rect 6920 5570 6950 5580
rect 7390 5570 7540 5580
rect 7550 5570 7610 5580
rect 7770 5570 7790 5580
rect 7950 5570 8020 5580
rect 8090 5570 8100 5580
rect 8110 5570 8120 5580
rect 8350 5570 8400 5580
rect 8900 5570 8960 5580
rect 9090 5570 9100 5580
rect 9990 5570 9990 5580
rect 660 5560 680 5570
rect 1870 5560 1930 5570
rect 2190 5560 2230 5570
rect 2430 5560 2620 5570
rect 2900 5560 2920 5570
rect 3260 5560 3310 5570
rect 3640 5560 3660 5570
rect 3670 5560 3680 5570
rect 3700 5560 3710 5570
rect 3730 5560 3740 5570
rect 3750 5560 3770 5570
rect 4200 5560 4210 5570
rect 5590 5560 5630 5570
rect 5850 5560 5880 5570
rect 6290 5560 6450 5570
rect 6890 5560 6900 5570
rect 6920 5560 6950 5570
rect 7370 5560 7610 5570
rect 7760 5560 7790 5570
rect 7940 5560 8020 5570
rect 8250 5560 8280 5570
rect 8320 5560 8330 5570
rect 8340 5560 8370 5570
rect 8860 5560 8870 5570
rect 8900 5560 8950 5570
rect 9030 5560 9040 5570
rect 9090 5560 9100 5570
rect 9990 5560 9990 5570
rect 660 5550 670 5560
rect 1870 5550 1940 5560
rect 2190 5550 2230 5560
rect 2430 5550 2530 5560
rect 2540 5550 2600 5560
rect 2920 5550 2940 5560
rect 3260 5550 3310 5560
rect 3650 5550 3660 5560
rect 3690 5550 3700 5560
rect 3770 5550 3780 5560
rect 5630 5550 5680 5560
rect 5850 5550 5900 5560
rect 6270 5550 6340 5560
rect 6400 5550 6500 5560
rect 6900 5550 6910 5560
rect 6930 5550 6960 5560
rect 7380 5550 7620 5560
rect 7750 5550 7790 5560
rect 7950 5550 8020 5560
rect 8190 5550 8200 5560
rect 8250 5550 8360 5560
rect 8840 5550 8850 5560
rect 8900 5550 8950 5560
rect 9000 5550 9060 5560
rect 9080 5550 9090 5560
rect 580 5540 600 5550
rect 1880 5540 1940 5550
rect 2190 5540 2230 5550
rect 2430 5540 2490 5550
rect 2500 5540 2590 5550
rect 2930 5540 2950 5550
rect 3260 5540 3310 5550
rect 3490 5540 3500 5550
rect 3650 5540 3660 5550
rect 3720 5540 3730 5550
rect 3740 5540 3750 5550
rect 3760 5540 3770 5550
rect 3780 5540 3790 5550
rect 5120 5540 5150 5550
rect 5650 5540 5760 5550
rect 5860 5540 5900 5550
rect 6260 5540 6300 5550
rect 6440 5540 6540 5550
rect 6900 5540 6950 5550
rect 7380 5540 7620 5550
rect 7720 5540 7790 5550
rect 7950 5540 8020 5550
rect 8110 5540 8120 5550
rect 8190 5540 8210 5550
rect 8240 5540 8300 5550
rect 8780 5540 8790 5550
rect 8850 5540 8860 5550
rect 8910 5540 8940 5550
rect 9000 5540 9050 5550
rect 9060 5540 9070 5550
rect 570 5530 600 5540
rect 650 5530 660 5540
rect 950 5530 960 5540
rect 1890 5530 1920 5540
rect 1930 5530 1940 5540
rect 2190 5530 2230 5540
rect 2420 5530 2480 5540
rect 2530 5530 2600 5540
rect 2940 5530 2960 5540
rect 3250 5530 3310 5540
rect 3650 5530 3660 5540
rect 5120 5530 5140 5540
rect 5250 5530 5260 5540
rect 5690 5530 5810 5540
rect 5850 5530 5910 5540
rect 6240 5530 6290 5540
rect 6470 5530 6550 5540
rect 6900 5530 6950 5540
rect 7380 5530 7530 5540
rect 7710 5530 7790 5540
rect 7960 5530 8030 5540
rect 8110 5530 8130 5540
rect 8180 5530 8230 5540
rect 8240 5530 8280 5540
rect 8760 5530 8770 5540
rect 8800 5530 8810 5540
rect 8840 5530 8860 5540
rect 8910 5530 8940 5540
rect 9000 5530 9070 5540
rect 1880 5520 1920 5530
rect 1930 5520 1940 5530
rect 2190 5520 2230 5530
rect 2420 5520 2470 5530
rect 2520 5520 2540 5530
rect 2550 5520 2560 5530
rect 2570 5520 2610 5530
rect 2950 5520 2970 5530
rect 3250 5520 3310 5530
rect 3500 5520 3510 5530
rect 3650 5520 3660 5530
rect 4170 5520 4190 5530
rect 5130 5520 5140 5530
rect 5740 5520 5920 5530
rect 6210 5520 6270 5530
rect 6480 5520 6550 5530
rect 6900 5520 6950 5530
rect 7380 5520 7510 5530
rect 7710 5520 7800 5530
rect 7950 5520 8030 5530
rect 8100 5520 8150 5530
rect 8170 5520 8190 5530
rect 8710 5520 8740 5530
rect 8750 5520 8760 5530
rect 8810 5520 8860 5530
rect 8910 5520 8940 5530
rect 9000 5520 9050 5530
rect 540 5510 570 5520
rect 580 5510 590 5520
rect 640 5510 650 5520
rect 1890 5510 1920 5520
rect 1930 5510 1960 5520
rect 2190 5510 2230 5520
rect 2410 5510 2470 5520
rect 2510 5510 2540 5520
rect 2550 5510 2600 5520
rect 3250 5510 3310 5520
rect 3520 5510 3540 5520
rect 5730 5510 5920 5520
rect 6210 5510 6260 5520
rect 6460 5510 6540 5520
rect 6900 5510 6940 5520
rect 7390 5510 7500 5520
rect 7710 5510 7800 5520
rect 7960 5510 8040 5520
rect 8100 5510 8150 5520
rect 8680 5510 8700 5520
rect 8720 5510 8750 5520
rect 8820 5510 8860 5520
rect 8920 5510 8940 5520
rect 9000 5510 9030 5520
rect 9110 5510 9130 5520
rect 490 5500 540 5510
rect 570 5500 590 5510
rect 620 5500 640 5510
rect 1890 5500 1920 5510
rect 1940 5500 1970 5510
rect 2190 5500 2230 5510
rect 2410 5500 2460 5510
rect 2480 5500 2590 5510
rect 2860 5500 2870 5510
rect 3240 5500 3320 5510
rect 3550 5500 3570 5510
rect 3710 5500 3720 5510
rect 3750 5500 3770 5510
rect 4160 5500 4170 5510
rect 5240 5500 5250 5510
rect 5730 5500 5930 5510
rect 6200 5500 6250 5510
rect 6370 5500 6510 5510
rect 6900 5500 6920 5510
rect 6930 5500 6950 5510
rect 7390 5500 7410 5510
rect 7420 5500 7500 5510
rect 7750 5500 7800 5510
rect 7960 5500 8040 5510
rect 8090 5500 8150 5510
rect 8160 5500 8170 5510
rect 8660 5500 8690 5510
rect 8730 5500 8740 5510
rect 8840 5500 8850 5510
rect 8920 5500 8950 5510
rect 9000 5500 9050 5510
rect 9120 5500 9130 5510
rect 420 5490 450 5500
rect 470 5490 540 5500
rect 570 5490 590 5500
rect 610 5490 640 5500
rect 1890 5490 1930 5500
rect 1940 5490 1970 5500
rect 2180 5490 2230 5500
rect 2400 5490 2590 5500
rect 3240 5490 3290 5500
rect 3300 5490 3320 5500
rect 3590 5490 3600 5500
rect 3610 5490 3630 5500
rect 3660 5490 3670 5500
rect 5110 5490 5130 5500
rect 5240 5490 5250 5500
rect 5730 5490 5760 5500
rect 5790 5490 5820 5500
rect 5840 5490 5930 5500
rect 6190 5490 6240 5500
rect 6350 5490 6460 5500
rect 7390 5490 7410 5500
rect 7420 5490 7500 5500
rect 7760 5490 7800 5500
rect 7960 5490 8150 5500
rect 8610 5490 8630 5500
rect 8650 5490 8690 5500
rect 8920 5490 8950 5500
rect 9000 5490 9040 5500
rect 430 5480 510 5490
rect 580 5480 590 5490
rect 610 5480 630 5490
rect 1900 5480 1970 5490
rect 2190 5480 2230 5490
rect 2400 5480 2490 5490
rect 2500 5480 2580 5490
rect 3240 5480 3290 5490
rect 3300 5480 3330 5490
rect 3550 5480 3580 5490
rect 3600 5480 3620 5490
rect 5760 5480 5790 5490
rect 5810 5480 5820 5490
rect 5840 5480 5920 5490
rect 6180 5480 6230 5490
rect 6350 5480 6450 5490
rect 7390 5480 7410 5490
rect 7420 5480 7500 5490
rect 7550 5480 7560 5490
rect 7750 5480 7800 5490
rect 7960 5480 8150 5490
rect 8600 5480 8620 5490
rect 8660 5480 8680 5490
rect 8930 5480 8940 5490
rect 9000 5480 9040 5490
rect 9120 5480 9130 5490
rect 460 5470 490 5480
rect 540 5470 550 5480
rect 580 5470 590 5480
rect 610 5470 620 5480
rect 1900 5470 1970 5480
rect 2180 5470 2230 5480
rect 2400 5470 2490 5480
rect 2510 5470 2530 5480
rect 2540 5470 2570 5480
rect 3240 5470 3290 5480
rect 3300 5470 3330 5480
rect 3560 5470 3570 5480
rect 3620 5470 3640 5480
rect 5110 5470 5120 5480
rect 5540 5470 5590 5480
rect 5620 5470 5800 5480
rect 5850 5470 5930 5480
rect 6180 5470 6240 5480
rect 6350 5470 6440 5480
rect 7400 5470 7500 5480
rect 7750 5470 7800 5480
rect 7960 5470 8150 5480
rect 8600 5470 8610 5480
rect 8660 5470 8680 5480
rect 8740 5470 8750 5480
rect 8930 5470 8940 5480
rect 9010 5470 9050 5480
rect 450 5460 460 5470
rect 540 5460 550 5470
rect 560 5460 590 5470
rect 1900 5460 1970 5470
rect 2190 5460 2230 5470
rect 2390 5460 2440 5470
rect 2460 5460 2470 5470
rect 2550 5460 2570 5470
rect 2910 5460 2930 5470
rect 3230 5460 3280 5470
rect 3300 5460 3330 5470
rect 3570 5460 3580 5470
rect 5110 5460 5120 5470
rect 5130 5460 5140 5470
rect 5520 5460 5540 5470
rect 5610 5460 5660 5470
rect 5750 5460 5930 5470
rect 6180 5460 6240 5470
rect 6360 5460 6440 5470
rect 7380 5460 7500 5470
rect 7730 5460 7810 5470
rect 7960 5460 8150 5470
rect 8520 5460 8530 5470
rect 8550 5460 8570 5470
rect 8590 5460 8610 5470
rect 8930 5460 8950 5470
rect 9010 5460 9070 5470
rect 450 5450 460 5460
rect 1900 5450 1970 5460
rect 2190 5450 2230 5460
rect 2430 5450 2460 5460
rect 2550 5450 2590 5460
rect 2850 5450 2910 5460
rect 3230 5450 3280 5460
rect 3300 5450 3320 5460
rect 3580 5450 3590 5460
rect 5110 5450 5140 5460
rect 5500 5450 5510 5460
rect 5570 5450 5590 5460
rect 5670 5450 5690 5460
rect 5770 5450 5920 5460
rect 6180 5450 6240 5460
rect 6250 5450 6270 5460
rect 6360 5450 6450 5460
rect 7390 5450 7510 5460
rect 7720 5450 7810 5460
rect 7960 5450 8150 5460
rect 8510 5450 8520 5460
rect 8570 5450 8610 5460
rect 8670 5450 8680 5460
rect 8930 5450 8950 5460
rect 9010 5450 9020 5460
rect 9030 5450 9070 5460
rect 9120 5450 9130 5460
rect 520 5440 530 5450
rect 580 5440 590 5450
rect 1910 5440 1930 5450
rect 1940 5440 1970 5450
rect 2190 5440 2220 5450
rect 2390 5440 2440 5450
rect 2540 5440 2550 5450
rect 2580 5440 2590 5450
rect 2600 5440 2630 5450
rect 2860 5440 2930 5450
rect 3230 5440 3270 5450
rect 3290 5440 3320 5450
rect 3580 5440 3590 5450
rect 5110 5440 5120 5450
rect 5480 5440 5490 5450
rect 5540 5440 5550 5450
rect 5680 5440 5710 5450
rect 5790 5440 5920 5450
rect 6180 5440 6240 5450
rect 6360 5440 6480 5450
rect 6920 5440 6940 5450
rect 7390 5440 7510 5450
rect 7720 5440 7810 5450
rect 7960 5440 8160 5450
rect 8500 5440 8510 5450
rect 8580 5440 8620 5450
rect 8670 5440 8680 5450
rect 8940 5440 8960 5450
rect 9020 5440 9030 5450
rect 9040 5440 9060 5450
rect 510 5430 520 5440
rect 1910 5430 1970 5440
rect 2190 5430 2230 5440
rect 2390 5430 2430 5440
rect 2580 5430 2600 5440
rect 2640 5430 2650 5440
rect 2860 5430 2950 5440
rect 3000 5430 3020 5440
rect 3220 5430 3270 5440
rect 3290 5430 3300 5440
rect 5110 5430 5120 5440
rect 5470 5430 5480 5440
rect 5520 5430 5530 5440
rect 5640 5430 5740 5440
rect 5800 5430 5920 5440
rect 6180 5430 6230 5440
rect 6480 5430 6510 5440
rect 6920 5430 6940 5440
rect 7390 5430 7470 5440
rect 7480 5430 7510 5440
rect 7630 5430 7640 5440
rect 7790 5430 7810 5440
rect 7960 5430 7990 5440
rect 8010 5430 8160 5440
rect 8430 5430 8450 5440
rect 8490 5430 8510 5440
rect 8590 5430 8620 5440
rect 8940 5430 8970 5440
rect 9110 5430 9120 5440
rect 9550 5430 9570 5440
rect 450 5420 460 5430
rect 500 5420 510 5430
rect 1920 5420 1970 5430
rect 2200 5420 2230 5430
rect 2390 5420 2420 5430
rect 2520 5420 2530 5430
rect 2610 5420 2660 5430
rect 2860 5420 3030 5430
rect 3200 5420 3280 5430
rect 5230 5420 5240 5430
rect 5460 5420 5470 5430
rect 5500 5420 5510 5430
rect 5550 5420 5580 5430
rect 5700 5420 5740 5430
rect 5840 5420 5920 5430
rect 6180 5420 6230 5430
rect 6530 5420 6540 5430
rect 6930 5420 6940 5430
rect 7390 5420 7470 5430
rect 7480 5420 7510 5430
rect 7630 5420 7640 5430
rect 7790 5420 7820 5430
rect 7850 5420 7860 5430
rect 7870 5420 7880 5430
rect 7960 5420 7980 5430
rect 8010 5420 8150 5430
rect 8470 5420 8510 5430
rect 8600 5420 8620 5430
rect 8940 5420 8980 5430
rect 9100 5420 9120 5430
rect 570 5410 580 5420
rect 1920 5410 1970 5420
rect 2200 5410 2220 5420
rect 2390 5410 2420 5420
rect 2520 5410 2530 5420
rect 2600 5410 2660 5420
rect 2720 5410 2730 5420
rect 2860 5410 2920 5420
rect 2960 5410 3040 5420
rect 3200 5410 3270 5420
rect 3570 5410 3580 5420
rect 5230 5410 5240 5420
rect 5450 5410 5460 5420
rect 5490 5410 5500 5420
rect 5530 5410 5540 5420
rect 5730 5410 5750 5420
rect 5860 5410 5920 5420
rect 6180 5410 6220 5420
rect 6410 5410 6430 5420
rect 6560 5410 6600 5420
rect 7400 5410 7520 5420
rect 7630 5410 7640 5420
rect 7790 5410 7880 5420
rect 7950 5410 8160 5420
rect 8480 5410 8510 5420
rect 8610 5410 8620 5420
rect 8940 5410 8990 5420
rect 9090 5410 9100 5420
rect 9480 5410 9500 5420
rect 9540 5410 9550 5420
rect 9580 5410 9590 5420
rect 430 5400 440 5410
rect 770 5400 780 5410
rect 830 5400 840 5410
rect 890 5400 910 5410
rect 920 5400 950 5410
rect 1920 5400 1980 5410
rect 2200 5400 2220 5410
rect 2390 5400 2420 5410
rect 2580 5400 2660 5410
rect 2720 5400 2730 5410
rect 2870 5400 2910 5410
rect 2990 5400 3050 5410
rect 3160 5400 3230 5410
rect 3570 5400 3580 5410
rect 5100 5400 5110 5410
rect 5440 5400 5450 5410
rect 5470 5400 5490 5410
rect 5870 5400 5920 5410
rect 6180 5400 6210 5410
rect 6600 5400 6620 5410
rect 7400 5400 7520 5410
rect 7780 5400 7890 5410
rect 7960 5400 8150 5410
rect 8340 5400 8350 5410
rect 8490 5400 8510 5410
rect 8830 5400 8840 5410
rect 8950 5400 9000 5410
rect 9070 5400 9080 5410
rect 9540 5400 9550 5410
rect 410 5390 420 5400
rect 760 5390 770 5400
rect 820 5390 830 5400
rect 980 5390 990 5400
rect 1920 5390 1990 5400
rect 2200 5390 2220 5400
rect 2380 5390 2420 5400
rect 2580 5390 2610 5400
rect 2620 5390 2680 5400
rect 2760 5390 2790 5400
rect 2890 5390 2930 5400
rect 3050 5390 3090 5400
rect 3130 5390 3210 5400
rect 3570 5390 3580 5400
rect 5430 5390 5440 5400
rect 5460 5390 5490 5400
rect 5880 5390 5910 5400
rect 6180 5390 6210 5400
rect 6620 5390 6640 5400
rect 7410 5390 7520 5400
rect 7750 5390 7890 5400
rect 7900 5390 7910 5400
rect 7960 5390 8140 5400
rect 8310 5390 8320 5400
rect 8340 5390 8350 5400
rect 8500 5390 8520 5400
rect 8840 5390 8860 5400
rect 8950 5390 8960 5400
rect 8980 5390 9050 5400
rect 9530 5390 9540 5400
rect 390 5380 400 5390
rect 460 5380 470 5390
rect 1920 5380 1990 5390
rect 2200 5380 2220 5390
rect 2380 5380 2430 5390
rect 2480 5380 2490 5390
rect 2580 5380 2610 5390
rect 2640 5380 2690 5390
rect 2740 5380 2840 5390
rect 2870 5380 2880 5390
rect 2900 5380 2910 5390
rect 2920 5380 2950 5390
rect 3080 5380 3190 5390
rect 5090 5380 5100 5390
rect 5410 5380 5450 5390
rect 5460 5380 5480 5390
rect 5880 5380 5920 5390
rect 6180 5380 6210 5390
rect 6630 5380 6670 5390
rect 7410 5380 7520 5390
rect 7720 5380 7890 5390
rect 7960 5380 8180 5390
rect 8240 5380 8350 5390
rect 8400 5380 8450 5390
rect 8500 5380 8520 5390
rect 8840 5380 8880 5390
rect 9400 5380 9410 5390
rect 9480 5380 9490 5390
rect 370 5370 380 5380
rect 560 5370 570 5380
rect 880 5370 920 5380
rect 1920 5370 1990 5380
rect 2380 5370 2420 5380
rect 2480 5370 2490 5380
rect 2580 5370 2610 5380
rect 2680 5370 2710 5380
rect 2720 5370 2740 5380
rect 2750 5370 2880 5380
rect 2940 5370 3000 5380
rect 3110 5370 3170 5380
rect 3490 5370 3510 5380
rect 5090 5370 5100 5380
rect 5130 5370 5140 5380
rect 5440 5370 5460 5380
rect 5720 5370 5750 5380
rect 5870 5370 5910 5380
rect 6180 5370 6200 5380
rect 6650 5370 6670 5380
rect 7410 5370 7510 5380
rect 7650 5370 7790 5380
rect 7820 5370 7900 5380
rect 7970 5370 8180 5380
rect 8220 5370 8230 5380
rect 8280 5370 8350 5380
rect 8400 5370 8440 5380
rect 8500 5370 8530 5380
rect 8840 5370 8880 5380
rect 8940 5370 8950 5380
rect 9400 5370 9410 5380
rect 9440 5370 9450 5380
rect 9490 5370 9500 5380
rect 350 5360 360 5370
rect 440 5360 450 5370
rect 540 5360 550 5370
rect 880 5360 900 5370
rect 1930 5360 1990 5370
rect 2390 5360 2420 5370
rect 2480 5360 2490 5370
rect 2590 5360 2610 5370
rect 2710 5360 2910 5370
rect 2930 5360 3010 5370
rect 3490 5360 3520 5370
rect 5090 5360 5100 5370
rect 5130 5360 5140 5370
rect 5430 5360 5440 5370
rect 5750 5360 5760 5370
rect 5820 5360 5900 5370
rect 6180 5360 6200 5370
rect 6550 5360 6560 5370
rect 6660 5360 6680 5370
rect 7420 5360 7520 5370
rect 7640 5360 7780 5370
rect 7830 5360 7920 5370
rect 7970 5360 8180 5370
rect 8210 5360 8230 5370
rect 8280 5360 8350 5370
rect 8400 5360 8440 5370
rect 8490 5360 8530 5370
rect 8840 5360 8870 5370
rect 8880 5360 8910 5370
rect 8930 5360 8940 5370
rect 9290 5360 9310 5370
rect 9350 5360 9360 5370
rect 9400 5360 9410 5370
rect 9500 5360 9510 5370
rect 9570 5360 9580 5370
rect 330 5350 350 5360
rect 400 5350 440 5360
rect 880 5350 900 5360
rect 1930 5350 2000 5360
rect 2390 5350 2420 5360
rect 2460 5350 2510 5360
rect 2600 5350 2620 5360
rect 2720 5350 3020 5360
rect 3490 5350 3520 5360
rect 3560 5350 3570 5360
rect 5090 5350 5100 5360
rect 5220 5350 5230 5360
rect 5410 5350 5430 5360
rect 5460 5350 5470 5360
rect 5550 5350 5570 5360
rect 5580 5350 5590 5360
rect 5600 5350 5650 5360
rect 5710 5350 5750 5360
rect 5830 5350 5860 5360
rect 6180 5350 6200 5360
rect 6370 5350 6390 5360
rect 6540 5350 6570 5360
rect 6680 5350 6700 5360
rect 7400 5350 7520 5360
rect 7580 5350 7760 5360
rect 7840 5350 7900 5360
rect 7970 5350 8140 5360
rect 8150 5350 8180 5360
rect 8200 5350 8230 5360
rect 8290 5350 8350 5360
rect 8400 5350 8420 5360
rect 8490 5350 8530 5360
rect 8770 5350 8780 5360
rect 8840 5350 8850 5360
rect 9270 5350 9280 5360
rect 9400 5350 9410 5360
rect 9510 5350 9520 5360
rect 9570 5350 9580 5360
rect 300 5340 330 5350
rect 360 5340 380 5350
rect 1930 5340 2000 5350
rect 2390 5340 2420 5350
rect 2460 5340 2520 5350
rect 2610 5340 2620 5350
rect 2720 5340 3030 5350
rect 3490 5340 3510 5350
rect 5140 5340 5150 5350
rect 5220 5340 5230 5350
rect 5400 5340 5420 5350
rect 5590 5340 5620 5350
rect 5670 5340 5750 5350
rect 5840 5340 5850 5350
rect 6200 5340 6210 5350
rect 6280 5340 6300 5350
rect 6360 5340 6380 5350
rect 6540 5340 6570 5350
rect 6690 5340 6710 5350
rect 7370 5340 7530 5350
rect 7570 5340 7720 5350
rect 7740 5340 7750 5350
rect 7840 5340 7900 5350
rect 7970 5340 8130 5350
rect 8170 5340 8220 5350
rect 8300 5340 8360 5350
rect 8510 5340 8530 5350
rect 8600 5340 8610 5350
rect 8690 5340 8700 5350
rect 8770 5340 8800 5350
rect 8840 5340 8850 5350
rect 9520 5340 9530 5350
rect 270 5330 290 5340
rect 320 5330 330 5340
rect 560 5330 570 5340
rect 1930 5330 2000 5340
rect 2390 5330 2420 5340
rect 2450 5330 2480 5340
rect 2520 5330 2530 5340
rect 2590 5330 2600 5340
rect 2720 5330 3050 5340
rect 3480 5330 3500 5340
rect 5090 5330 5110 5340
rect 5140 5330 5160 5340
rect 5220 5330 5230 5340
rect 5700 5330 5770 5340
rect 5850 5330 5860 5340
rect 6190 5330 6210 5340
rect 6250 5330 6290 5340
rect 6350 5330 6370 5340
rect 6690 5330 6720 5340
rect 7360 5330 7480 5340
rect 7490 5330 7730 5340
rect 7840 5330 7900 5340
rect 7980 5330 8080 5340
rect 8100 5330 8110 5340
rect 8170 5330 8220 5340
rect 8300 5330 8360 5340
rect 8510 5330 8530 5340
rect 8590 5330 8610 5340
rect 8770 5330 8830 5340
rect 9410 5330 9420 5340
rect 9520 5330 9530 5340
rect 9580 5330 9590 5340
rect 250 5320 270 5330
rect 570 5320 580 5330
rect 1930 5320 2000 5330
rect 2390 5320 2430 5330
rect 2440 5320 2480 5330
rect 2520 5320 2540 5330
rect 2590 5320 2600 5330
rect 2650 5320 2660 5330
rect 2730 5320 2790 5330
rect 2800 5320 3050 5330
rect 5130 5320 5150 5330
rect 5160 5320 5170 5330
rect 5210 5320 5220 5330
rect 5750 5320 5840 5330
rect 5850 5320 5860 5330
rect 6190 5320 6220 5330
rect 6240 5320 6290 5330
rect 6340 5320 6400 5330
rect 6700 5320 6730 5330
rect 7360 5320 7700 5330
rect 7840 5320 7890 5330
rect 7980 5320 8060 5330
rect 8180 5320 8220 5330
rect 8310 5320 8360 5330
rect 8460 5320 8490 5330
rect 8520 5320 8530 5330
rect 8590 5320 8620 5330
rect 8710 5320 8720 5330
rect 8770 5320 8790 5330
rect 9310 5320 9330 5330
rect 9520 5320 9530 5330
rect 9590 5320 9600 5330
rect 240 5310 290 5320
rect 580 5310 590 5320
rect 1940 5310 2000 5320
rect 2390 5310 2470 5320
rect 2530 5310 2550 5320
rect 2590 5310 2600 5320
rect 2630 5310 2680 5320
rect 2740 5310 2810 5320
rect 2830 5310 3050 5320
rect 5160 5310 5170 5320
rect 5180 5310 5190 5320
rect 5200 5310 5220 5320
rect 5770 5310 5790 5320
rect 5800 5310 5810 5320
rect 6200 5310 6280 5320
rect 6370 5310 6460 5320
rect 6490 5310 6510 5320
rect 6560 5310 6590 5320
rect 6640 5310 6660 5320
rect 6720 5310 6740 5320
rect 7360 5310 7640 5320
rect 7650 5310 7670 5320
rect 7690 5310 7700 5320
rect 7830 5310 7900 5320
rect 7980 5310 8010 5320
rect 8030 5310 8060 5320
rect 8180 5310 8220 5320
rect 8310 5310 8370 5320
rect 8520 5310 8540 5320
rect 8590 5310 8630 5320
rect 8700 5310 8740 5320
rect 8750 5310 8790 5320
rect 9120 5310 9130 5320
rect 9250 5310 9260 5320
rect 9310 5310 9320 5320
rect 230 5300 240 5310
rect 570 5300 580 5310
rect 1940 5300 2010 5310
rect 2390 5300 2460 5310
rect 2530 5300 2570 5310
rect 2590 5300 2600 5310
rect 2630 5300 2660 5310
rect 2740 5300 3060 5310
rect 5150 5300 5170 5310
rect 5180 5300 5190 5310
rect 5200 5300 5210 5310
rect 6200 5300 6290 5310
rect 6350 5300 6390 5310
rect 6400 5300 6430 5310
rect 6480 5300 6540 5310
rect 6680 5300 6690 5310
rect 6730 5300 6770 5310
rect 7350 5300 7690 5310
rect 7840 5300 7910 5310
rect 7980 5300 8000 5310
rect 8180 5300 8200 5310
rect 8320 5300 8370 5310
rect 8480 5300 8490 5310
rect 8530 5300 8540 5310
rect 8590 5300 8640 5310
rect 8690 5300 8730 5310
rect 8770 5300 8780 5310
rect 9250 5300 9260 5310
rect 9300 5300 9330 5310
rect 9360 5300 9370 5310
rect 9420 5300 9430 5310
rect 210 5290 230 5300
rect 1940 5290 2010 5300
rect 2400 5290 2460 5300
rect 2570 5290 2580 5300
rect 2590 5290 2600 5300
rect 2610 5290 2630 5300
rect 2640 5290 2660 5300
rect 2760 5290 2840 5300
rect 2860 5290 2990 5300
rect 5150 5290 5160 5300
rect 5180 5290 5190 5300
rect 5200 5290 5210 5300
rect 6210 5290 6320 5300
rect 6330 5290 6380 5300
rect 6400 5290 6460 5300
rect 6480 5290 6490 5300
rect 6700 5290 6720 5300
rect 6740 5290 6770 5300
rect 7340 5290 7640 5300
rect 7680 5290 7690 5300
rect 7840 5290 7910 5300
rect 7990 5290 8000 5300
rect 8200 5290 8210 5300
rect 8320 5290 8370 5300
rect 8490 5290 8500 5300
rect 8530 5290 8550 5300
rect 8590 5290 8640 5300
rect 9110 5290 9120 5300
rect 9250 5290 9260 5300
rect 9510 5290 9520 5300
rect 9560 5290 9570 5300
rect 9940 5290 9950 5300
rect 9970 5290 9980 5300
rect 600 5280 610 5290
rect 1940 5280 2010 5290
rect 2400 5280 2460 5290
rect 2580 5280 2640 5290
rect 2800 5280 2970 5290
rect 5110 5280 5120 5290
rect 5140 5280 5150 5290
rect 5200 5280 5220 5290
rect 6220 5280 6290 5290
rect 6300 5280 6380 5290
rect 6740 5280 6760 5290
rect 7330 5280 7570 5290
rect 7580 5280 7620 5290
rect 7650 5280 7660 5290
rect 7830 5280 7910 5290
rect 8190 5280 8200 5290
rect 8330 5280 8370 5290
rect 8430 5280 8440 5290
rect 8530 5280 8550 5290
rect 8590 5280 8610 5290
rect 8650 5280 8660 5290
rect 9030 5280 9040 5290
rect 9070 5280 9080 5290
rect 9100 5280 9120 5290
rect 9260 5280 9270 5290
rect 9510 5280 9520 5290
rect 9580 5280 9590 5290
rect 9940 5280 9950 5290
rect 610 5270 630 5280
rect 1400 5270 1410 5280
rect 1950 5270 2010 5280
rect 2410 5270 2450 5280
rect 2590 5270 2650 5280
rect 2810 5270 2970 5280
rect 5190 5270 5200 5280
rect 6310 5270 6330 5280
rect 7330 5270 7570 5280
rect 7600 5270 7610 5280
rect 7670 5270 7680 5280
rect 7840 5270 7910 5280
rect 8190 5270 8200 5280
rect 8330 5270 8370 5280
rect 8420 5270 8450 5280
rect 8510 5270 8520 5280
rect 8550 5270 8560 5280
rect 8590 5270 8610 5280
rect 9020 5270 9040 5280
rect 9100 5270 9130 5280
rect 9270 5270 9280 5280
rect 9390 5270 9400 5280
rect 9510 5270 9520 5280
rect 9940 5270 9950 5280
rect 730 5260 740 5270
rect 1390 5260 1400 5270
rect 1950 5260 2020 5270
rect 2410 5260 2440 5270
rect 2600 5260 2610 5270
rect 2630 5260 2650 5270
rect 2730 5260 2750 5270
rect 2820 5260 2860 5270
rect 2870 5260 2910 5270
rect 2920 5260 2960 5270
rect 3490 5260 3500 5270
rect 5080 5260 5100 5270
rect 5180 5260 5210 5270
rect 6300 5260 6330 5270
rect 7340 5260 7430 5270
rect 7440 5260 7470 5270
rect 7480 5260 7500 5270
rect 7510 5260 7550 5270
rect 7600 5260 7610 5270
rect 7620 5260 7630 5270
rect 7650 5260 7660 5270
rect 7850 5260 7940 5270
rect 8190 5260 8200 5270
rect 8340 5260 8370 5270
rect 8420 5260 8450 5270
rect 8960 5260 8970 5270
rect 9030 5260 9040 5270
rect 9100 5260 9130 5270
rect 9170 5260 9180 5270
rect 9350 5260 9360 5270
rect 9430 5260 9440 5270
rect 9470 5260 9480 5270
rect 9540 5260 9550 5270
rect 9940 5260 9950 5270
rect 9980 5260 9990 5270
rect 350 5250 360 5260
rect 610 5250 620 5260
rect 1380 5250 1390 5260
rect 1950 5250 2020 5260
rect 2610 5250 2620 5260
rect 2640 5250 2650 5260
rect 2730 5250 2740 5260
rect 2820 5250 2850 5260
rect 2890 5250 2910 5260
rect 3500 5250 3510 5260
rect 5090 5250 5100 5260
rect 5180 5250 5190 5260
rect 5730 5250 5750 5260
rect 6340 5250 6370 5260
rect 7340 5250 7450 5260
rect 7460 5250 7480 5260
rect 7490 5250 7500 5260
rect 7580 5250 7600 5260
rect 7610 5250 7630 5260
rect 7650 5250 7680 5260
rect 7850 5250 7860 5260
rect 7870 5250 7930 5260
rect 8190 5250 8220 5260
rect 8340 5250 8370 5260
rect 8430 5250 8470 5260
rect 8920 5250 8940 5260
rect 8970 5250 8980 5260
rect 9030 5250 9040 5260
rect 9110 5250 9130 5260
rect 9350 5250 9360 5260
rect 9760 5250 9790 5260
rect 620 5240 630 5250
rect 1370 5240 1380 5250
rect 1950 5240 2020 5250
rect 2620 5240 2630 5250
rect 2830 5240 2840 5250
rect 2890 5240 2920 5250
rect 3500 5240 3510 5250
rect 5080 5240 5120 5250
rect 5700 5240 5750 5250
rect 6370 5240 6380 5250
rect 6390 5240 6410 5250
rect 6420 5240 6430 5250
rect 7330 5240 7440 5250
rect 7580 5240 7600 5250
rect 7610 5240 7630 5250
rect 7640 5240 7680 5250
rect 7850 5240 7860 5250
rect 7870 5240 7940 5250
rect 8190 5240 8220 5250
rect 8350 5240 8380 5250
rect 8430 5240 8490 5250
rect 8500 5240 8510 5250
rect 8840 5240 8850 5250
rect 8890 5240 8900 5250
rect 8910 5240 8930 5250
rect 9030 5240 9040 5250
rect 9120 5240 9140 5250
rect 9300 5240 9310 5250
rect 9350 5240 9360 5250
rect 9440 5240 9450 5250
rect 9950 5240 9960 5250
rect 620 5230 630 5240
rect 1360 5230 1370 5240
rect 1950 5230 2030 5240
rect 2640 5230 2650 5240
rect 2810 5230 2830 5240
rect 2900 5230 2930 5240
rect 3500 5230 3510 5240
rect 6380 5230 6450 5240
rect 6460 5230 6480 5240
rect 6540 5230 6560 5240
rect 7340 5230 7450 5240
rect 7540 5230 7550 5240
rect 7580 5230 7590 5240
rect 7640 5230 7660 5240
rect 7670 5230 7680 5240
rect 7860 5230 7930 5240
rect 8190 5230 8220 5240
rect 8350 5230 8370 5240
rect 8830 5230 8840 5240
rect 8860 5230 8890 5240
rect 8900 5230 8930 5240
rect 9040 5230 9050 5240
rect 9720 5230 9730 5240
rect 1950 5220 2030 5230
rect 2720 5220 2730 5230
rect 2810 5220 2820 5230
rect 2900 5220 2950 5230
rect 5070 5220 5110 5230
rect 5130 5220 5140 5230
rect 6390 5220 6550 5230
rect 7340 5220 7420 5230
rect 7430 5220 7440 5230
rect 7450 5220 7460 5230
rect 7520 5220 7550 5230
rect 7560 5220 7600 5230
rect 7620 5220 7640 5230
rect 7650 5220 7660 5230
rect 7670 5220 7680 5230
rect 7850 5220 7930 5230
rect 8190 5220 8200 5230
rect 8360 5220 8380 5230
rect 8870 5220 8930 5230
rect 8990 5220 9000 5230
rect 9040 5220 9050 5230
rect 9850 5220 9860 5230
rect 9940 5220 9950 5230
rect 9990 5220 9990 5230
rect 1960 5210 2030 5220
rect 2710 5210 2720 5220
rect 2910 5210 2960 5220
rect 5080 5210 5110 5220
rect 5120 5210 5140 5220
rect 6470 5210 6480 5220
rect 7340 5210 7420 5220
rect 7430 5210 7440 5220
rect 7530 5210 7600 5220
rect 7610 5210 7640 5220
rect 7650 5210 7670 5220
rect 7860 5210 7940 5220
rect 8190 5210 8200 5220
rect 8290 5210 8300 5220
rect 8360 5210 8380 5220
rect 8750 5210 8780 5220
rect 8820 5210 8830 5220
rect 8870 5210 8880 5220
rect 8900 5210 8930 5220
rect 9040 5210 9050 5220
rect 9180 5210 9190 5220
rect 9290 5210 9300 5220
rect 9370 5210 9380 5220
rect 9830 5210 9840 5220
rect 9990 5210 9990 5220
rect 680 5200 690 5210
rect 1960 5200 2030 5210
rect 2670 5200 2680 5210
rect 2910 5200 3000 5210
rect 5080 5200 5100 5210
rect 5130 5200 5140 5210
rect 5160 5200 5170 5210
rect 7350 5200 7440 5210
rect 7530 5200 7540 5210
rect 7550 5200 7620 5210
rect 7630 5200 7640 5210
rect 7650 5200 7660 5210
rect 7860 5200 7950 5210
rect 8010 5200 8020 5210
rect 8190 5200 8200 5210
rect 8270 5200 8310 5210
rect 8350 5200 8360 5210
rect 8780 5200 8790 5210
rect 8810 5200 8830 5210
rect 8870 5200 8890 5210
rect 8910 5200 8930 5210
rect 9050 5200 9060 5210
rect 9100 5200 9110 5210
rect 9310 5200 9320 5210
rect 9350 5200 9360 5210
rect 9790 5200 9800 5210
rect 9830 5200 9840 5210
rect 9860 5200 9870 5210
rect 9910 5200 9920 5210
rect 690 5190 700 5200
rect 1830 5190 1840 5200
rect 1960 5190 2030 5200
rect 2680 5190 2690 5200
rect 2730 5190 2740 5200
rect 2910 5190 3010 5200
rect 3350 5190 3360 5200
rect 3480 5190 3490 5200
rect 5080 5190 5100 5200
rect 5130 5190 5140 5200
rect 5160 5190 5170 5200
rect 7350 5190 7440 5200
rect 7540 5190 7550 5200
rect 7560 5190 7590 5200
rect 7610 5190 7670 5200
rect 7860 5190 7950 5200
rect 8010 5190 8030 5200
rect 8270 5190 8330 5200
rect 8680 5190 8690 5200
rect 8720 5190 8730 5200
rect 8740 5190 8750 5200
rect 8790 5190 8810 5200
rect 8820 5190 8840 5200
rect 8900 5190 8930 5200
rect 9040 5190 9060 5200
rect 9110 5190 9130 5200
rect 9550 5190 9560 5200
rect 9590 5190 9600 5200
rect 9790 5190 9800 5200
rect 620 5180 630 5190
rect 670 5180 710 5190
rect 1810 5180 1850 5190
rect 1960 5180 2040 5190
rect 2740 5180 2750 5190
rect 2910 5180 2940 5190
rect 2990 5180 3020 5190
rect 5070 5180 5080 5190
rect 5090 5180 5170 5190
rect 7350 5180 7440 5190
rect 7540 5180 7600 5190
rect 7610 5180 7630 5190
rect 7870 5180 7960 5190
rect 8010 5180 8030 5190
rect 8260 5180 8270 5190
rect 8650 5180 8660 5190
rect 8730 5180 8750 5190
rect 8790 5180 8840 5190
rect 8900 5180 8910 5190
rect 8920 5180 8930 5190
rect 9050 5180 9060 5190
rect 9100 5180 9110 5190
rect 9130 5180 9140 5190
rect 9900 5180 9910 5190
rect 9940 5180 9950 5190
rect 620 5170 630 5180
rect 680 5170 700 5180
rect 1800 5170 1860 5180
rect 1960 5170 2040 5180
rect 2700 5170 2720 5180
rect 2910 5170 2930 5180
rect 2990 5170 3010 5180
rect 3330 5170 3340 5180
rect 3470 5170 3480 5180
rect 5110 5170 5170 5180
rect 7340 5170 7440 5180
rect 7540 5170 7590 5180
rect 7680 5170 7690 5180
rect 7870 5170 7950 5180
rect 8010 5170 8030 5180
rect 8100 5170 8110 5180
rect 8190 5170 8230 5180
rect 8250 5170 8260 5180
rect 8620 5170 8630 5180
rect 8730 5170 8750 5180
rect 8790 5170 8800 5180
rect 8820 5170 8840 5180
rect 8880 5170 8890 5180
rect 8910 5170 8930 5180
rect 8970 5170 8980 5180
rect 9020 5170 9030 5180
rect 9060 5170 9070 5180
rect 9100 5170 9110 5180
rect 9750 5170 9760 5180
rect 9800 5170 9810 5180
rect 9870 5170 9880 5180
rect 620 5160 630 5170
rect 640 5160 650 5170
rect 690 5160 710 5170
rect 1800 5160 1860 5170
rect 1960 5160 2040 5170
rect 2720 5160 2730 5170
rect 2790 5160 2800 5170
rect 2900 5160 2920 5170
rect 2990 5160 3010 5170
rect 5080 5160 5090 5170
rect 5100 5160 5130 5170
rect 5140 5160 5170 5170
rect 7330 5160 7450 5170
rect 7550 5160 7560 5170
rect 7890 5160 7960 5170
rect 8010 5160 8030 5170
rect 8100 5160 8120 5170
rect 8190 5160 8230 5170
rect 8710 5160 8720 5170
rect 8740 5160 8760 5170
rect 8910 5160 8930 5170
rect 9060 5160 9070 5170
rect 9440 5160 9450 5170
rect 9460 5160 9470 5170
rect 9840 5160 9850 5170
rect 9910 5160 9920 5170
rect 640 5150 660 5160
rect 680 5150 720 5160
rect 1790 5150 1830 5160
rect 1850 5150 1860 5160
rect 1960 5150 2050 5160
rect 2730 5150 2740 5160
rect 2900 5150 2920 5160
rect 3000 5150 3010 5160
rect 5090 5150 5130 5160
rect 5140 5150 5160 5160
rect 7340 5150 7450 5160
rect 7890 5150 7960 5160
rect 8010 5150 8040 5160
rect 8100 5150 8140 5160
rect 8180 5150 8230 5160
rect 8600 5150 8610 5160
rect 8690 5150 8700 5160
rect 8740 5150 8760 5160
rect 8910 5150 8930 5160
rect 9400 5150 9410 5160
rect 9470 5150 9480 5160
rect 9500 5150 9510 5160
rect 9580 5150 9590 5160
rect 9980 5150 9990 5160
rect 610 5140 620 5150
rect 640 5140 740 5150
rect 1800 5140 1840 5150
rect 1960 5140 2040 5150
rect 2740 5140 2750 5150
rect 2890 5140 2910 5150
rect 2990 5140 3040 5150
rect 3450 5140 3460 5150
rect 5110 5140 5120 5150
rect 5140 5140 5150 5150
rect 5180 5140 5190 5150
rect 7340 5140 7450 5150
rect 7570 5140 7610 5150
rect 7620 5140 7640 5150
rect 7880 5140 7970 5150
rect 8000 5140 8040 5150
rect 8100 5140 8170 5150
rect 8180 5140 8210 5150
rect 8600 5140 8620 5150
rect 8690 5140 8700 5150
rect 8740 5140 8760 5150
rect 8900 5140 8930 5150
rect 9040 5140 9050 5150
rect 9370 5140 9380 5150
rect 9470 5140 9480 5150
rect 9500 5140 9510 5150
rect 9580 5140 9590 5150
rect 130 5130 140 5140
rect 610 5130 620 5140
rect 650 5130 740 5140
rect 1800 5130 1840 5140
rect 1970 5130 2060 5140
rect 2750 5130 2760 5140
rect 2830 5130 2840 5140
rect 2890 5130 2910 5140
rect 2980 5130 3040 5140
rect 5140 5130 5150 5140
rect 5170 5130 5190 5140
rect 7330 5130 7450 5140
rect 7560 5130 7590 5140
rect 7610 5130 7640 5140
rect 7880 5130 7970 5140
rect 8010 5130 8050 5140
rect 8090 5130 8200 5140
rect 8470 5130 8480 5140
rect 8650 5130 8660 5140
rect 8690 5130 8700 5140
rect 8750 5130 8760 5140
rect 8820 5130 8830 5140
rect 8890 5130 8900 5140
rect 8910 5130 8930 5140
rect 8990 5130 9010 5140
rect 9040 5130 9050 5140
rect 9460 5130 9470 5140
rect 9500 5130 9510 5140
rect 9720 5130 9730 5140
rect 9760 5130 9770 5140
rect 9920 5130 9930 5140
rect 580 5120 590 5130
rect 610 5120 620 5130
rect 660 5120 740 5130
rect 1800 5120 1880 5130
rect 1890 5120 1900 5130
rect 1970 5120 2060 5130
rect 2770 5120 2780 5130
rect 2860 5120 2910 5130
rect 2960 5120 3000 5130
rect 3010 5120 3030 5130
rect 3310 5120 3320 5130
rect 5120 5120 5140 5130
rect 5180 5120 5200 5130
rect 7330 5120 7450 5130
rect 7520 5120 7530 5130
rect 7580 5120 7590 5130
rect 7600 5120 7620 5130
rect 7630 5120 7640 5130
rect 7870 5120 7970 5130
rect 8010 5120 8080 5130
rect 8090 5120 8130 5130
rect 8140 5120 8220 5130
rect 8430 5120 8440 5130
rect 8650 5120 8660 5130
rect 8760 5120 8770 5130
rect 8800 5120 8810 5130
rect 8850 5120 8860 5130
rect 8890 5120 8900 5130
rect 8910 5120 8920 5130
rect 9010 5120 9020 5130
rect 9280 5120 9290 5130
rect 9360 5120 9370 5130
rect 9590 5120 9600 5130
rect 9720 5120 9730 5130
rect 9890 5120 9900 5130
rect 580 5110 600 5120
rect 620 5110 630 5120
rect 670 5110 740 5120
rect 1780 5110 1860 5120
rect 1890 5110 1900 5120
rect 1970 5110 2070 5120
rect 2780 5110 2800 5120
rect 2900 5110 2910 5120
rect 2960 5110 2990 5120
rect 3000 5110 3030 5120
rect 3430 5110 3440 5120
rect 5180 5110 5200 5120
rect 7320 5110 7450 5120
rect 7870 5110 7970 5120
rect 8010 5110 8030 5120
rect 8110 5110 8220 5120
rect 8510 5110 8520 5120
rect 8650 5110 8660 5120
rect 8850 5110 8860 5120
rect 8900 5110 8910 5120
rect 8920 5110 8930 5120
rect 9250 5110 9260 5120
rect 9360 5110 9370 5120
rect 9510 5110 9520 5120
rect 580 5100 630 5110
rect 670 5100 750 5110
rect 1800 5100 1860 5110
rect 1970 5100 2080 5110
rect 2810 5100 2820 5110
rect 2930 5100 2940 5110
rect 2970 5100 2990 5110
rect 3000 5100 3030 5110
rect 3460 5100 3470 5110
rect 5170 5100 5180 5110
rect 5190 5100 5200 5110
rect 7310 5100 7450 5110
rect 7460 5100 7470 5110
rect 7540 5100 7550 5110
rect 7560 5100 7570 5110
rect 7880 5100 7970 5110
rect 8010 5100 8030 5110
rect 8110 5100 8210 5110
rect 8410 5100 8420 5110
rect 8490 5100 8500 5110
rect 8660 5100 8670 5110
rect 9550 5100 9560 5110
rect 9730 5100 9740 5110
rect 540 5090 550 5100
rect 580 5090 630 5100
rect 680 5090 750 5100
rect 1800 5090 1860 5100
rect 1880 5090 1890 5100
rect 1980 5090 2090 5100
rect 2830 5090 2850 5100
rect 2960 5090 2980 5100
rect 3010 5090 3030 5100
rect 5170 5090 5180 5100
rect 5190 5090 5210 5100
rect 7320 5090 7450 5100
rect 7880 5090 7980 5100
rect 8010 5090 8040 5100
rect 8130 5090 8170 5100
rect 8180 5090 8210 5100
rect 8220 5090 8230 5100
rect 8320 5090 8330 5100
rect 8370 5090 8380 5100
rect 8400 5090 8420 5100
rect 8460 5090 8470 5100
rect 8660 5090 8670 5100
rect 8700 5090 8710 5100
rect 8770 5090 8780 5100
rect 8810 5090 8820 5100
rect 8860 5090 8870 5100
rect 9220 5090 9230 5100
rect 9410 5090 9420 5100
rect 9740 5090 9750 5100
rect 590 5080 640 5090
rect 690 5080 750 5090
rect 1790 5080 1810 5090
rect 1820 5080 1880 5090
rect 1980 5080 2100 5090
rect 2860 5080 2870 5090
rect 3410 5080 3420 5090
rect 5170 5080 5180 5090
rect 5200 5080 5210 5090
rect 7310 5080 7450 5090
rect 7880 5080 7990 5090
rect 8020 5080 8040 5090
rect 8110 5080 8120 5090
rect 8130 5080 8140 5090
rect 8150 5080 8170 5090
rect 8190 5080 8220 5090
rect 8390 5080 8420 5090
rect 8460 5080 8470 5090
rect 8760 5080 8780 5090
rect 9130 5080 9140 5090
rect 9370 5080 9380 5090
rect 9520 5080 9530 5090
rect 9770 5080 9790 5090
rect 600 5070 650 5080
rect 700 5070 740 5080
rect 1770 5070 1870 5080
rect 1970 5070 2080 5080
rect 2860 5070 2870 5080
rect 2880 5070 2890 5080
rect 5170 5070 5200 5080
rect 7310 5070 7450 5080
rect 7880 5070 7990 5080
rect 8030 5070 8040 5080
rect 8120 5070 8140 5080
rect 8160 5070 8210 5080
rect 8270 5070 8280 5080
rect 8400 5070 8430 5080
rect 8470 5070 8490 5080
rect 8660 5070 8680 5080
rect 8770 5070 8780 5080
rect 9200 5070 9210 5080
rect 9370 5070 9380 5080
rect 9600 5070 9610 5080
rect 430 5060 480 5070
rect 490 5060 500 5070
rect 610 5060 650 5070
rect 1760 5060 1880 5070
rect 1980 5060 2080 5070
rect 2870 5060 2980 5070
rect 5180 5060 5200 5070
rect 7310 5060 7450 5070
rect 7890 5060 7990 5070
rect 8030 5060 8050 5070
rect 8130 5060 8170 5070
rect 8180 5060 8240 5070
rect 8250 5060 8280 5070
rect 8410 5060 8430 5070
rect 8520 5060 8530 5070
rect 8670 5060 8680 5070
rect 8710 5060 8720 5070
rect 8780 5060 8790 5070
rect 9090 5060 9100 5070
rect 9380 5060 9390 5070
rect 9440 5060 9450 5070
rect 9580 5060 9590 5070
rect 380 5050 650 5060
rect 1770 5050 1880 5060
rect 1990 5050 2090 5060
rect 2890 5050 3040 5060
rect 3300 5050 3310 5060
rect 3320 5050 3330 5060
rect 5180 5050 5200 5060
rect 7320 5050 7450 5060
rect 7900 5050 7990 5060
rect 8030 5050 8050 5060
rect 8110 5050 8120 5060
rect 8130 5050 8180 5060
rect 8250 5050 8280 5060
rect 8340 5050 8370 5060
rect 8410 5050 8430 5060
rect 8670 5050 8680 5060
rect 9090 5050 9100 5060
rect 9270 5050 9280 5060
rect 380 5040 480 5050
rect 500 5040 620 5050
rect 1780 5040 1880 5050
rect 1990 5040 2100 5050
rect 2860 5040 2870 5050
rect 2890 5040 2940 5050
rect 2960 5040 3050 5050
rect 3080 5040 3090 5050
rect 3310 5040 3330 5050
rect 3380 5040 3390 5050
rect 5180 5040 5200 5050
rect 7370 5040 7390 5050
rect 7420 5040 7430 5050
rect 7900 5040 7980 5050
rect 8030 5040 8050 5050
rect 8110 5040 8160 5050
rect 8260 5040 8280 5050
rect 8340 5040 8350 5050
rect 8360 5040 8370 5050
rect 8420 5040 8430 5050
rect 8710 5040 8720 5050
rect 9090 5040 9110 5050
rect 9270 5040 9280 5050
rect 9420 5040 9430 5050
rect 9530 5040 9540 5050
rect 380 5030 470 5040
rect 1760 5030 1780 5040
rect 1790 5030 1890 5040
rect 1990 5030 2110 5040
rect 2830 5030 2870 5040
rect 2890 5030 2940 5040
rect 2960 5030 3050 5040
rect 3330 5030 3340 5040
rect 3370 5030 3400 5040
rect 5180 5030 5200 5040
rect 7310 5030 7350 5040
rect 7400 5030 7440 5040
rect 7900 5030 7980 5040
rect 8030 5030 8090 5040
rect 8100 5030 8150 5040
rect 8270 5030 8280 5040
rect 8350 5030 8360 5040
rect 8400 5030 8440 5040
rect 8700 5030 8710 5040
rect 9020 5030 9030 5040
rect 9130 5030 9140 5040
rect 9470 5030 9480 5040
rect 9490 5030 9500 5040
rect 180 5020 190 5030
rect 380 5020 470 5030
rect 1750 5020 1790 5030
rect 1800 5020 1880 5030
rect 1990 5020 2110 5030
rect 2830 5020 2940 5030
rect 2960 5020 3050 5030
rect 3360 5020 3370 5030
rect 3390 5020 3400 5030
rect 5180 5020 5200 5030
rect 7320 5020 7350 5030
rect 7390 5020 7400 5030
rect 7440 5020 7460 5030
rect 7900 5020 7990 5030
rect 8030 5020 8090 5030
rect 8110 5020 8140 5030
rect 8270 5020 8290 5030
rect 8430 5020 8440 5030
rect 8960 5020 8970 5030
rect 9000 5020 9010 5030
rect 9070 5020 9080 5030
rect 9130 5020 9140 5030
rect 9280 5020 9290 5030
rect 9390 5020 9400 5030
rect 400 5010 460 5020
rect 1750 5010 1800 5020
rect 1810 5010 1870 5020
rect 2000 5010 2120 5020
rect 2820 5010 2940 5020
rect 2950 5010 3040 5020
rect 3350 5010 3360 5020
rect 5180 5010 5200 5020
rect 7310 5010 7350 5020
rect 7430 5010 7450 5020
rect 7460 5010 7480 5020
rect 7880 5010 7990 5020
rect 8040 5010 8080 5020
rect 8120 5010 8140 5020
rect 8190 5010 8230 5020
rect 8270 5010 8290 5020
rect 8390 5010 8400 5020
rect 8430 5010 8440 5020
rect 8480 5010 8490 5020
rect 8880 5010 8890 5020
rect 9030 5010 9040 5020
rect 9130 5010 9140 5020
rect 9180 5010 9190 5020
rect 9280 5010 9290 5020
rect 9390 5010 9400 5020
rect 9500 5010 9510 5020
rect 190 5000 210 5010
rect 410 5000 430 5010
rect 440 5000 460 5010
rect 1760 5000 1820 5010
rect 2020 5000 2120 5010
rect 2760 5000 3030 5010
rect 3340 5000 3360 5010
rect 3370 5000 3390 5010
rect 5180 5000 5200 5010
rect 7320 5000 7340 5010
rect 7370 5000 7380 5010
rect 7470 5000 7500 5010
rect 7890 5000 7910 5010
rect 7930 5000 7990 5010
rect 8050 5000 8080 5010
rect 8120 5000 8130 5010
rect 8190 5000 8220 5010
rect 8270 5000 8290 5010
rect 8430 5000 8440 5010
rect 8860 5000 8880 5010
rect 8930 5000 8940 5010
rect 8950 5000 8960 5010
rect 9030 5000 9040 5010
rect 9140 5000 9150 5010
rect 9480 5000 9490 5010
rect 210 4990 220 5000
rect 410 4990 430 5000
rect 450 4990 460 5000
rect 1770 4990 1820 5000
rect 1830 4990 1840 5000
rect 2020 4990 2030 5000
rect 2040 4990 2050 5000
rect 2060 4990 2120 5000
rect 2760 4990 3000 5000
rect 3330 4990 3350 5000
rect 3370 4990 3390 5000
rect 5750 4990 5760 5000
rect 7320 4990 7350 5000
rect 7500 4990 7530 5000
rect 7890 4990 7990 5000
rect 8050 4990 8070 5000
rect 8130 4990 8150 5000
rect 8190 4990 8230 5000
rect 8280 4990 8300 5000
rect 8390 4990 8400 5000
rect 8440 4990 8450 5000
rect 8540 4990 8550 5000
rect 8870 4990 8880 5000
rect 8930 4990 8960 5000
rect 9010 4990 9040 5000
rect 9400 4990 9410 5000
rect 9440 4990 9450 5000
rect 420 4980 440 4990
rect 450 4980 480 4990
rect 1780 4980 1830 4990
rect 2060 4980 2130 4990
rect 2760 4980 2990 4990
rect 3260 4980 3270 4990
rect 3330 4980 3350 4990
rect 5720 4980 5760 4990
rect 7320 4980 7350 4990
rect 7860 4980 7870 4990
rect 7890 4980 7990 4990
rect 8190 4980 8230 4990
rect 8280 4980 8300 4990
rect 8440 4980 8450 4990
rect 8520 4980 8530 4990
rect 8830 4980 8840 4990
rect 8870 4980 8880 4990
rect 8940 4980 8960 4990
rect 9010 4980 9020 4990
rect 9030 4980 9040 4990
rect 9140 4980 9150 4990
rect 9690 4980 9700 4990
rect 420 4970 440 4980
rect 450 4970 500 4980
rect 1800 4970 1830 4980
rect 2060 4970 2140 4980
rect 2680 4970 2690 4980
rect 2760 4970 2970 4980
rect 3350 4970 3370 4980
rect 4010 4970 4020 4980
rect 4030 4970 4040 4980
rect 4050 4970 4060 4980
rect 4210 4970 4270 4980
rect 4320 4970 4330 4980
rect 4350 4970 4360 4980
rect 4530 4970 4540 4980
rect 4550 4970 4560 4980
rect 4570 4970 4580 4980
rect 5720 4970 5750 4980
rect 7320 4970 7350 4980
rect 7840 4970 7990 4980
rect 8130 4970 8140 4980
rect 8200 4970 8230 4980
rect 8280 4970 8300 4980
rect 8410 4970 8420 4980
rect 8480 4970 8490 4980
rect 8740 4970 8750 4980
rect 8870 4970 8880 4980
rect 8950 4970 8960 4980
rect 9030 4970 9050 4980
rect 9080 4970 9090 4980
rect 9150 4970 9160 4980
rect 9190 4970 9200 4980
rect 9650 4970 9660 4980
rect 9710 4970 9720 4980
rect 420 4960 440 4970
rect 450 4960 550 4970
rect 1820 4960 1830 4970
rect 2100 4960 2150 4970
rect 2640 4960 2690 4970
rect 2700 4960 2710 4970
rect 2760 4960 2950 4970
rect 3340 4960 3350 4970
rect 3360 4960 3380 4970
rect 4200 4960 4210 4970
rect 4340 4960 4350 4970
rect 4370 4960 4380 4970
rect 5700 4960 5740 4970
rect 6350 4960 6370 4970
rect 7330 4960 7350 4970
rect 7840 4960 7850 4970
rect 7920 4960 7990 4970
rect 8210 4960 8230 4970
rect 8280 4960 8300 4970
rect 8340 4960 8350 4970
rect 8360 4960 8370 4970
rect 8670 4960 8710 4970
rect 8870 4960 8880 4970
rect 9040 4960 9050 4970
rect 9150 4960 9160 4970
rect 9310 4960 9330 4970
rect 9620 4960 9630 4970
rect 270 4950 280 4960
rect 420 4950 440 4960
rect 450 4950 560 4960
rect 1850 4950 1890 4960
rect 2120 4950 2160 4960
rect 2640 4950 2910 4960
rect 2920 4950 2940 4960
rect 3230 4950 3250 4960
rect 3340 4950 3350 4960
rect 3360 4950 3370 4960
rect 4040 4950 4050 4960
rect 4070 4950 4080 4960
rect 4190 4950 4200 4960
rect 4330 4950 4350 4960
rect 4360 4950 4380 4960
rect 5690 4950 5730 4960
rect 6350 4950 6380 4960
rect 7330 4950 7340 4960
rect 7940 4950 7990 4960
rect 8130 4950 8150 4960
rect 8200 4950 8230 4960
rect 8280 4950 8310 4960
rect 8640 4950 8650 4960
rect 8710 4950 8720 4960
rect 8730 4950 8740 4960
rect 8780 4950 8820 4960
rect 8880 4950 8890 4960
rect 9150 4950 9160 4960
rect 9200 4950 9210 4960
rect 9700 4950 9710 4960
rect 280 4940 330 4950
rect 400 4940 430 4950
rect 440 4940 590 4950
rect 1040 4940 1050 4950
rect 1860 4940 1890 4950
rect 2130 4940 2170 4950
rect 2270 4940 2320 4950
rect 2650 4940 2900 4950
rect 2920 4940 2930 4950
rect 3220 4940 3230 4950
rect 3330 4940 3360 4950
rect 4080 4940 4090 4950
rect 4190 4940 4200 4950
rect 4410 4940 4420 4950
rect 4670 4940 4700 4950
rect 5670 4940 5730 4950
rect 6350 4940 6400 4950
rect 7330 4940 7340 4950
rect 7940 4940 7990 4950
rect 8140 4940 8160 4950
rect 8200 4940 8220 4950
rect 8280 4940 8310 4950
rect 8340 4940 8350 4950
rect 8730 4940 8740 4950
rect 8800 4940 8820 4950
rect 8880 4940 8890 4950
rect 9020 4940 9030 4950
rect 9050 4940 9060 4950
rect 9140 4940 9160 4950
rect 9250 4940 9260 4950
rect 9540 4940 9550 4950
rect 9570 4940 9580 4950
rect 9670 4940 9680 4950
rect 260 4930 320 4940
rect 360 4930 610 4940
rect 1040 4930 1060 4940
rect 1860 4930 1890 4940
rect 2150 4930 2170 4940
rect 2190 4930 2210 4940
rect 2260 4930 2320 4940
rect 2640 4930 2890 4940
rect 3220 4930 3230 4940
rect 3340 4930 3360 4940
rect 4000 4930 4010 4940
rect 4350 4930 4360 4940
rect 4370 4930 4380 4940
rect 4430 4930 4440 4940
rect 4520 4930 4540 4940
rect 5650 4930 5720 4940
rect 5860 4930 5880 4940
rect 6350 4930 6400 4940
rect 7330 4930 7340 4940
rect 7760 4930 7770 4940
rect 7790 4930 7830 4940
rect 7950 4930 7990 4940
rect 8140 4930 8160 4940
rect 8310 4930 8320 4940
rect 8780 4930 8800 4940
rect 8810 4930 8820 4940
rect 8890 4930 8900 4940
rect 9090 4930 9100 4940
rect 9130 4930 9140 4940
rect 9270 4930 9280 4940
rect 9650 4930 9660 4940
rect 220 4920 320 4930
rect 380 4920 640 4930
rect 1040 4920 1060 4930
rect 2160 4920 2210 4930
rect 2250 4920 2280 4930
rect 2290 4920 2330 4930
rect 2660 4920 2880 4930
rect 3210 4920 3220 4930
rect 3300 4920 3310 4930
rect 3340 4920 3360 4930
rect 4000 4920 4010 4930
rect 4040 4920 4050 4930
rect 4400 4920 4410 4930
rect 4450 4920 4470 4930
rect 4550 4920 4580 4930
rect 5650 4920 5690 4930
rect 5700 4920 5720 4930
rect 5830 4920 5840 4930
rect 5900 4920 5910 4930
rect 6280 4920 6290 4930
rect 6340 4920 6410 4930
rect 7330 4920 7340 4930
rect 7800 4920 7820 4930
rect 7870 4920 7890 4930
rect 7950 4920 8000 4930
rect 8140 4920 8160 4930
rect 8670 4920 8690 4930
rect 8780 4920 8810 4930
rect 8990 4920 9000 4930
rect 9120 4920 9130 4930
rect 9280 4920 9290 4930
rect 9470 4920 9480 4930
rect 9610 4920 9620 4930
rect 90 4910 150 4920
rect 190 4910 330 4920
rect 410 4910 670 4920
rect 680 4910 690 4920
rect 1040 4910 1070 4920
rect 2160 4910 2240 4920
rect 2250 4910 2280 4920
rect 2290 4910 2330 4920
rect 2650 4910 2880 4920
rect 3210 4910 3220 4920
rect 3320 4910 3360 4920
rect 3910 4910 3920 4920
rect 3980 4910 3990 4920
rect 4140 4910 4150 4920
rect 4190 4910 4210 4920
rect 4390 4910 4410 4920
rect 4430 4910 4440 4920
rect 4470 4910 4490 4920
rect 4590 4910 4630 4920
rect 5630 4910 5710 4920
rect 5820 4910 5840 4920
rect 5920 4910 5930 4920
rect 6220 4910 6230 4920
rect 6290 4910 6420 4920
rect 7330 4910 7340 4920
rect 7720 4910 7730 4920
rect 7750 4910 7760 4920
rect 7800 4910 7820 4920
rect 7870 4910 7890 4920
rect 7950 4910 8000 4920
rect 8140 4910 8170 4920
rect 8500 4910 8510 4920
rect 8550 4910 8560 4920
rect 8590 4910 8600 4920
rect 8740 4910 8750 4920
rect 8940 4910 8950 4920
rect 8980 4910 8990 4920
rect 9110 4910 9120 4920
rect 9290 4910 9300 4920
rect 9530 4910 9540 4920
rect 9580 4910 9590 4920
rect 9670 4910 9680 4920
rect 70 4900 380 4910
rect 420 4900 720 4910
rect 1070 4900 1090 4910
rect 2170 4900 2200 4910
rect 2220 4900 2270 4910
rect 2300 4900 2330 4910
rect 2640 4900 2860 4910
rect 3190 4900 3220 4910
rect 3980 4900 3990 4910
rect 4000 4900 4010 4910
rect 4020 4900 4030 4910
rect 4180 4900 4200 4910
rect 4490 4900 4520 4910
rect 4540 4900 4550 4910
rect 4630 4900 4710 4910
rect 5610 4900 5700 4910
rect 5820 4900 5860 4910
rect 5940 4900 5950 4910
rect 6140 4900 6170 4910
rect 6290 4900 6430 4910
rect 7330 4900 7350 4910
rect 7680 4900 7690 4910
rect 7730 4900 7760 4910
rect 7810 4900 7820 4910
rect 7870 4900 7900 4910
rect 7950 4900 8000 4910
rect 8150 4900 8180 4910
rect 8230 4900 8260 4910
rect 8470 4900 8480 4910
rect 8570 4900 8610 4910
rect 8740 4900 8750 4910
rect 8840 4900 8850 4910
rect 8900 4900 8910 4910
rect 8940 4900 8960 4910
rect 9030 4900 9040 4910
rect 9090 4900 9110 4910
rect 50 4890 740 4900
rect 1070 4890 1080 4900
rect 2180 4890 2200 4900
rect 2220 4890 2240 4900
rect 2250 4890 2260 4900
rect 2310 4890 2340 4900
rect 2640 4890 2830 4900
rect 3170 4890 3210 4900
rect 3290 4890 3310 4900
rect 3900 4890 3910 4900
rect 4160 4890 4170 4900
rect 4190 4890 4200 4900
rect 4470 4890 4490 4900
rect 4500 4890 4540 4900
rect 4550 4890 4600 4900
rect 4670 4890 4700 4900
rect 4740 4890 4750 4900
rect 5600 4890 5690 4900
rect 5820 4890 5880 4900
rect 5950 4890 5960 4900
rect 6130 4890 6180 4900
rect 6300 4890 6440 4900
rect 7330 4890 7360 4900
rect 7670 4890 7690 4900
rect 7740 4890 7770 4900
rect 7810 4890 7830 4900
rect 7870 4890 7900 4900
rect 7950 4890 8000 4900
rect 8090 4890 8100 4900
rect 8200 4890 8210 4900
rect 8590 4890 8610 4900
rect 8650 4890 8660 4900
rect 8700 4890 8710 4900
rect 9500 4890 9510 4900
rect 9710 4890 9720 4900
rect 40 4880 490 4890
rect 500 4880 740 4890
rect 1040 4880 1050 4890
rect 1060 4880 1080 4890
rect 2190 4880 2240 4890
rect 2250 4880 2260 4890
rect 2280 4880 2360 4890
rect 2660 4880 2810 4890
rect 3160 4880 3200 4890
rect 3310 4880 3320 4890
rect 3730 4880 3740 4890
rect 3900 4880 3910 4890
rect 3940 4880 3950 4890
rect 3970 4880 3980 4890
rect 4000 4880 4010 4890
rect 4170 4880 4180 4890
rect 4190 4880 4200 4890
rect 4510 4880 4550 4890
rect 4580 4880 4620 4890
rect 4640 4880 4650 4890
rect 4670 4880 4680 4890
rect 4740 4880 4790 4890
rect 5590 4880 5680 4890
rect 5830 4880 5890 4890
rect 5960 4880 5970 4890
rect 6050 4880 6090 4890
rect 6120 4880 6160 4890
rect 6300 4880 6440 4890
rect 7350 4880 7370 4890
rect 7670 4880 7690 4890
rect 7750 4880 7770 4890
rect 7810 4880 7830 4890
rect 7870 4880 7900 4890
rect 7950 4880 8000 4890
rect 8070 4880 8080 4890
rect 8100 4880 8110 4890
rect 8460 4880 8470 4890
rect 8590 4880 8610 4890
rect 8750 4880 8760 4890
rect 9090 4880 9100 4890
rect 9450 4880 9460 4890
rect 9620 4880 9630 4890
rect 9690 4880 9700 4890
rect 30 4870 760 4880
rect 1060 4870 1090 4880
rect 2200 4870 2210 4880
rect 2220 4870 2240 4880
rect 2250 4870 2260 4880
rect 2270 4870 2300 4880
rect 2340 4870 2350 4880
rect 2660 4870 2800 4880
rect 3150 4870 3190 4880
rect 3710 4870 3740 4880
rect 3870 4870 3890 4880
rect 3940 4870 3970 4880
rect 4180 4870 4200 4880
rect 4570 4870 4610 4880
rect 4780 4870 4830 4880
rect 5590 4870 5680 4880
rect 5850 4870 5980 4880
rect 6030 4870 6140 4880
rect 6300 4870 6410 4880
rect 6440 4870 6450 4880
rect 7340 4870 7350 4880
rect 7670 4870 7690 4880
rect 7810 4870 7830 4880
rect 7880 4870 7910 4880
rect 7960 4870 8000 4880
rect 8070 4870 8090 4880
rect 8100 4870 8110 4880
rect 8460 4870 8470 4880
rect 8510 4870 8550 4880
rect 8600 4870 8610 4880
rect 8700 4870 8710 4880
rect 8750 4870 8760 4880
rect 8790 4870 8800 4880
rect 8860 4870 8870 4880
rect 8910 4870 8920 4880
rect 9080 4870 9090 4880
rect 9380 4870 9390 4880
rect 9420 4870 9430 4880
rect 9450 4870 9460 4880
rect 9590 4870 9600 4880
rect 9620 4870 9630 4880
rect 30 4860 40 4870
rect 70 4860 760 4870
rect 1010 4860 1020 4870
rect 1060 4860 1100 4870
rect 2240 4860 2250 4870
rect 2260 4860 2280 4870
rect 2330 4860 2350 4870
rect 2660 4860 2790 4870
rect 3100 4860 3120 4870
rect 3140 4860 3190 4870
rect 3690 4860 3710 4870
rect 3720 4860 3730 4870
rect 3920 4860 3930 4870
rect 3970 4860 3980 4870
rect 4190 4860 4200 4870
rect 4850 4860 4870 4870
rect 4920 4860 4940 4870
rect 5580 4860 5680 4870
rect 5850 4860 5910 4870
rect 5920 4860 5980 4870
rect 6010 4860 6120 4870
rect 6220 4860 6230 4870
rect 6300 4860 6370 4870
rect 6380 4860 6420 4870
rect 6440 4860 6460 4870
rect 7360 4860 7390 4870
rect 7470 4860 7480 4870
rect 7680 4860 7690 4870
rect 7820 4860 7830 4870
rect 7880 4860 7900 4870
rect 7960 4860 8010 4870
rect 8070 4860 8090 4870
rect 8320 4860 8340 4870
rect 8350 4860 8360 4870
rect 8460 4860 8470 4870
rect 8510 4860 8540 4870
rect 8600 4860 8620 4870
rect 8680 4860 8690 4870
rect 8870 4860 8880 4870
rect 8920 4860 8930 4870
rect 80 4850 350 4860
rect 370 4850 750 4860
rect 1070 4850 1120 4860
rect 2330 4850 2350 4860
rect 2670 4850 2780 4860
rect 3100 4850 3180 4860
rect 3320 4850 3330 4860
rect 3680 4850 3690 4860
rect 3840 4850 3850 4860
rect 3860 4850 3870 4860
rect 3960 4850 3970 4860
rect 4890 4850 4900 4860
rect 4940 4850 4950 4860
rect 5570 4850 5670 4860
rect 5960 4850 6120 4860
rect 6160 4850 6230 4860
rect 6280 4850 6360 4860
rect 6370 4850 6420 4860
rect 6430 4850 6460 4860
rect 7360 4850 7380 4860
rect 7390 4850 7410 4860
rect 7680 4850 7700 4860
rect 7820 4850 7830 4860
rect 7880 4850 7890 4860
rect 7950 4850 8020 4860
rect 8060 4850 8080 4860
rect 8250 4850 8280 4860
rect 8510 4850 8540 4860
rect 8580 4850 8590 4860
rect 8650 4850 8660 4860
rect 8830 4850 8840 4860
rect 9060 4850 9080 4860
rect 9330 4850 9340 4860
rect 9720 4850 9740 4860
rect 80 4840 90 4850
rect 100 4840 790 4850
rect 1030 4840 1100 4850
rect 1110 4840 1120 4850
rect 2330 4840 2350 4850
rect 2680 4840 2780 4850
rect 3090 4840 3130 4850
rect 3150 4840 3160 4850
rect 3240 4840 3250 4850
rect 3260 4840 3270 4850
rect 3320 4840 3330 4850
rect 3340 4840 3360 4850
rect 3670 4840 3680 4850
rect 3860 4840 3870 4850
rect 3950 4840 3960 4850
rect 3980 4840 3990 4850
rect 4260 4840 4270 4850
rect 4950 4840 4960 4850
rect 5560 4840 5670 4850
rect 5990 4840 6120 4850
rect 6140 4840 6220 4850
rect 6270 4840 6470 4850
rect 7340 4840 7350 4850
rect 7680 4840 7700 4850
rect 7820 4840 7830 4850
rect 7950 4840 8050 4850
rect 8060 4840 8090 4850
rect 8250 4840 8280 4850
rect 8370 4840 8380 4850
rect 8470 4840 8480 4850
rect 8760 4840 8770 4850
rect 8850 4840 8870 4850
rect 9060 4840 9070 4850
rect 9390 4840 9400 4850
rect 9460 4840 9470 4850
rect 9560 4840 9570 4850
rect 9600 4840 9610 4850
rect 9630 4840 9640 4850
rect 9680 4840 9690 4850
rect 170 4830 350 4840
rect 390 4830 790 4840
rect 1030 4830 1070 4840
rect 1100 4830 1110 4840
rect 2340 4830 2350 4840
rect 2690 4830 2790 4840
rect 3080 4830 3130 4840
rect 3140 4830 3150 4840
rect 3160 4830 3170 4840
rect 3230 4830 3240 4840
rect 3260 4830 3270 4840
rect 3320 4830 3360 4840
rect 3670 4830 3680 4840
rect 3700 4830 3710 4840
rect 3720 4830 3750 4840
rect 3810 4830 3820 4840
rect 3850 4830 3860 4840
rect 4910 4830 4960 4840
rect 4970 4830 4980 4840
rect 5550 4830 5600 4840
rect 5620 4830 5660 4840
rect 5980 4830 6230 4840
rect 6250 4830 6370 4840
rect 6380 4830 6480 4840
rect 7340 4830 7350 4840
rect 7680 4830 7700 4840
rect 7740 4830 7750 4840
rect 7820 4830 7830 4840
rect 7940 4830 8090 4840
rect 8220 4830 8230 4840
rect 8240 4830 8270 4840
rect 8470 4830 8480 4840
rect 8680 4830 8700 4840
rect 9390 4830 9400 4840
rect 9430 4830 9440 4840
rect 9560 4830 9570 4840
rect 9750 4830 9760 4840
rect 0 4820 40 4830
rect 200 4820 330 4830
rect 470 4820 490 4830
rect 510 4820 730 4830
rect 1020 4820 1090 4830
rect 1140 4820 1150 4830
rect 2350 4820 2360 4830
rect 2710 4820 2790 4830
rect 3070 4820 3120 4830
rect 3140 4820 3150 4830
rect 3230 4820 3250 4830
rect 3330 4820 3350 4830
rect 3650 4820 3660 4830
rect 3700 4820 3750 4830
rect 3770 4820 3780 4830
rect 3800 4820 3810 4830
rect 3960 4820 3970 4830
rect 4910 4820 4920 4830
rect 4930 4820 4940 4830
rect 4950 4820 4970 4830
rect 5550 4820 5600 4830
rect 5620 4820 5670 4830
rect 5980 4820 6370 4830
rect 6380 4820 6480 4830
rect 7360 4820 7370 4830
rect 7570 4820 7590 4830
rect 7690 4820 7710 4830
rect 7750 4820 7760 4830
rect 7830 4820 7850 4830
rect 7930 4820 8080 4830
rect 8190 4820 8200 4830
rect 8230 4820 8270 4830
rect 8620 4820 8630 4830
rect 9520 4820 9530 4830
rect 220 4810 280 4820
rect 290 4810 310 4820
rect 540 4810 680 4820
rect 840 4810 870 4820
rect 980 4810 990 4820
rect 1030 4810 1100 4820
rect 2350 4810 2360 4820
rect 2710 4810 2810 4820
rect 3050 4810 3140 4820
rect 3210 4810 3220 4820
rect 3320 4810 3360 4820
rect 3640 4810 3650 4820
rect 3690 4810 3710 4820
rect 3720 4810 3740 4820
rect 3760 4810 3770 4820
rect 3780 4810 3790 4820
rect 3800 4810 3810 4820
rect 3910 4810 3920 4820
rect 4910 4810 4930 4820
rect 4970 4810 4980 4820
rect 5210 4810 5240 4820
rect 5520 4810 5590 4820
rect 5620 4810 5660 4820
rect 5980 4810 6490 4820
rect 7350 4810 7370 4820
rect 7450 4810 7460 4820
rect 7690 4810 7710 4820
rect 7750 4810 7770 4820
rect 7830 4810 7860 4820
rect 7900 4810 7910 4820
rect 7930 4810 7940 4820
rect 7950 4810 7970 4820
rect 7980 4810 8090 4820
rect 8120 4810 8130 4820
rect 8190 4810 8200 4820
rect 8240 4810 8270 4820
rect 8310 4810 8320 4820
rect 8530 4810 8540 4820
rect 8620 4810 8630 4820
rect 9040 4810 9050 4820
rect 9330 4810 9340 4820
rect 9470 4810 9480 4820
rect 9510 4810 9520 4820
rect 130 4800 150 4810
rect 230 4800 290 4810
rect 330 4800 460 4810
rect 550 4800 580 4810
rect 600 4800 630 4810
rect 740 4800 880 4810
rect 1030 4800 1040 4810
rect 1050 4800 1100 4810
rect 1140 4800 1150 4810
rect 2350 4800 2370 4810
rect 2750 4800 2840 4810
rect 3040 4800 3130 4810
rect 3140 4800 3150 4810
rect 3220 4800 3250 4810
rect 3310 4800 3370 4810
rect 3630 4800 3640 4810
rect 3680 4800 3690 4810
rect 3780 4800 3790 4810
rect 3900 4800 3910 4810
rect 4910 4800 4960 4810
rect 4970 4800 5000 4810
rect 5010 4800 5020 4810
rect 5210 4800 5240 4810
rect 5510 4800 5560 4810
rect 5620 4800 5660 4810
rect 5980 4800 6250 4810
rect 6290 4800 6320 4810
rect 6360 4800 6510 4810
rect 7350 4800 7370 4810
rect 7520 4800 7540 4810
rect 7690 4800 7710 4810
rect 7750 4800 7780 4810
rect 7930 4800 7940 4810
rect 7980 4800 8120 4810
rect 8160 4800 8200 4810
rect 8240 4800 8270 4810
rect 8310 4800 8360 4810
rect 8480 4800 8490 4810
rect 8520 4800 8530 4810
rect 8710 4800 8720 4810
rect 9020 4800 9030 4810
rect 9400 4800 9410 4810
rect 9570 4800 9580 4810
rect 110 4790 140 4800
rect 150 4790 160 4800
rect 170 4790 180 4800
rect 210 4790 250 4800
rect 300 4790 480 4800
rect 550 4790 580 4800
rect 600 4790 880 4800
rect 890 4790 900 4800
rect 1030 4790 1100 4800
rect 2360 4790 2390 4800
rect 2760 4790 2920 4800
rect 3040 4790 3130 4800
rect 3240 4790 3260 4800
rect 3270 4790 3280 4800
rect 3320 4790 3360 4800
rect 3620 4790 3630 4800
rect 3880 4790 3890 4800
rect 4930 4790 4940 4800
rect 4990 4790 5000 4800
rect 5190 4790 5230 4800
rect 5500 4790 5560 4800
rect 5610 4790 5650 4800
rect 5990 4790 6230 4800
rect 6360 4790 6510 4800
rect 7350 4790 7370 4800
rect 7510 4790 7520 4800
rect 7690 4790 7710 4800
rect 7750 4790 7780 4800
rect 7790 4790 7800 4800
rect 7810 4790 7820 4800
rect 7920 4790 7940 4800
rect 7980 4790 8030 4800
rect 8070 4790 8120 4800
rect 8170 4790 8200 4800
rect 8250 4790 8270 4800
rect 8630 4790 8640 4800
rect 8670 4790 8680 4800
rect 8990 4790 9000 4800
rect 110 4780 130 4790
rect 180 4780 320 4790
rect 460 4780 520 4790
rect 600 4780 880 4790
rect 900 4780 920 4790
rect 1040 4780 1100 4790
rect 2360 4780 2370 4790
rect 2430 4780 2440 4790
rect 2800 4780 2930 4790
rect 3030 4780 3120 4790
rect 3320 4780 3340 4790
rect 3870 4780 3880 4790
rect 3890 4780 3900 4790
rect 5210 4780 5220 4790
rect 5490 4780 5550 4790
rect 5610 4780 5640 4790
rect 5990 4780 6210 4790
rect 6380 4780 6520 4790
rect 7350 4780 7370 4790
rect 7500 4780 7510 4790
rect 7700 4780 7710 4790
rect 7990 4780 8010 4790
rect 8090 4780 8120 4790
rect 8180 4780 8200 4790
rect 8250 4780 8280 4790
rect 9480 4780 9490 4790
rect 140 4770 310 4780
rect 480 4770 550 4780
rect 590 4770 850 4780
rect 880 4770 900 4780
rect 1050 4770 1060 4780
rect 1070 4770 1110 4780
rect 2390 4770 2420 4780
rect 2430 4770 2440 4780
rect 2820 4770 2930 4780
rect 3020 4770 3110 4780
rect 3120 4770 3130 4780
rect 3280 4770 3290 4780
rect 3330 4770 3340 4780
rect 3620 4770 3630 4780
rect 3800 4770 3810 4780
rect 3880 4770 3890 4780
rect 5040 4770 5050 4780
rect 5480 4770 5530 4780
rect 5600 4770 5630 4780
rect 6010 4770 6130 4780
rect 6140 4770 6190 4780
rect 6390 4770 6530 4780
rect 7350 4770 7360 4780
rect 7480 4770 7500 4780
rect 7710 4770 7720 4780
rect 7960 4770 8000 4780
rect 8110 4770 8120 4780
rect 8250 4770 8290 4780
rect 8490 4770 8500 4780
rect 8530 4770 8540 4780
rect 9410 4770 9420 4780
rect 160 4760 320 4770
rect 500 4760 960 4770
rect 990 4760 1010 4770
rect 1080 4760 1130 4770
rect 2380 4760 2420 4770
rect 2430 4760 2450 4770
rect 2830 4760 2940 4770
rect 3000 4760 3100 4770
rect 3290 4760 3300 4770
rect 3330 4760 3340 4770
rect 3590 4760 3600 4770
rect 3610 4760 3620 4770
rect 3790 4760 3810 4770
rect 5060 4760 5070 4770
rect 5470 4760 5530 4770
rect 5580 4760 5620 4770
rect 6030 4760 6110 4770
rect 6400 4760 6540 4770
rect 7470 4760 7480 4770
rect 7930 4760 7950 4770
rect 7960 4760 7990 4770
rect 8250 4760 8260 4770
rect 8300 4760 8360 4770
rect 8820 4760 8830 4770
rect 8850 4760 8860 4770
rect 9000 4760 9010 4770
rect 9300 4760 9310 4770
rect 9410 4760 9420 4770
rect 150 4750 350 4760
rect 530 4750 950 4760
rect 990 4750 1010 4760
rect 1070 4750 1140 4760
rect 2380 4750 2410 4760
rect 2420 4750 2450 4760
rect 2830 4750 3100 4760
rect 3580 4750 3590 4760
rect 3780 4750 3800 4760
rect 3830 4750 3840 4760
rect 3870 4750 3880 4760
rect 5070 4750 5080 4760
rect 5470 4750 5510 4760
rect 5580 4750 5610 4760
rect 6410 4750 6550 4760
rect 7360 4750 7380 4760
rect 7390 4750 7400 4760
rect 7450 4750 7470 4760
rect 7890 4750 7900 4760
rect 7940 4750 7990 4760
rect 8250 4750 8260 4760
rect 8300 4750 8310 4760
rect 8350 4750 8360 4760
rect 8510 4750 8520 4760
rect 8800 4750 8810 4760
rect 8910 4750 8920 4760
rect 9000 4750 9010 4760
rect 9300 4750 9310 4760
rect 9420 4750 9430 4760
rect 9920 4750 9960 4760
rect 150 4740 370 4750
rect 550 4740 960 4750
rect 980 4740 1000 4750
rect 1010 4740 1020 4750
rect 1090 4740 1110 4750
rect 1140 4740 1170 4750
rect 2400 4740 2410 4750
rect 2420 4740 2450 4750
rect 2470 4740 2480 4750
rect 2850 4740 3090 4750
rect 3290 4740 3300 4750
rect 3340 4740 3350 4750
rect 3520 4740 3530 4750
rect 3780 4740 3800 4750
rect 3820 4740 3830 4750
rect 3840 4740 3850 4750
rect 3910 4740 3930 4750
rect 3980 4740 3990 4750
rect 5080 4740 5090 4750
rect 5470 4740 5510 4750
rect 5570 4740 5600 4750
rect 6420 4740 6560 4750
rect 7440 4740 7460 4750
rect 7870 4740 7880 4750
rect 7960 4740 7980 4750
rect 8260 4740 8290 4750
rect 8320 4740 8330 4750
rect 8340 4740 8350 4750
rect 8390 4740 8400 4750
rect 8910 4740 8920 4750
rect 8980 4740 8990 4750
rect 9000 4740 9010 4750
rect 9310 4740 9320 4750
rect 9870 4740 9880 4750
rect 160 4730 410 4740
rect 570 4730 650 4740
rect 670 4730 1000 4740
rect 1010 4730 1030 4740
rect 1090 4730 1120 4740
rect 1140 4730 1150 4740
rect 2410 4730 2420 4740
rect 2430 4730 2450 4740
rect 2480 4730 2500 4740
rect 2850 4730 3100 4740
rect 3290 4730 3300 4740
rect 3340 4730 3350 4740
rect 3510 4730 3530 4740
rect 3790 4730 3800 4740
rect 3820 4730 3830 4740
rect 5080 4730 5090 4740
rect 5470 4730 5510 4740
rect 5550 4730 5600 4740
rect 6430 4730 6570 4740
rect 7440 4730 7450 4740
rect 7860 4730 7870 4740
rect 7960 4730 7980 4740
rect 8110 4730 8130 4740
rect 8260 4730 8290 4740
rect 8780 4730 8790 4740
rect 9000 4730 9010 4740
rect 9290 4730 9300 4740
rect 9850 4730 9860 4740
rect 150 4720 430 4730
rect 620 4720 640 4730
rect 690 4720 1020 4730
rect 1030 4720 1040 4730
rect 1060 4720 1070 4730
rect 1090 4720 1160 4730
rect 2430 4720 2450 4730
rect 2480 4720 2500 4730
rect 2860 4720 2990 4730
rect 3010 4720 3060 4730
rect 3080 4720 3090 4730
rect 3290 4720 3300 4730
rect 3510 4720 3530 4730
rect 3580 4720 3600 4730
rect 3780 4720 3800 4730
rect 5090 4720 5110 4730
rect 5470 4720 5500 4730
rect 5550 4720 5600 4730
rect 6440 4720 6570 4730
rect 7430 4720 7440 4730
rect 7770 4720 7800 4730
rect 7850 4720 7860 4730
rect 7950 4720 7980 4730
rect 8110 4720 8130 4730
rect 8180 4720 8190 4730
rect 8260 4720 8290 4730
rect 8820 4720 8830 4730
rect 8850 4720 8860 4730
rect 8890 4720 8900 4730
rect 9340 4720 9350 4730
rect 9840 4720 9850 4730
rect 150 4710 450 4720
rect 630 4710 650 4720
rect 710 4710 1040 4720
rect 1100 4710 1170 4720
rect 2430 4710 2460 4720
rect 2470 4710 2530 4720
rect 2850 4710 2980 4720
rect 3010 4710 3060 4720
rect 3080 4710 3090 4720
rect 3290 4710 3310 4720
rect 3500 4710 3530 4720
rect 3550 4710 3560 4720
rect 3580 4710 3600 4720
rect 3770 4710 3800 4720
rect 5110 4710 5130 4720
rect 5460 4710 5500 4720
rect 5550 4710 5600 4720
rect 6440 4710 6580 4720
rect 7410 4710 7440 4720
rect 7730 4710 7740 4720
rect 7810 4710 7820 4720
rect 7830 4710 7850 4720
rect 7900 4710 7980 4720
rect 8110 4710 8130 4720
rect 8180 4710 8200 4720
rect 8270 4710 8290 4720
rect 8850 4710 8860 4720
rect 8920 4710 8930 4720
rect 160 4700 470 4710
rect 660 4700 670 4710
rect 730 4700 990 4710
rect 1000 4700 1030 4710
rect 1080 4700 1090 4710
rect 1100 4700 1170 4710
rect 2440 4700 2450 4710
rect 2470 4700 2540 4710
rect 2840 4700 2850 4710
rect 2890 4700 2960 4710
rect 3020 4700 3060 4710
rect 3090 4700 3100 4710
rect 3170 4700 3180 4710
rect 3290 4700 3320 4710
rect 3500 4700 3520 4710
rect 3540 4700 3550 4710
rect 3770 4700 3790 4710
rect 5120 4700 5130 4710
rect 5460 4700 5500 4710
rect 5570 4700 5610 4710
rect 6460 4700 6580 4710
rect 7400 4700 7430 4710
rect 7720 4700 7730 4710
rect 7830 4700 7850 4710
rect 7900 4700 7990 4710
rect 8040 4700 8060 4710
rect 8120 4700 8140 4710
rect 8180 4700 8210 4710
rect 8300 4700 8310 4710
rect 8340 4700 8350 4710
rect 8600 4700 8610 4710
rect 8670 4700 8680 4710
rect 8970 4700 8980 4710
rect 150 4690 500 4700
rect 670 4690 680 4700
rect 740 4690 1030 4700
rect 1060 4690 1090 4700
rect 1110 4690 1170 4700
rect 2440 4690 2450 4700
rect 2480 4690 2540 4700
rect 2630 4690 2670 4700
rect 2720 4690 2730 4700
rect 2750 4690 2780 4700
rect 2830 4690 2860 4700
rect 2880 4690 2960 4700
rect 3000 4690 3080 4700
rect 3090 4690 3110 4700
rect 3170 4690 3190 4700
rect 3290 4690 3310 4700
rect 3510 4690 3550 4700
rect 3620 4690 3640 4700
rect 5150 4690 5160 4700
rect 5470 4690 5500 4700
rect 5580 4690 5630 4700
rect 6460 4690 6570 4700
rect 7380 4690 7390 4700
rect 7400 4690 7420 4700
rect 7660 4690 7690 4700
rect 7700 4690 7720 4700
rect 7830 4690 7850 4700
rect 7950 4690 8000 4700
rect 8030 4690 8060 4700
rect 8120 4690 8140 4700
rect 8180 4690 8220 4700
rect 8260 4690 8270 4700
rect 8970 4690 8990 4700
rect 140 4680 510 4690
rect 750 4680 1040 4690
rect 1120 4680 1170 4690
rect 2480 4680 2530 4690
rect 2540 4680 2550 4690
rect 2600 4680 2800 4690
rect 2820 4680 2960 4690
rect 3000 4680 3060 4690
rect 3100 4680 3110 4690
rect 3130 4680 3150 4690
rect 3180 4680 3190 4690
rect 3490 4680 3540 4690
rect 3600 4680 3610 4690
rect 3630 4680 3640 4690
rect 5160 4680 5170 4690
rect 5470 4680 5510 4690
rect 5580 4680 5630 4690
rect 6460 4680 6530 4690
rect 6550 4680 6570 4690
rect 7390 4680 7410 4690
rect 7700 4680 7720 4690
rect 7970 4680 7990 4690
rect 8040 4680 8060 4690
rect 8120 4680 8150 4690
rect 8190 4680 8210 4690
rect 8240 4680 8260 4690
rect 8560 4680 8570 4690
rect 8650 4680 8660 4690
rect 8780 4680 8790 4690
rect 8820 4680 8830 4690
rect 8860 4680 8870 4690
rect 8970 4680 9000 4690
rect 130 4670 520 4680
rect 760 4670 1010 4680
rect 1030 4670 1050 4680
rect 1160 4670 1180 4680
rect 2510 4670 2520 4680
rect 2540 4670 2620 4680
rect 2630 4670 2670 4680
rect 2680 4670 2970 4680
rect 2990 4670 3060 4680
rect 3110 4670 3140 4680
rect 3170 4670 3190 4680
rect 3260 4670 3270 4680
rect 3340 4670 3350 4680
rect 3600 4670 3610 4680
rect 3700 4670 3720 4680
rect 5170 4670 5180 4680
rect 5480 4670 5520 4680
rect 5590 4670 5650 4680
rect 6430 4670 6540 4680
rect 6550 4670 6570 4680
rect 7390 4670 7400 4680
rect 7700 4670 7720 4680
rect 7770 4670 7780 4680
rect 7840 4670 7860 4680
rect 7980 4670 8000 4680
rect 8040 4670 8050 4680
rect 8120 4670 8130 4680
rect 8140 4670 8150 4680
rect 8180 4670 8190 4680
rect 8530 4670 8540 4680
rect 8560 4670 8570 4680
rect 8930 4670 8940 4680
rect 8970 4670 8990 4680
rect 9800 4670 9810 4680
rect 90 4660 100 4670
rect 110 4660 540 4670
rect 800 4660 1040 4670
rect 1170 4660 1180 4670
rect 2500 4660 2510 4670
rect 2550 4660 2620 4670
rect 2640 4660 2730 4670
rect 2760 4660 3030 4670
rect 3050 4660 3060 4670
rect 3110 4660 3130 4670
rect 3170 4660 3180 4670
rect 3250 4660 3260 4670
rect 3340 4660 3350 4670
rect 3480 4660 3490 4670
rect 3610 4660 3620 4670
rect 3780 4660 3790 4670
rect 5150 4660 5160 4670
rect 5180 4660 5190 4670
rect 5490 4660 5520 4670
rect 5590 4660 5740 4670
rect 6420 4660 6520 4670
rect 6560 4660 6580 4670
rect 7690 4660 7720 4670
rect 7770 4660 7790 4670
rect 7840 4660 7880 4670
rect 7980 4660 8000 4670
rect 8150 4660 8180 4670
rect 8590 4660 8610 4670
rect 8640 4660 8650 4670
rect 8930 4660 8940 4670
rect 9790 4660 9800 4670
rect 90 4650 560 4660
rect 830 4650 1070 4660
rect 1140 4650 1180 4660
rect 2480 4650 2490 4660
rect 2540 4650 2720 4660
rect 2780 4650 3010 4660
rect 3050 4650 3060 4660
rect 3090 4650 3100 4660
rect 3110 4650 3120 4660
rect 3170 4650 3180 4660
rect 3480 4650 3500 4660
rect 5500 4650 5520 4660
rect 5730 4650 5770 4660
rect 6420 4650 6520 4660
rect 6560 4650 6580 4660
rect 7510 4650 7520 4660
rect 7700 4650 7730 4660
rect 7910 4650 7940 4660
rect 7980 4650 8010 4660
rect 8110 4650 8120 4660
rect 8870 4650 8880 4660
rect 8980 4650 8990 4660
rect 9780 4650 9790 4660
rect 0 4640 30 4650
rect 40 4640 580 4650
rect 840 4640 1090 4650
rect 1100 4640 1110 4650
rect 2490 4640 2500 4650
rect 2540 4640 2550 4650
rect 2560 4640 2720 4650
rect 2770 4640 3010 4650
rect 3030 4640 3070 4650
rect 3110 4640 3130 4650
rect 3150 4640 3180 4650
rect 3470 4640 3490 4650
rect 5140 4640 5150 4650
rect 5190 4640 5200 4650
rect 5500 4640 5530 4650
rect 5760 4640 5830 4650
rect 6080 4640 6190 4650
rect 6200 4640 6230 4650
rect 6410 4640 6510 4650
rect 6560 4640 6580 4650
rect 7380 4640 7390 4650
rect 7570 4640 7580 4650
rect 7590 4640 7600 4650
rect 7640 4640 7650 4650
rect 7710 4640 7730 4650
rect 7920 4640 7940 4650
rect 7980 4640 8010 4650
rect 8100 4640 8110 4650
rect 8790 4640 8800 4650
rect 8830 4640 8840 4650
rect 9770 4640 9780 4650
rect 0 4630 600 4640
rect 840 4630 1120 4640
rect 1180 4630 1190 4640
rect 2490 4630 2500 4640
rect 2590 4630 2720 4640
rect 2780 4630 2800 4640
rect 2810 4630 2820 4640
rect 2830 4630 3000 4640
rect 3020 4630 3030 4640
rect 3040 4630 3050 4640
rect 3080 4630 3090 4640
rect 3100 4630 3110 4640
rect 3130 4630 3160 4640
rect 3170 4630 3180 4640
rect 3460 4630 3480 4640
rect 5150 4630 5160 4640
rect 5170 4630 5180 4640
rect 5510 4630 5540 4640
rect 5750 4630 5760 4640
rect 5790 4630 5860 4640
rect 5870 4630 5960 4640
rect 6050 4630 6240 4640
rect 6410 4630 6500 4640
rect 6560 4630 6580 4640
rect 7380 4630 7390 4640
rect 7580 4630 7590 4640
rect 7640 4630 7700 4640
rect 7720 4630 7730 4640
rect 7870 4630 7880 4640
rect 7910 4630 7930 4640
rect 7980 4630 7990 4640
rect 8010 4630 8020 4640
rect 8080 4630 8120 4640
rect 8300 4630 8310 4640
rect 8360 4630 8370 4640
rect 8490 4630 8500 4640
rect 8850 4630 8860 4640
rect 9760 4630 9770 4640
rect 0 4620 620 4630
rect 850 4620 1120 4630
rect 1130 4620 1200 4630
rect 2600 4620 2710 4630
rect 2720 4620 2800 4630
rect 2880 4620 2890 4630
rect 2910 4620 2970 4630
rect 2980 4620 3000 4630
rect 3010 4620 3030 4630
rect 3120 4620 3130 4630
rect 3140 4620 3160 4630
rect 3460 4620 3480 4630
rect 5160 4620 5170 4630
rect 5200 4620 5210 4630
rect 5520 4620 5540 4630
rect 5610 4620 5630 4630
rect 5750 4620 5770 4630
rect 5800 4620 5970 4630
rect 5980 4620 5990 4630
rect 6020 4620 6490 4630
rect 6560 4620 6570 4630
rect 7380 4620 7400 4630
rect 7470 4620 7480 4630
rect 7590 4620 7600 4630
rect 7720 4620 7730 4630
rect 7970 4620 7990 4630
rect 8080 4620 8120 4630
rect 8370 4620 8380 4630
rect 8490 4620 8500 4630
rect 8560 4620 8570 4630
rect 8650 4620 8660 4630
rect 8800 4620 8810 4630
rect 8900 4620 8910 4630
rect 0 4610 630 4620
rect 860 4610 1220 4620
rect 2730 4610 2750 4620
rect 2840 4610 2890 4620
rect 2920 4610 2960 4620
rect 2970 4610 3000 4620
rect 3010 4610 3020 4620
rect 3130 4610 3170 4620
rect 3230 4610 3240 4620
rect 3290 4610 3300 4620
rect 3460 4610 3480 4620
rect 5520 4610 5540 4620
rect 5600 4610 5640 4620
rect 5750 4610 5770 4620
rect 5780 4610 5800 4620
rect 5810 4610 5890 4620
rect 5900 4610 6110 4620
rect 6160 4610 6360 4620
rect 6380 4610 6480 4620
rect 6530 4610 6570 4620
rect 7390 4610 7400 4620
rect 7470 4610 7480 4620
rect 7520 4610 7550 4620
rect 7590 4610 7610 4620
rect 7730 4610 7740 4620
rect 7830 4610 7840 4620
rect 7860 4610 7870 4620
rect 7960 4610 7980 4620
rect 8070 4610 8120 4620
rect 8230 4610 8240 4620
rect 8270 4610 8280 4620
rect 8380 4610 8390 4620
rect 8490 4610 8500 4620
rect 8650 4610 8660 4620
rect 8890 4610 8900 4620
rect 0 4600 650 4610
rect 870 4600 1220 4610
rect 2850 4600 2930 4610
rect 2990 4600 3000 4610
rect 3010 4600 3020 4610
rect 3030 4600 3040 4610
rect 3050 4600 3060 4610
rect 3130 4600 3160 4610
rect 3220 4600 3240 4610
rect 3360 4600 3370 4610
rect 3450 4600 3470 4610
rect 5180 4600 5190 4610
rect 5530 4600 5540 4610
rect 5570 4600 5610 4610
rect 5640 4600 5650 4610
rect 5750 4600 5790 4610
rect 6000 4600 6080 4610
rect 6180 4600 6190 4610
rect 6510 4600 6560 4610
rect 7390 4600 7410 4610
rect 7470 4600 7480 4610
rect 7540 4600 7550 4610
rect 7590 4600 7600 4610
rect 7730 4600 7740 4610
rect 7840 4600 7850 4610
rect 7870 4600 7880 4610
rect 7950 4600 7960 4610
rect 7970 4600 7980 4610
rect 8070 4600 8130 4610
rect 8190 4600 8210 4610
rect 8260 4600 8280 4610
rect 8490 4600 8500 4610
rect 8870 4600 8880 4610
rect 9240 4600 9250 4610
rect 9730 4600 9740 4610
rect 0 4590 660 4600
rect 870 4590 1210 4600
rect 2820 4590 2830 4600
rect 2850 4590 2870 4600
rect 3030 4590 3050 4600
rect 3130 4590 3170 4600
rect 3200 4590 3220 4600
rect 3230 4590 3240 4600
rect 3270 4590 3280 4600
rect 3360 4590 3370 4600
rect 3450 4590 3460 4600
rect 5180 4590 5190 4600
rect 5530 4590 5540 4600
rect 5570 4590 5600 4600
rect 5750 4590 5780 4600
rect 6030 4590 6080 4600
rect 6110 4590 6200 4600
rect 6510 4590 6560 4600
rect 7390 4590 7420 4600
rect 7470 4590 7480 4600
rect 7520 4590 7540 4600
rect 7730 4590 7740 4600
rect 7910 4590 7930 4600
rect 8080 4590 8130 4600
rect 8160 4590 8170 4600
rect 8260 4590 8280 4600
rect 8320 4590 8350 4600
rect 8530 4590 8540 4600
rect 8960 4590 8970 4600
rect 9720 4590 9730 4600
rect 0 4580 670 4590
rect 890 4580 1210 4590
rect 2810 4580 2830 4590
rect 3110 4580 3120 4590
rect 3140 4580 3220 4590
rect 3450 4580 3460 4590
rect 5220 4580 5230 4590
rect 5530 4580 5550 4590
rect 5570 4580 5600 4590
rect 5650 4580 5660 4590
rect 5760 4580 5780 4590
rect 6170 4580 6260 4590
rect 6500 4580 6550 4590
rect 7580 4580 7590 4590
rect 7610 4580 7620 4590
rect 7650 4580 7660 4590
rect 7720 4580 7740 4590
rect 7790 4580 7800 4590
rect 7840 4580 7850 4590
rect 8070 4580 8130 4590
rect 8150 4580 8160 4590
rect 8250 4580 8280 4590
rect 8320 4580 8350 4590
rect 8390 4580 8400 4590
rect 8530 4580 8550 4590
rect 8620 4580 8630 4590
rect 9710 4580 9720 4590
rect 0 4570 700 4580
rect 910 4570 1220 4580
rect 3020 4570 3040 4580
rect 3130 4570 3200 4580
rect 3220 4570 3230 4580
rect 3450 4570 3460 4580
rect 5530 4570 5550 4580
rect 5570 4570 5600 4580
rect 5760 4570 5780 4580
rect 6210 4570 6290 4580
rect 6310 4570 6320 4580
rect 6480 4570 6530 4580
rect 7470 4570 7490 4580
rect 7570 4570 7580 4580
rect 7610 4570 7620 4580
rect 7690 4570 7700 4580
rect 7710 4570 7720 4580
rect 7730 4570 7740 4580
rect 7780 4570 7830 4580
rect 8070 4570 8090 4580
rect 8130 4570 8150 4580
rect 8230 4570 8240 4580
rect 8260 4570 8280 4580
rect 8330 4570 8340 4580
rect 8390 4570 8400 4580
rect 8590 4570 8600 4580
rect 9700 4570 9710 4580
rect 0 4560 700 4570
rect 920 4560 1230 4570
rect 3030 4560 3040 4570
rect 3150 4560 3170 4570
rect 3180 4560 3200 4570
rect 3220 4560 3230 4570
rect 3250 4560 3260 4570
rect 5540 4560 5550 4570
rect 5570 4560 5600 4570
rect 5670 4560 5680 4570
rect 6210 4560 6240 4570
rect 6280 4560 6330 4570
rect 6480 4560 6520 4570
rect 7380 4560 7390 4570
rect 7480 4560 7490 4570
rect 7560 4560 7570 4570
rect 7610 4560 7620 4570
rect 7720 4560 7740 4570
rect 7780 4560 7810 4570
rect 8080 4560 8090 4570
rect 8140 4560 8160 4570
rect 8270 4560 8290 4570
rect 8390 4560 8400 4570
rect 8950 4560 8960 4570
rect 9690 4560 9700 4570
rect 0 4550 710 4560
rect 930 4550 1200 4560
rect 1210 4550 1240 4560
rect 2800 4550 2810 4560
rect 2980 4550 2990 4560
rect 3030 4550 3040 4560
rect 3050 4550 3080 4560
rect 3130 4550 3140 4560
rect 3150 4550 3160 4560
rect 3190 4550 3200 4560
rect 3210 4550 3230 4560
rect 5540 4550 5550 4560
rect 5560 4550 5580 4560
rect 5670 4550 5680 4560
rect 6210 4550 6230 4560
rect 6280 4550 6330 4560
rect 6470 4550 6520 4560
rect 7610 4550 7620 4560
rect 7720 4550 7740 4560
rect 8040 4550 8050 4560
rect 8060 4550 8080 4560
rect 8140 4550 8160 4560
rect 8260 4550 8290 4560
rect 8380 4550 8390 4560
rect 8480 4550 8490 4560
rect 8600 4550 8610 4560
rect 8950 4550 8960 4560
rect 9230 4550 9240 4560
rect 0 4540 720 4550
rect 940 4540 1170 4550
rect 2980 4540 2990 4550
rect 3050 4540 3060 4550
rect 3150 4540 3160 4550
rect 3200 4540 3230 4550
rect 3240 4540 3250 4550
rect 5540 4540 5580 4550
rect 5680 4540 5690 4550
rect 5790 4540 5800 4550
rect 6210 4540 6220 4550
rect 6280 4540 6320 4550
rect 6450 4540 6520 4550
rect 7530 4540 7540 4550
rect 7610 4540 7620 4550
rect 7710 4540 7720 4550
rect 8000 4540 8010 4550
rect 8050 4540 8060 4550
rect 8140 4540 8160 4550
rect 8250 4540 8290 4550
rect 8370 4540 8380 4550
rect 8480 4540 8490 4550
rect 0 4530 730 4540
rect 950 4530 1160 4540
rect 2970 4530 2980 4540
rect 3030 4530 3060 4540
rect 3070 4530 3080 4540
rect 3190 4530 3240 4540
rect 5240 4530 5250 4540
rect 5540 4530 5580 4540
rect 5680 4530 5690 4540
rect 5800 4530 5810 4540
rect 6270 4530 6280 4540
rect 6290 4530 6310 4540
rect 6460 4530 6510 4540
rect 7390 4530 7400 4540
rect 7910 4530 7920 4540
rect 7970 4530 8010 4540
rect 8140 4530 8160 4540
rect 8250 4530 8290 4540
rect 8480 4530 8490 4540
rect 8520 4530 8530 4540
rect 8580 4530 8590 4540
rect 8940 4530 8950 4540
rect 9670 4530 9680 4540
rect 0 4520 770 4530
rect 980 4520 1160 4530
rect 2980 4520 2990 4530
rect 3040 4520 3060 4530
rect 3070 4520 3090 4530
rect 3200 4520 3210 4530
rect 3220 4520 3240 4530
rect 5250 4520 5260 4530
rect 5540 4520 5580 4530
rect 5690 4520 5700 4530
rect 6270 4520 6300 4530
rect 6470 4520 6510 4530
rect 7480 4520 7500 4530
rect 7640 4520 7650 4530
rect 7890 4520 7900 4530
rect 7990 4520 8010 4530
rect 8140 4520 8160 4530
rect 8280 4520 8300 4530
rect 8390 4520 8400 4530
rect 9660 4520 9670 4530
rect 0 4510 680 4520
rect 690 4510 770 4520
rect 980 4510 1170 4520
rect 1180 4510 1200 4520
rect 2980 4510 3000 4520
rect 3050 4510 3060 4520
rect 3070 4510 3090 4520
rect 3210 4510 3220 4520
rect 3870 4510 3920 4520
rect 5260 4510 5270 4520
rect 5540 4510 5580 4520
rect 5770 4510 5810 4520
rect 6260 4510 6290 4520
rect 6420 4510 6510 4520
rect 7400 4510 7410 4520
rect 7830 4510 7850 4520
rect 7880 4510 7890 4520
rect 8000 4510 8010 4520
rect 8140 4510 8160 4520
rect 8240 4510 8250 4520
rect 8280 4510 8300 4520
rect 8500 4510 8510 4520
rect 9650 4510 9660 4520
rect 9990 4510 9990 4520
rect 0 4500 780 4510
rect 990 4500 1170 4510
rect 1190 4500 1200 4510
rect 2990 4500 3010 4510
rect 3410 4500 3420 4510
rect 3870 4500 3940 4510
rect 5260 4500 5270 4510
rect 5540 4500 5570 4510
rect 5710 4500 5720 4510
rect 5770 4500 5810 4510
rect 6260 4500 6290 4510
rect 6410 4500 6510 4510
rect 7340 4500 7350 4510
rect 7780 4500 7800 4510
rect 7860 4500 7890 4510
rect 8000 4500 8010 4510
rect 8150 4500 8170 4510
rect 8210 4500 8220 4510
rect 8280 4500 8300 4510
rect 8350 4500 8360 4510
rect 9220 4500 9230 4510
rect 9640 4500 9650 4510
rect 9980 4500 9990 4510
rect 0 4490 600 4500
rect 610 4490 650 4500
rect 670 4490 690 4500
rect 730 4490 770 4500
rect 1000 4490 1160 4500
rect 1180 4490 1190 4500
rect 3000 4490 3010 4500
rect 3060 4490 3090 4500
rect 3250 4490 3260 4500
rect 3860 4490 3910 4500
rect 3930 4490 3950 4500
rect 5270 4490 5280 4500
rect 5540 4490 5570 4500
rect 5760 4490 5800 4500
rect 5840 4490 5850 4500
rect 6250 4490 6280 4500
rect 6410 4490 6510 4500
rect 7340 4490 7350 4500
rect 7520 4490 7530 4500
rect 7760 4490 7770 4500
rect 7860 4490 7880 4500
rect 7930 4490 7950 4500
rect 8000 4490 8020 4500
rect 8150 4490 8170 4500
rect 8210 4490 8220 4500
rect 8290 4490 8300 4500
rect 8340 4490 8370 4500
rect 8400 4490 8410 4500
rect 9630 4490 9640 4500
rect 0 4480 590 4490
rect 610 4480 640 4490
rect 1010 4480 1140 4490
rect 1150 4480 1160 4490
rect 1170 4480 1180 4490
rect 2880 4480 2890 4490
rect 2990 4480 3000 4490
rect 3030 4480 3040 4490
rect 3050 4480 3070 4490
rect 3080 4480 3090 4490
rect 3100 4480 3110 4490
rect 3260 4480 3270 4490
rect 3860 4480 3910 4490
rect 3930 4480 3950 4490
rect 5730 4480 5740 4490
rect 5760 4480 5800 4490
rect 6400 4480 6410 4490
rect 6420 4480 6510 4490
rect 7420 4480 7430 4490
rect 7750 4480 7760 4490
rect 7860 4480 7880 4490
rect 7920 4480 7950 4490
rect 8000 4480 8020 4490
rect 8150 4480 8170 4490
rect 8210 4480 8240 4490
rect 8280 4480 8300 4490
rect 8340 4480 8370 4490
rect 9620 4480 9630 4490
rect 0 4470 580 4480
rect 600 4470 620 4480
rect 1010 4470 1100 4480
rect 1120 4470 1170 4480
rect 2990 4470 3000 4480
rect 3030 4470 3040 4480
rect 3050 4470 3080 4480
rect 3860 4470 3890 4480
rect 5320 4470 5330 4480
rect 6230 4470 6240 4480
rect 6390 4470 6400 4480
rect 6430 4470 6510 4480
rect 7340 4470 7350 4480
rect 7750 4470 7760 4480
rect 7840 4470 7850 4480
rect 7860 4470 7880 4480
rect 7930 4470 7960 4480
rect 8010 4470 8030 4480
rect 8150 4470 8170 4480
rect 8290 4470 8310 4480
rect 9610 4470 9620 4480
rect 0 4460 470 4470
rect 520 4460 580 4470
rect 590 4460 620 4470
rect 1030 4460 1130 4470
rect 1140 4460 1170 4470
rect 2990 4460 3000 4470
rect 3050 4460 3080 4470
rect 3120 4460 3130 4470
rect 3140 4460 3150 4470
rect 3170 4460 3180 4470
rect 3270 4460 3280 4470
rect 3390 4460 3400 4470
rect 3870 4460 3940 4470
rect 5780 4460 5790 4470
rect 6180 4460 6190 4470
rect 6210 4460 6220 4470
rect 6380 4460 6390 4470
rect 6430 4460 6500 4470
rect 7760 4460 7770 4470
rect 7870 4460 7880 4470
rect 7930 4460 7960 4470
rect 8010 4460 8030 4470
rect 8150 4460 8180 4470
rect 8280 4460 8290 4470
rect 8910 4460 8920 4470
rect 9210 4460 9220 4470
rect 9600 4460 9610 4470
rect 0 4450 440 4460
rect 460 4450 470 4460
rect 520 4450 570 4460
rect 600 4450 610 4460
rect 690 4450 700 4460
rect 1040 4450 1160 4460
rect 2980 4450 3000 4460
rect 3050 4450 3090 4460
rect 3120 4450 3160 4460
rect 3170 4450 3200 4460
rect 3230 4450 3250 4460
rect 3270 4450 3290 4460
rect 5780 4450 5790 4460
rect 6180 4450 6200 4460
rect 6360 4450 6380 4460
rect 6430 4450 6500 4460
rect 7790 4450 7800 4460
rect 7870 4450 7890 4460
rect 7930 4450 7960 4460
rect 8010 4450 8040 4460
rect 8150 4450 8180 4460
rect 9590 4450 9600 4460
rect 9940 4450 9950 4460
rect 0 4440 460 4450
rect 540 4440 600 4450
rect 680 4440 690 4450
rect 1060 4440 1160 4450
rect 2850 4440 2860 4450
rect 2990 4440 3000 4450
rect 3060 4440 3070 4450
rect 3090 4440 3100 4450
rect 3110 4440 3170 4450
rect 3180 4440 3190 4450
rect 3220 4440 3230 4450
rect 3240 4440 3250 4450
rect 3260 4440 3280 4450
rect 3900 4440 3910 4450
rect 4620 4440 4630 4450
rect 5770 4440 5780 4450
rect 6140 4440 6170 4450
rect 6200 4440 6210 4450
rect 6220 4440 6250 4450
rect 6340 4440 6370 4450
rect 6430 4440 6500 4450
rect 7780 4440 7800 4450
rect 7840 4440 7850 4450
rect 7880 4440 7890 4450
rect 7930 4440 7960 4450
rect 8010 4440 8040 4450
rect 8150 4440 8190 4450
rect 8230 4440 8240 4450
rect 8880 4440 8900 4450
rect 9580 4440 9590 4450
rect 9930 4440 9940 4450
rect 0 4430 450 4440
rect 500 4430 510 4440
rect 560 4430 580 4440
rect 1070 4430 1110 4440
rect 1140 4430 1170 4440
rect 2850 4430 2860 4440
rect 2980 4430 2990 4440
rect 3070 4430 3140 4440
rect 3150 4430 3170 4440
rect 3230 4430 3250 4440
rect 3280 4430 3300 4440
rect 3380 4430 3390 4440
rect 3860 4430 3910 4440
rect 3940 4430 3950 4440
rect 4610 4430 4650 4440
rect 6090 4430 6100 4440
rect 6200 4430 6250 4440
rect 6340 4430 6360 4440
rect 6440 4430 6490 4440
rect 7780 4430 7800 4440
rect 7840 4430 7850 4440
rect 7870 4430 7890 4440
rect 7930 4430 7970 4440
rect 8010 4430 8020 4440
rect 8030 4430 8040 4440
rect 8090 4430 8100 4440
rect 8150 4430 8180 4440
rect 8850 4430 8860 4440
rect 9570 4430 9580 4440
rect 9920 4430 9930 4440
rect 0 4420 290 4430
rect 310 4420 410 4430
rect 460 4420 490 4430
rect 1080 4420 1110 4430
rect 1140 4420 1150 4430
rect 2630 4420 2640 4430
rect 2750 4420 2760 4430
rect 2970 4420 2980 4430
rect 3070 4420 3100 4430
rect 3130 4420 3150 4430
rect 3160 4420 3200 4430
rect 3230 4420 3250 4430
rect 3290 4420 3310 4430
rect 3850 4420 3920 4430
rect 3940 4420 3950 4430
rect 4230 4420 4280 4430
rect 4610 4420 4670 4430
rect 4780 4420 4790 4430
rect 5300 4420 5310 4430
rect 6090 4420 6100 4430
rect 6200 4420 6250 4430
rect 6320 4420 6340 4430
rect 6350 4420 6360 4430
rect 6440 4420 6490 4430
rect 7790 4420 7800 4430
rect 7880 4420 7890 4430
rect 7940 4420 7970 4430
rect 8010 4420 8020 4430
rect 8030 4420 8050 4430
rect 8080 4420 8100 4430
rect 8110 4420 8120 4430
rect 8140 4420 8170 4430
rect 9560 4420 9570 4430
rect 9900 4420 9920 4430
rect 0 4410 280 4420
rect 320 4410 350 4420
rect 360 4410 400 4420
rect 410 4410 420 4420
rect 460 4410 480 4420
rect 1090 4410 1100 4420
rect 2740 4410 2750 4420
rect 2840 4410 2850 4420
rect 2960 4410 2970 4420
rect 3070 4410 3110 4420
rect 3130 4410 3180 4420
rect 3190 4410 3210 4420
rect 3220 4410 3240 4420
rect 3370 4410 3380 4420
rect 3830 4410 3920 4420
rect 3940 4410 3950 4420
rect 4230 4410 4300 4420
rect 4600 4410 4620 4420
rect 4660 4410 4690 4420
rect 4780 4410 4790 4420
rect 6210 4410 6250 4420
rect 6300 4410 6330 4420
rect 6440 4410 6490 4420
rect 7420 4410 7430 4420
rect 7790 4410 7810 4420
rect 7850 4410 7860 4420
rect 7880 4410 7900 4420
rect 8010 4410 8020 4420
rect 8030 4410 8040 4420
rect 8080 4410 8090 4420
rect 8120 4410 8170 4420
rect 8880 4410 8890 4420
rect 9550 4410 9560 4420
rect 9890 4410 9910 4420
rect 0 4400 280 4410
rect 330 4400 360 4410
rect 2650 4400 2660 4410
rect 2840 4400 2860 4410
rect 2870 4400 2880 4410
rect 3060 4400 3110 4410
rect 3130 4400 3180 4410
rect 3190 4400 3240 4410
rect 3290 4400 3300 4410
rect 3310 4400 3320 4410
rect 3820 4400 3910 4410
rect 3920 4400 3940 4410
rect 4240 4400 4310 4410
rect 4600 4400 4610 4410
rect 4700 4400 4710 4410
rect 6200 4400 6250 4410
rect 6290 4400 6300 4410
rect 6440 4400 6480 4410
rect 7790 4400 7810 4410
rect 7850 4400 7860 4410
rect 7890 4400 7900 4410
rect 8000 4400 8010 4410
rect 8130 4400 8170 4410
rect 8880 4400 8890 4410
rect 9870 4400 9900 4410
rect 0 4390 220 4400
rect 230 4390 260 4400
rect 350 4390 370 4400
rect 380 4390 400 4400
rect 2640 4390 2670 4400
rect 2800 4390 2810 4400
rect 2940 4390 2950 4400
rect 3070 4390 3180 4400
rect 3200 4390 3210 4400
rect 3220 4390 3240 4400
rect 3360 4390 3370 4400
rect 3820 4390 3920 4400
rect 4250 4390 4310 4400
rect 4590 4390 4610 4400
rect 4710 4390 4730 4400
rect 4820 4390 4860 4400
rect 4880 4390 4890 4400
rect 5310 4390 5320 4400
rect 6200 4390 6240 4400
rect 6280 4390 6290 4400
rect 6450 4390 6470 4400
rect 7790 4390 7810 4400
rect 7850 4390 7860 4400
rect 7890 4390 7910 4400
rect 8120 4390 8170 4400
rect 9870 4390 9890 4400
rect 0 4380 220 4390
rect 370 4380 380 4390
rect 2700 4380 2710 4390
rect 2820 4380 2840 4390
rect 2870 4380 2880 4390
rect 2930 4380 2940 4390
rect 3080 4380 3190 4390
rect 3210 4380 3220 4390
rect 3820 4380 3920 4390
rect 4260 4380 4320 4390
rect 4590 4380 4600 4390
rect 4730 4380 4740 4390
rect 4800 4380 4900 4390
rect 5950 4380 5960 4390
rect 6080 4380 6100 4390
rect 6150 4380 6160 4390
rect 6190 4380 6210 4390
rect 6270 4380 6280 4390
rect 7790 4380 7810 4390
rect 7890 4380 7900 4390
rect 7910 4380 7920 4390
rect 7980 4380 7990 4390
rect 8130 4380 8170 4390
rect 8720 4380 8730 4390
rect 8850 4380 8860 4390
rect 9190 4380 9200 4390
rect 9510 4380 9520 4390
rect 9870 4380 9880 4390
rect 0 4370 220 4380
rect 2630 4370 2640 4380
rect 2710 4370 2720 4380
rect 2820 4370 2830 4380
rect 2840 4370 2850 4380
rect 2870 4370 2880 4380
rect 2950 4370 2960 4380
rect 3090 4370 3130 4380
rect 3170 4370 3200 4380
rect 3830 4370 3930 4380
rect 4270 4370 4320 4380
rect 4580 4370 4590 4380
rect 4740 4370 4780 4380
rect 4790 4370 4840 4380
rect 4850 4370 4900 4380
rect 5330 4370 5340 4380
rect 5960 4370 5980 4380
rect 5990 4370 6050 4380
rect 6070 4370 6190 4380
rect 6220 4370 6260 4380
rect 7800 4370 7810 4380
rect 8130 4370 8170 4380
rect 8600 4370 8620 4380
rect 8720 4370 8730 4380
rect 8850 4370 8860 4380
rect 9500 4370 9510 4380
rect 0 4360 220 4370
rect 2590 4360 2600 4370
rect 2620 4360 2630 4370
rect 2700 4360 2710 4370
rect 2930 4360 2950 4370
rect 3080 4360 3090 4370
rect 3170 4360 3210 4370
rect 3220 4360 3230 4370
rect 3300 4360 3310 4370
rect 3350 4360 3360 4370
rect 3840 4360 3920 4370
rect 4280 4360 4330 4370
rect 4570 4360 4580 4370
rect 4820 4360 4900 4370
rect 5330 4360 5340 4370
rect 5980 4360 6240 4370
rect 7800 4360 7820 4370
rect 8140 4360 8170 4370
rect 8540 4360 8550 4370
rect 8590 4360 8600 4370
rect 8850 4360 8860 4370
rect 0 4350 240 4360
rect 2830 4350 2840 4360
rect 3070 4350 3080 4360
rect 3180 4350 3200 4360
rect 3230 4350 3250 4360
rect 3350 4350 3360 4360
rect 3850 4350 3900 4360
rect 4280 4350 4310 4360
rect 4570 4350 4580 4360
rect 4840 4350 4860 4360
rect 4890 4350 4920 4360
rect 5330 4350 5340 4360
rect 6080 4350 6150 4360
rect 7360 4350 7380 4360
rect 7850 4350 7860 4360
rect 8140 4350 8170 4360
rect 9850 4350 9860 4360
rect 9970 4350 9980 4360
rect 0 4340 240 4350
rect 2580 4340 2590 4350
rect 2740 4340 2750 4350
rect 2820 4340 2830 4350
rect 2920 4340 2930 4350
rect 3050 4340 3060 4350
rect 3160 4340 3210 4350
rect 3240 4340 3260 4350
rect 3300 4340 3310 4350
rect 3330 4340 3340 4350
rect 3850 4340 3860 4350
rect 4170 4340 4190 4350
rect 4200 4340 4230 4350
rect 4300 4340 4310 4350
rect 4560 4340 4570 4350
rect 4890 4340 4930 4350
rect 8140 4340 8180 4350
rect 8580 4340 8590 4350
rect 9180 4340 9190 4350
rect 9840 4340 9850 4350
rect 0 4330 80 4340
rect 90 4330 240 4340
rect 260 4330 270 4340
rect 2580 4330 2590 4340
rect 2630 4330 2640 4340
rect 2740 4330 2750 4340
rect 2920 4330 2930 4340
rect 3030 4330 3040 4340
rect 3090 4330 3100 4340
rect 3140 4330 3210 4340
rect 3240 4330 3260 4340
rect 3300 4330 3310 4340
rect 4170 4330 4240 4340
rect 4300 4330 4330 4340
rect 4560 4330 4570 4340
rect 4900 4330 4940 4340
rect 5340 4330 5350 4340
rect 7370 4330 7410 4340
rect 8140 4330 8180 4340
rect 8510 4330 8520 4340
rect 0 4320 70 4330
rect 90 4320 120 4330
rect 130 4320 270 4330
rect 2810 4320 2820 4330
rect 2840 4320 2860 4330
rect 3020 4320 3030 4330
rect 3100 4320 3110 4330
rect 3120 4320 3140 4330
rect 3190 4320 3210 4330
rect 3240 4320 3260 4330
rect 3270 4320 3280 4330
rect 3300 4320 3310 4330
rect 4150 4320 4160 4330
rect 4170 4320 4230 4330
rect 4240 4320 4260 4330
rect 4330 4320 4340 4330
rect 4550 4320 4560 4330
rect 4910 4320 4940 4330
rect 7350 4320 7360 4330
rect 8150 4320 8180 4330
rect 8430 4320 8440 4330
rect 8680 4320 8700 4330
rect 0 4310 140 4320
rect 150 4310 170 4320
rect 180 4310 210 4320
rect 230 4310 260 4320
rect 2690 4310 2700 4320
rect 2800 4310 2810 4320
rect 2820 4310 2840 4320
rect 2850 4310 2860 4320
rect 3010 4310 3020 4320
rect 3090 4310 3140 4320
rect 3200 4310 3210 4320
rect 3220 4310 3230 4320
rect 3260 4310 3280 4320
rect 4150 4310 4220 4320
rect 4250 4310 4270 4320
rect 4330 4310 4340 4320
rect 4910 4310 4940 4320
rect 5320 4310 5330 4320
rect 7330 4310 7340 4320
rect 8160 4310 8180 4320
rect 8430 4310 8440 4320
rect 9440 4310 9450 4320
rect 9920 4310 9950 4320
rect 0 4300 80 4310
rect 100 4300 120 4310
rect 2800 4300 2810 4310
rect 2820 4300 2830 4310
rect 2850 4300 2860 4310
rect 3000 4300 3010 4310
rect 3050 4300 3130 4310
rect 3180 4300 3190 4310
rect 3200 4300 3210 4310
rect 3260 4300 3290 4310
rect 4140 4300 4200 4310
rect 4270 4300 4280 4310
rect 4540 4300 4550 4310
rect 4920 4300 4950 4310
rect 5320 4300 5330 4310
rect 7260 4300 7290 4310
rect 8160 4300 8180 4310
rect 9180 4300 9190 4310
rect 9930 4300 9940 4310
rect 9950 4300 9960 4310
rect 0 4290 70 4300
rect 2560 4290 2590 4300
rect 2830 4290 2840 4300
rect 2990 4290 3000 4300
rect 3040 4290 3050 4300
rect 3060 4290 3080 4300
rect 3100 4290 3140 4300
rect 3150 4290 3160 4300
rect 3240 4290 3250 4300
rect 3260 4290 3270 4300
rect 3280 4290 3290 4300
rect 4140 4290 4180 4300
rect 4530 4290 4550 4300
rect 4920 4290 4960 4300
rect 6090 4290 6100 4300
rect 6150 4290 6170 4300
rect 7230 4290 7250 4300
rect 7350 4290 7370 4300
rect 8160 4290 8180 4300
rect 8520 4290 8530 4300
rect 8660 4290 8670 4300
rect 8730 4290 8740 4300
rect 9180 4290 9190 4300
rect 9930 4290 9950 4300
rect 0 4280 80 4290
rect 2580 4280 2590 4290
rect 2810 4280 2820 4290
rect 2910 4280 2920 4290
rect 2990 4280 3000 4290
rect 3030 4280 3040 4290
rect 3090 4280 3120 4290
rect 3130 4280 3140 4290
rect 3150 4280 3170 4290
rect 3190 4280 3210 4290
rect 3240 4280 3260 4290
rect 4130 4280 4180 4290
rect 4300 4280 4310 4290
rect 4530 4280 4540 4290
rect 4940 4280 4960 4290
rect 5350 4280 5360 4290
rect 6080 4280 6180 4290
rect 7200 4280 7220 4290
rect 8160 4280 8180 4290
rect 8710 4280 8720 4290
rect 8850 4280 8860 4290
rect 9180 4280 9190 4290
rect 9930 4280 9940 4290
rect 0 4270 80 4280
rect 2830 4270 2860 4280
rect 2870 4270 2880 4280
rect 2890 4270 2920 4280
rect 2980 4270 2990 4280
rect 3110 4270 3140 4280
rect 3160 4270 3180 4280
rect 3200 4270 3210 4280
rect 3240 4270 3260 4280
rect 3290 4270 3300 4280
rect 4140 4270 4170 4280
rect 4520 4270 4540 4280
rect 4950 4270 4980 4280
rect 7160 4270 7180 4280
rect 7200 4270 7220 4280
rect 8170 4270 8190 4280
rect 8580 4270 8590 4280
rect 9180 4270 9190 4280
rect 9810 4270 9820 4280
rect 9920 4270 9930 4280
rect 0 4260 80 4270
rect 2810 4260 2820 4270
rect 2850 4260 2860 4270
rect 2930 4260 2940 4270
rect 3020 4260 3030 4270
rect 3100 4260 3140 4270
rect 3170 4260 3180 4270
rect 3240 4260 3290 4270
rect 4140 4260 4160 4270
rect 4320 4260 4330 4270
rect 4510 4260 4520 4270
rect 4960 4260 4970 4270
rect 5460 4260 5470 4270
rect 7170 4260 7240 4270
rect 7400 4260 7420 4270
rect 8170 4260 8190 4270
rect 8440 4260 8450 4270
rect 9180 4260 9190 4270
rect 9780 4260 9790 4270
rect 9800 4260 9820 4270
rect 9860 4260 9880 4270
rect 9910 4260 9930 4270
rect 0 4250 90 4260
rect 2800 4250 2810 4260
rect 2830 4250 2850 4260
rect 2880 4250 2890 4260
rect 2930 4250 2940 4260
rect 2970 4250 2980 4260
rect 3010 4250 3030 4260
rect 3080 4250 3130 4260
rect 3150 4250 3160 4260
rect 3180 4250 3190 4260
rect 3240 4250 3280 4260
rect 4130 4250 4160 4260
rect 4330 4250 4340 4260
rect 4510 4250 4520 4260
rect 4970 4250 4990 4260
rect 5470 4250 5480 4260
rect 7080 4250 7150 4260
rect 7190 4250 7230 4260
rect 7350 4250 7370 4260
rect 7440 4250 7450 4260
rect 8170 4250 8200 4260
rect 8440 4250 8450 4260
rect 9180 4250 9190 4260
rect 9770 4250 9780 4260
rect 9860 4250 9870 4260
rect 0 4240 120 4250
rect 2540 4240 2550 4250
rect 2740 4240 2760 4250
rect 2790 4240 2800 4250
rect 2830 4240 2870 4250
rect 2890 4240 2910 4250
rect 2960 4240 2990 4250
rect 3010 4240 3070 4250
rect 3150 4240 3170 4250
rect 3190 4240 3200 4250
rect 3250 4240 3270 4250
rect 4120 4240 4160 4250
rect 4340 4240 4350 4250
rect 4490 4240 4500 4250
rect 4980 4240 5000 4250
rect 5370 4240 5380 4250
rect 5480 4240 5490 4250
rect 7090 4240 7110 4250
rect 7180 4240 7190 4250
rect 7280 4240 7290 4250
rect 7410 4240 7450 4250
rect 8160 4240 8200 4250
rect 8510 4240 8520 4250
rect 9180 4240 9190 4250
rect 9390 4240 9400 4250
rect 9850 4240 9870 4250
rect 10 4230 110 4240
rect 2510 4230 2520 4240
rect 2530 4230 2550 4240
rect 2830 4230 2870 4240
rect 2890 4230 2900 4240
rect 2960 4230 2970 4240
rect 2980 4230 2990 4240
rect 3060 4230 3070 4240
rect 3090 4230 3130 4240
rect 3150 4230 3160 4240
rect 3220 4230 3240 4240
rect 4120 4230 4140 4240
rect 4350 4230 4360 4240
rect 4480 4230 4490 4240
rect 4990 4230 5000 4240
rect 7150 4230 7170 4240
rect 7250 4230 7260 4240
rect 7370 4230 7380 4240
rect 7390 4230 7420 4240
rect 8170 4230 8200 4240
rect 8470 4230 8480 4240
rect 9180 4230 9190 4240
rect 9800 4230 9810 4240
rect 9830 4230 9870 4240
rect 9990 4230 9990 4240
rect 10 4220 110 4230
rect 2530 4220 2550 4230
rect 2600 4220 2610 4230
rect 2790 4220 2810 4230
rect 2860 4220 2890 4230
rect 2950 4220 2990 4230
rect 3010 4220 3040 4230
rect 3100 4220 3110 4230
rect 3130 4220 3140 4230
rect 3230 4220 3240 4230
rect 4110 4220 4130 4230
rect 4360 4220 4370 4230
rect 4460 4220 4490 4230
rect 4990 4220 5010 4230
rect 5490 4220 5500 4230
rect 7130 4220 7140 4230
rect 7210 4220 7220 4230
rect 8160 4220 8200 4230
rect 8830 4220 8840 4230
rect 9950 4220 9980 4230
rect 20 4210 130 4220
rect 2800 4210 2810 4220
rect 2840 4210 2890 4220
rect 2910 4210 2970 4220
rect 3000 4210 3030 4220
rect 3150 4210 3160 4220
rect 3170 4210 3180 4220
rect 3210 4210 3220 4220
rect 3230 4210 3240 4220
rect 3250 4210 3260 4220
rect 4110 4210 4130 4220
rect 4360 4210 4370 4220
rect 4450 4210 4470 4220
rect 5000 4210 5010 4220
rect 5500 4210 5530 4220
rect 7300 4210 7340 4220
rect 7460 4210 7470 4220
rect 8170 4210 8200 4220
rect 9320 4210 9330 4220
rect 9970 4210 9990 4220
rect 60 4200 120 4210
rect 2780 4200 2790 4210
rect 2950 4200 2960 4210
rect 3010 4200 3030 4210
rect 3100 4200 3140 4210
rect 3160 4200 3170 4210
rect 3210 4200 3230 4210
rect 4110 4200 4120 4210
rect 4360 4200 4390 4210
rect 4440 4200 4450 4210
rect 5000 4200 5010 4210
rect 5390 4200 5410 4210
rect 5500 4200 5540 4210
rect 8180 4200 8210 4210
rect 9760 4200 9770 4210
rect 9970 4200 9980 4210
rect 9990 4200 9990 4210
rect 0 4190 10 4200
rect 70 4190 130 4200
rect 150 4190 200 4200
rect 2550 4190 2560 4200
rect 2570 4190 2600 4200
rect 2650 4190 2660 4200
rect 2760 4190 2790 4200
rect 2870 4190 2910 4200
rect 2990 4190 3050 4200
rect 3080 4190 3150 4200
rect 3210 4190 3230 4200
rect 3240 4190 3250 4200
rect 4100 4190 4120 4200
rect 4380 4190 4400 4200
rect 4440 4190 4450 4200
rect 5010 4190 5020 4200
rect 5490 4190 5500 4200
rect 5510 4190 5550 4200
rect 7230 4190 7260 4200
rect 7470 4190 7480 4200
rect 8180 4190 8200 4200
rect 9790 4190 9800 4200
rect 9810 4190 9820 4200
rect 9880 4190 9900 4200
rect 0 4180 20 4190
rect 30 4180 40 4190
rect 80 4180 130 4190
rect 2570 4180 2590 4190
rect 2600 4180 2610 4190
rect 2640 4180 2660 4190
rect 2760 4180 2790 4190
rect 2820 4180 2860 4190
rect 2890 4180 2930 4190
rect 3000 4180 3020 4190
rect 3080 4180 3090 4190
rect 3130 4180 3140 4190
rect 3170 4180 3190 4190
rect 3200 4180 3220 4190
rect 3230 4180 3240 4190
rect 4100 4180 4110 4190
rect 4440 4180 4450 4190
rect 5020 4180 5030 4190
rect 5390 4180 5400 4190
rect 5490 4180 5500 4190
rect 5540 4180 5560 4190
rect 7290 4180 7310 4190
rect 7470 4180 7480 4190
rect 8180 4180 8210 4190
rect 9180 4180 9190 4190
rect 9290 4180 9310 4190
rect 9810 4180 9840 4190
rect 0 4170 30 4180
rect 70 4170 130 4180
rect 2570 4170 2590 4180
rect 2630 4170 2660 4180
rect 2670 4170 2690 4180
rect 2700 4170 2710 4180
rect 2760 4170 2790 4180
rect 2810 4170 2840 4180
rect 2870 4170 2900 4180
rect 2940 4170 2950 4180
rect 3000 4170 3020 4180
rect 3170 4170 3200 4180
rect 3220 4170 3230 4180
rect 4090 4170 4100 4180
rect 4410 4170 4440 4180
rect 5020 4170 5030 4180
rect 5380 4170 5390 4180
rect 5490 4170 5500 4180
rect 5540 4170 5570 4180
rect 7310 4170 7330 4180
rect 7470 4170 7480 4180
rect 8180 4170 8210 4180
rect 9290 4170 9310 4180
rect 9820 4170 9830 4180
rect 9860 4170 9870 4180
rect 0 4160 30 4170
rect 60 4160 130 4170
rect 2580 4160 2610 4170
rect 2650 4160 2660 4170
rect 2680 4160 2780 4170
rect 2810 4160 2840 4170
rect 2850 4160 2860 4170
rect 2870 4160 2890 4170
rect 2950 4160 2970 4170
rect 2990 4160 3010 4170
rect 3130 4160 3170 4170
rect 3180 4160 3190 4170
rect 4090 4160 4100 4170
rect 5030 4160 5040 4170
rect 5400 4160 5410 4170
rect 5560 4160 5580 4170
rect 7260 4160 7270 4170
rect 7310 4160 7340 4170
rect 8190 4160 8200 4170
rect 9830 4160 9840 4170
rect 9870 4160 9880 4170
rect 10 4150 40 4160
rect 50 4150 110 4160
rect 2580 4150 2620 4160
rect 2670 4150 2690 4160
rect 2700 4150 2730 4160
rect 2740 4150 2760 4160
rect 2770 4150 2780 4160
rect 2810 4150 2860 4160
rect 2880 4150 2900 4160
rect 2920 4150 2930 4160
rect 2970 4150 3010 4160
rect 3090 4150 3120 4160
rect 3170 4150 3180 4160
rect 3200 4150 3210 4160
rect 3230 4150 3240 4160
rect 4080 4150 4100 4160
rect 5030 4150 5040 4160
rect 5490 4150 5500 4160
rect 5570 4150 5590 4160
rect 7250 4150 7260 4160
rect 7350 4150 7360 4160
rect 9280 4150 9290 4160
rect 9850 4150 9860 4160
rect 9880 4150 9890 4160
rect 50 4140 150 4150
rect 2580 4140 2590 4150
rect 2600 4140 2630 4150
rect 2670 4140 2680 4150
rect 2690 4140 2720 4150
rect 2740 4140 2790 4150
rect 2810 4140 2870 4150
rect 2880 4140 2900 4150
rect 2920 4140 2930 4150
rect 2970 4140 3040 4150
rect 3090 4140 3110 4150
rect 3140 4140 3150 4150
rect 3190 4140 3230 4150
rect 3280 4140 3290 4150
rect 4080 4140 4090 4150
rect 5040 4140 5060 4150
rect 5430 4140 5440 4150
rect 5590 4140 5600 4150
rect 7370 4140 7380 4150
rect 8200 4140 8210 4150
rect 8810 4140 8820 4150
rect 9870 4140 9880 4150
rect 60 4130 150 4140
rect 2480 4130 2490 4140
rect 2580 4130 2620 4140
rect 2680 4130 2790 4140
rect 2810 4130 2900 4140
rect 2910 4130 2950 4140
rect 2990 4130 3020 4140
rect 3040 4130 3060 4140
rect 3070 4130 3120 4140
rect 3170 4130 3190 4140
rect 3210 4130 3220 4140
rect 3230 4130 3260 4140
rect 4760 4130 4800 4140
rect 4880 4130 4920 4140
rect 5040 4130 5090 4140
rect 5600 4130 5610 4140
rect 7390 4130 7420 4140
rect 7460 4130 7480 4140
rect 8200 4130 8210 4140
rect 9880 4130 9890 4140
rect 9940 4130 9950 4140
rect 90 4120 120 4130
rect 130 4120 150 4130
rect 2590 4120 2630 4130
rect 2680 4120 2790 4130
rect 2820 4120 2870 4130
rect 2880 4120 2970 4130
rect 2990 4120 3000 4130
rect 3010 4120 3020 4130
rect 3070 4120 3160 4130
rect 3200 4120 3210 4130
rect 3220 4120 3240 4130
rect 4070 4120 4080 4130
rect 4730 4120 4760 4130
rect 4920 4120 4950 4130
rect 5030 4120 5100 4130
rect 5610 4120 5620 4130
rect 7240 4120 7250 4130
rect 8200 4120 8210 4130
rect 9890 4120 9900 4130
rect 9950 4120 9960 4130
rect 90 4110 150 4120
rect 2600 4110 2640 4120
rect 2680 4110 2790 4120
rect 2810 4110 2840 4120
rect 2860 4110 2870 4120
rect 2890 4110 2970 4120
rect 3000 4110 3020 4120
rect 3080 4110 3130 4120
rect 3180 4110 3210 4120
rect 4070 4110 4080 4120
rect 4710 4110 4730 4120
rect 4940 4110 5030 4120
rect 5080 4110 5110 4120
rect 5620 4110 5630 4120
rect 7430 4110 7440 4120
rect 9910 4110 9920 4120
rect 9960 4110 9970 4120
rect 100 4100 150 4110
rect 2610 4100 2650 4110
rect 2680 4100 2790 4110
rect 2820 4100 2830 4110
rect 2840 4100 2860 4110
rect 2870 4100 2960 4110
rect 3010 4100 3090 4110
rect 3170 4100 3200 4110
rect 4670 4100 4700 4110
rect 4920 4100 5010 4110
rect 5080 4100 5120 4110
rect 5630 4100 5640 4110
rect 7450 4100 7470 4110
rect 7480 4100 7490 4110
rect 8800 4100 8810 4110
rect 9920 4100 9930 4110
rect 9980 4100 9990 4110
rect 110 4090 150 4100
rect 2610 4090 2800 4100
rect 2810 4090 2820 4100
rect 2840 4090 2950 4100
rect 2960 4090 2970 4100
rect 3010 4090 3030 4100
rect 3050 4090 3060 4100
rect 3070 4090 3190 4100
rect 4060 4090 4070 4100
rect 4670 4090 4680 4100
rect 4890 4090 4900 4100
rect 5090 4090 5130 4100
rect 5640 4090 5660 4100
rect 7470 4090 7480 4100
rect 7510 4090 7520 4100
rect 9940 4090 9950 4100
rect 9990 4090 9990 4100
rect 110 4080 140 4090
rect 2600 4080 2610 4090
rect 2620 4080 2800 4090
rect 2820 4080 2830 4090
rect 2850 4080 2970 4090
rect 2990 4080 3020 4090
rect 3030 4080 3070 4090
rect 4650 4080 4670 4090
rect 5100 4080 5130 4090
rect 5660 4080 5670 4090
rect 7570 4080 7580 4090
rect 8790 4080 8800 4090
rect 9210 4080 9220 4090
rect 9950 4080 9970 4090
rect 130 4070 150 4080
rect 2610 4070 2650 4080
rect 2660 4070 2810 4080
rect 2820 4070 2830 4080
rect 2880 4070 3020 4080
rect 3050 4070 3060 4080
rect 3080 4070 3090 4080
rect 3270 4070 3280 4080
rect 4050 4070 4060 4080
rect 4640 4070 4660 4080
rect 5110 4070 5140 4080
rect 5660 4070 5670 4080
rect 7550 4070 7560 4080
rect 8730 4070 8750 4080
rect 8770 4070 8790 4080
rect 9970 4070 9980 4080
rect 140 4060 160 4070
rect 2620 4060 2650 4070
rect 2660 4060 2810 4070
rect 2820 4060 2840 4070
rect 2850 4060 2870 4070
rect 2880 4060 2930 4070
rect 2950 4060 3010 4070
rect 3080 4060 3090 4070
rect 3110 4060 3130 4070
rect 4640 4060 4650 4070
rect 4810 4060 4820 4070
rect 5110 4060 5140 4070
rect 5670 4060 5680 4070
rect 7640 4060 7650 4070
rect 8730 4060 8750 4070
rect 8760 4060 8770 4070
rect 9990 4060 9990 4070
rect 2620 4050 2820 4060
rect 2830 4050 2850 4060
rect 2870 4050 2940 4060
rect 2950 4050 2970 4060
rect 2990 4050 3010 4060
rect 3120 4050 3150 4060
rect 3270 4050 3280 4060
rect 4040 4050 4050 4060
rect 4630 4050 4640 4060
rect 5110 4050 5150 4060
rect 5500 4050 5510 4060
rect 5690 4050 5700 4060
rect 8660 4050 8670 4060
rect 8690 4050 8700 4060
rect 8750 4050 8770 4060
rect 150 4040 160 4050
rect 2620 4040 2870 4050
rect 2880 4040 2960 4050
rect 2990 4040 3030 4050
rect 3150 4040 3170 4050
rect 4030 4040 4040 4050
rect 4630 4040 4640 4050
rect 4780 4040 4790 4050
rect 5110 4040 5150 4050
rect 5410 4040 5420 4050
rect 5500 4040 5510 4050
rect 5700 4040 5710 4050
rect 7690 4040 7700 4050
rect 8580 4040 8620 4050
rect 8760 4040 8770 4050
rect 150 4030 160 4040
rect 2600 4030 2640 4040
rect 2650 4030 2770 4040
rect 2820 4030 2870 4040
rect 2880 4030 2950 4040
rect 2980 4030 3050 4040
rect 3160 4030 3170 4040
rect 3270 4030 3280 4040
rect 4030 4030 4040 4040
rect 4620 4030 4630 4040
rect 4760 4030 4770 4040
rect 5110 4030 5160 4040
rect 5500 4030 5510 4040
rect 5710 4030 5720 4040
rect 7200 4030 7210 4040
rect 7670 4030 7690 4040
rect 8620 4030 8630 4040
rect 8730 4030 8750 4040
rect 150 4020 180 4030
rect 2600 4020 2770 4030
rect 2790 4020 2810 4030
rect 2820 4020 2870 4030
rect 2880 4020 2950 4030
rect 2980 4020 3060 4030
rect 3270 4020 3280 4030
rect 4620 4020 4630 4030
rect 5120 4020 5160 4030
rect 5500 4020 5510 4030
rect 5720 4020 5730 4030
rect 7700 4020 7710 4030
rect 7740 4020 7750 4030
rect 8480 4020 8500 4030
rect 8680 4020 8690 4030
rect 8730 4020 8740 4030
rect 160 4010 180 4020
rect 2590 4010 2780 4020
rect 2790 4010 2950 4020
rect 2980 4010 3070 4020
rect 3170 4010 3180 4020
rect 3270 4010 3280 4020
rect 4020 4010 4030 4020
rect 4620 4010 4630 4020
rect 4730 4010 4740 4020
rect 5130 4010 5160 4020
rect 5500 4010 5510 4020
rect 5730 4010 5740 4020
rect 7720 4010 7730 4020
rect 8530 4010 8540 4020
rect 8700 4010 8710 4020
rect 8760 4010 8770 4020
rect 160 4000 180 4010
rect 2600 4000 2770 4010
rect 2790 4000 2840 4010
rect 2850 4000 2950 4010
rect 2980 4000 3080 4010
rect 4010 4000 4030 4010
rect 5140 4000 5170 4010
rect 5500 4000 5510 4010
rect 5740 4000 5760 4010
rect 7790 4000 7800 4010
rect 8390 4000 8400 4010
rect 8430 4000 8440 4010
rect 8520 4000 8530 4010
rect 8540 4000 8560 4010
rect 8690 4000 8700 4010
rect 8720 4000 8730 4010
rect 2610 3990 2770 4000
rect 2800 3990 2840 4000
rect 2850 3990 2950 4000
rect 2970 3990 3090 4000
rect 4000 3990 4010 4000
rect 4680 3990 4690 4000
rect 5150 3990 5170 4000
rect 5500 3990 5510 4000
rect 5760 3990 5780 4000
rect 6300 3990 6310 4000
rect 7180 3990 7190 4000
rect 8340 3990 8350 4000
rect 8400 3990 8410 4000
rect 8430 3990 8440 4000
rect 8490 3990 8500 4000
rect 8670 3990 8680 4000
rect 8700 3990 8710 4000
rect 2610 3980 2770 3990
rect 2800 3980 2950 3990
rect 2970 3980 3100 3990
rect 3130 3980 3140 3990
rect 3270 3980 3280 3990
rect 4000 3980 4010 3990
rect 4820 3980 4840 3990
rect 5150 3980 5180 3990
rect 5780 3980 5800 3990
rect 6280 3980 6310 3990
rect 7800 3980 7810 3990
rect 7840 3980 7850 3990
rect 8310 3980 8330 3990
rect 8410 3980 8430 3990
rect 8500 3980 8520 3990
rect 8550 3980 8570 3990
rect 8710 3980 8720 3990
rect 2610 3970 2890 3980
rect 2900 3970 2950 3980
rect 2970 3970 3130 3980
rect 3180 3970 3190 3980
rect 3270 3970 3280 3980
rect 3980 3970 4000 3980
rect 4640 3970 4650 3980
rect 4790 3970 4830 3980
rect 5150 3970 5180 3980
rect 5490 3970 5500 3980
rect 5790 3970 5830 3980
rect 5860 3970 5870 3980
rect 5890 3970 5900 3980
rect 5930 3970 5950 3980
rect 6260 3970 6310 3980
rect 7170 3970 7180 3980
rect 7820 3970 7830 3980
rect 7870 3970 7880 3980
rect 8240 3970 8280 3980
rect 8300 3970 8310 3980
rect 8410 3970 8420 3980
rect 8540 3970 8550 3980
rect 8720 3970 8740 3980
rect 2610 3960 2890 3970
rect 2900 3960 2950 3970
rect 2970 3960 3130 3970
rect 3270 3960 3280 3970
rect 3960 3960 3990 3970
rect 4770 3960 4790 3970
rect 5160 3960 5200 3970
rect 5490 3960 5500 3970
rect 5820 3960 6000 3970
rect 6230 3960 6240 3970
rect 6250 3960 6310 3970
rect 7850 3960 7860 3970
rect 8200 3960 8220 3970
rect 8280 3960 8320 3970
rect 8410 3960 8430 3970
rect 8520 3960 8530 3970
rect 2610 3950 2820 3960
rect 2830 3950 2940 3960
rect 2970 3950 3120 3960
rect 3270 3950 3280 3960
rect 3950 3950 3980 3960
rect 4750 3950 4760 3960
rect 5170 3950 5210 3960
rect 5490 3950 5500 3960
rect 5860 3950 6040 3960
rect 6060 3950 6140 3960
rect 6150 3950 6320 3960
rect 7910 3950 7920 3960
rect 8160 3950 8170 3960
rect 8320 3950 8330 3960
rect 8410 3950 8420 3960
rect 8520 3950 8540 3960
rect 2610 3940 2950 3950
rect 2970 3940 3110 3950
rect 3270 3940 3280 3950
rect 3930 3940 3950 3950
rect 5180 3940 5220 3950
rect 5410 3940 5420 3950
rect 5490 3940 5500 3950
rect 5910 3940 5920 3950
rect 5960 3940 6320 3950
rect 7900 3940 7910 3950
rect 8120 3940 8130 3950
rect 8520 3940 8530 3950
rect 8540 3940 8550 3950
rect 8570 3940 8580 3950
rect 9690 3940 9700 3950
rect 2610 3930 2930 3940
rect 2970 3930 3050 3940
rect 3060 3930 3120 3940
rect 3170 3930 3180 3940
rect 3270 3930 3280 3940
rect 3910 3930 3940 3940
rect 4200 3930 4250 3940
rect 4260 3930 4270 3940
rect 5190 3930 5220 3940
rect 5420 3930 5490 3940
rect 6010 3930 6320 3940
rect 8100 3930 8110 3940
rect 8330 3930 8340 3940
rect 8420 3930 8430 3940
rect 8450 3930 8460 3940
rect 8510 3930 8520 3940
rect 8530 3930 8540 3940
rect 8630 3930 8640 3940
rect 9650 3930 9660 3940
rect 9680 3930 9690 3940
rect 2610 3920 2930 3930
rect 2960 3920 3020 3930
rect 3060 3920 3100 3930
rect 3160 3920 3180 3930
rect 3210 3920 3220 3930
rect 3260 3920 3280 3930
rect 3910 3920 3920 3930
rect 4160 3920 4170 3930
rect 4190 3920 4260 3930
rect 5200 3920 5230 3930
rect 5420 3920 5440 3930
rect 5460 3920 5480 3930
rect 6050 3920 6080 3930
rect 6090 3920 6130 3930
rect 6160 3920 6320 3930
rect 6330 3920 6340 3930
rect 7940 3920 7950 3930
rect 7970 3920 7980 3930
rect 8090 3920 8120 3930
rect 8130 3920 8140 3930
rect 8680 3920 8690 3930
rect 9640 3920 9660 3930
rect 9720 3920 9730 3930
rect 2610 3910 2860 3920
rect 2880 3910 2940 3920
rect 2960 3910 3030 3920
rect 3150 3910 3170 3920
rect 3200 3910 3220 3920
rect 3260 3910 3280 3920
rect 3900 3910 3910 3920
rect 4190 3910 4270 3920
rect 5200 3910 5230 3920
rect 5420 3910 5440 3920
rect 6160 3910 6330 3920
rect 7950 3910 7960 3920
rect 8060 3910 8070 3920
rect 8100 3910 8110 3920
rect 8120 3910 8140 3920
rect 8180 3910 8190 3920
rect 8280 3910 8310 3920
rect 8560 3910 8590 3920
rect 8650 3910 8660 3920
rect 9650 3910 9670 3920
rect 9710 3910 9730 3920
rect 9740 3910 9750 3920
rect 2590 3900 2860 3910
rect 2920 3900 2940 3910
rect 2960 3900 3030 3910
rect 3140 3900 3170 3910
rect 3200 3900 3220 3910
rect 3270 3900 3280 3910
rect 3900 3900 3910 3910
rect 4140 3900 4290 3910
rect 5220 3900 5230 3910
rect 6000 3900 6010 3910
rect 6140 3900 6330 3910
rect 7970 3900 7980 3910
rect 8280 3900 8300 3910
rect 8320 3900 8330 3910
rect 8590 3900 8600 3910
rect 8650 3900 8670 3910
rect 8700 3900 8710 3910
rect 9650 3900 9660 3910
rect 9740 3900 9760 3910
rect 2570 3890 2810 3900
rect 2820 3890 2860 3900
rect 2920 3890 2940 3900
rect 2960 3890 3000 3900
rect 3120 3890 3150 3900
rect 3270 3890 3280 3900
rect 3890 3890 3900 3900
rect 4110 3890 4300 3900
rect 5220 3890 5240 3900
rect 6020 3890 6030 3900
rect 6040 3890 6330 3900
rect 7970 3890 8000 3900
rect 8070 3890 8080 3900
rect 8280 3890 8300 3900
rect 8510 3890 8520 3900
rect 8550 3890 8560 3900
rect 8600 3890 8610 3900
rect 8620 3890 8640 3900
rect 9590 3890 9610 3900
rect 9640 3890 9650 3900
rect 9730 3890 9740 3900
rect 2550 3880 2860 3890
rect 2920 3880 2930 3890
rect 2980 3880 3010 3890
rect 3090 3880 3110 3890
rect 3120 3880 3130 3890
rect 3270 3880 3280 3890
rect 4110 3880 4300 3890
rect 5220 3880 5240 3890
rect 6040 3880 6340 3890
rect 7970 3880 8010 3890
rect 8290 3880 8310 3890
rect 8320 3880 8330 3890
rect 8520 3880 8560 3890
rect 8570 3880 8580 3890
rect 8600 3880 8610 3890
rect 9480 3880 9490 3890
rect 9550 3880 9560 3890
rect 2530 3870 2870 3880
rect 2980 3870 2990 3880
rect 3070 3870 3100 3880
rect 3110 3870 3120 3880
rect 3880 3870 3890 3880
rect 4110 3870 4310 3880
rect 5230 3870 5250 3880
rect 5990 3870 6000 3880
rect 6020 3870 6040 3880
rect 6060 3870 6340 3880
rect 7970 3870 8010 3880
rect 8020 3870 8030 3880
rect 8210 3870 8220 3880
rect 8300 3870 8320 3880
rect 8430 3870 8440 3880
rect 8460 3870 8470 3880
rect 8530 3870 8540 3880
rect 8670 3870 8690 3880
rect 9480 3870 9490 3880
rect 9800 3870 9810 3880
rect 9830 3870 9840 3880
rect 2230 3860 2300 3870
rect 2430 3860 2460 3870
rect 2540 3860 2800 3870
rect 2820 3860 2880 3870
rect 3070 3860 3100 3870
rect 3150 3860 3160 3870
rect 4110 3860 4300 3870
rect 5230 3860 5250 3870
rect 5990 3860 6310 3870
rect 6320 3860 6340 3870
rect 7980 3860 8010 3870
rect 8030 3860 8040 3870
rect 8210 3860 8220 3870
rect 8430 3860 8440 3870
rect 9440 3860 9450 3870
rect 9520 3860 9530 3870
rect 9550 3860 9560 3870
rect 9810 3860 9820 3870
rect 9850 3860 9860 3870
rect 2020 3850 2050 3860
rect 2230 3850 2290 3860
rect 2310 3850 2330 3860
rect 2390 3850 2460 3860
rect 2540 3850 2880 3860
rect 3050 3850 3070 3860
rect 3170 3850 3180 3860
rect 3870 3850 3880 3860
rect 4120 3850 4180 3860
rect 4230 3850 4280 3860
rect 5240 3850 5250 3860
rect 5980 3850 6340 3860
rect 7110 3850 7120 3860
rect 7980 3850 8010 3860
rect 8040 3850 8070 3860
rect 8210 3850 8230 3860
rect 9430 3850 9460 3860
rect 9570 3850 9580 3860
rect 9800 3850 9810 3860
rect 9860 3850 9870 3860
rect 2020 3840 2040 3850
rect 2240 3840 2300 3850
rect 2320 3840 2340 3850
rect 2400 3840 2470 3850
rect 2570 3840 2890 3850
rect 3030 3840 3060 3850
rect 3140 3840 3150 3850
rect 3860 3840 3870 3850
rect 4120 3840 4150 3850
rect 4250 3840 4280 3850
rect 5240 3840 5260 3850
rect 5970 3840 5980 3850
rect 5990 3840 6340 3850
rect 7990 3840 8020 3850
rect 8060 3840 8080 3850
rect 8210 3840 8230 3850
rect 9580 3840 9590 3850
rect 9720 3840 9730 3850
rect 2040 3830 2050 3840
rect 2410 3830 2470 3840
rect 2580 3830 2690 3840
rect 2700 3830 2900 3840
rect 2940 3830 2950 3840
rect 2980 3830 3040 3840
rect 3100 3830 3120 3840
rect 3140 3830 3150 3840
rect 3860 3830 3870 3840
rect 4100 3830 4130 3840
rect 4280 3830 4290 3840
rect 5250 3830 5260 3840
rect 5980 3830 6340 3840
rect 7100 3830 7110 3840
rect 8000 3830 8020 3840
rect 8080 3830 8100 3840
rect 8170 3830 8220 3840
rect 8470 3830 8490 3840
rect 9600 3830 9610 3840
rect 9720 3830 9730 3840
rect 9840 3830 9850 3840
rect 2420 3820 2450 3830
rect 2590 3820 2690 3830
rect 2700 3820 2890 3830
rect 2940 3820 2970 3830
rect 2980 3820 3000 3830
rect 3070 3820 3120 3830
rect 3140 3820 3160 3830
rect 3270 3820 3280 3830
rect 3850 3820 3870 3830
rect 4090 3820 4110 3830
rect 5980 3820 6310 3830
rect 8010 3820 8020 3830
rect 8070 3820 8090 3830
rect 8100 3820 8120 3830
rect 8170 3820 8220 3830
rect 8490 3820 8500 3830
rect 8610 3820 8630 3830
rect 9730 3820 9740 3830
rect 9800 3820 9820 3830
rect 2600 3810 2700 3820
rect 2710 3810 2950 3820
rect 2970 3810 2980 3820
rect 3130 3810 3160 3820
rect 3860 3810 3870 3820
rect 4080 3810 4090 3820
rect 4290 3810 4300 3820
rect 5260 3810 5270 3820
rect 5970 3810 6300 3820
rect 8080 3810 8090 3820
rect 8130 3810 8140 3820
rect 8170 3810 8180 3820
rect 8190 3810 8220 3820
rect 8500 3810 8520 3820
rect 8620 3810 8630 3820
rect 8640 3810 8650 3820
rect 9750 3810 9760 3820
rect 9770 3810 9780 3820
rect 9810 3810 9820 3820
rect 2620 3800 2700 3810
rect 2720 3800 2900 3810
rect 2920 3800 2960 3810
rect 3130 3800 3150 3810
rect 3160 3800 3200 3810
rect 3260 3800 3280 3810
rect 3860 3800 3870 3810
rect 4060 3800 4070 3810
rect 4290 3800 4300 3810
rect 5960 3800 6300 3810
rect 8020 3800 8030 3810
rect 8140 3800 8150 3810
rect 8290 3800 8300 3810
rect 8450 3800 8470 3810
rect 2540 3790 2560 3800
rect 2600 3790 2610 3800
rect 2620 3790 2700 3800
rect 2720 3790 2730 3800
rect 2740 3790 2810 3800
rect 2820 3790 2900 3800
rect 2920 3790 2940 3800
rect 3160 3790 3200 3800
rect 3270 3790 3290 3800
rect 3870 3790 3880 3800
rect 4050 3790 4060 3800
rect 5270 3790 5280 3800
rect 5970 3790 6300 3800
rect 8020 3790 8030 3800
rect 8110 3790 8120 3800
rect 8180 3790 8190 3800
rect 8200 3790 8250 3800
rect 8260 3790 8270 3800
rect 8460 3790 8470 3800
rect 8480 3790 8490 3800
rect 9750 3790 9760 3800
rect 2530 3780 2570 3790
rect 2620 3780 2940 3790
rect 3150 3780 3200 3790
rect 3270 3780 3290 3790
rect 3870 3780 3890 3790
rect 4030 3780 4050 3790
rect 4240 3780 4250 3790
rect 5270 3780 5280 3790
rect 5980 3780 6300 3790
rect 8020 3780 8030 3790
rect 8120 3780 8130 3790
rect 8150 3780 8160 3790
rect 8190 3780 8230 3790
rect 8470 3780 8480 3790
rect 1700 3770 1720 3780
rect 2540 3770 2580 3780
rect 2630 3770 2930 3780
rect 3130 3770 3190 3780
rect 3270 3770 3280 3780
rect 3290 3770 3300 3780
rect 3870 3770 3890 3780
rect 4020 3770 4040 3780
rect 5280 3770 5290 3780
rect 6010 3770 6050 3780
rect 6060 3770 6310 3780
rect 8150 3770 8160 3780
rect 8180 3770 8190 3780
rect 8330 3770 8360 3780
rect 8490 3770 8510 3780
rect 9720 3770 9730 3780
rect 9800 3770 9820 3780
rect 9840 3770 9850 3780
rect 1680 3760 1720 3770
rect 2550 3760 2590 3770
rect 2640 3760 2930 3770
rect 3130 3760 3190 3770
rect 3280 3760 3290 3770
rect 3880 3760 3900 3770
rect 4010 3760 4020 3770
rect 4180 3760 4190 3770
rect 5280 3760 5290 3770
rect 6000 3760 6010 3770
rect 6020 3760 6320 3770
rect 8140 3760 8150 3770
rect 8320 3760 8370 3770
rect 8510 3760 8530 3770
rect 9650 3760 9660 3770
rect 9710 3760 9720 3770
rect 9740 3760 9750 3770
rect 9860 3760 9870 3770
rect 1660 3750 1720 3760
rect 2560 3750 2600 3760
rect 2650 3750 2730 3760
rect 2740 3750 2770 3760
rect 2780 3750 2850 3760
rect 2870 3750 2900 3760
rect 3120 3750 3190 3760
rect 3280 3750 3290 3760
rect 3880 3750 3890 3760
rect 4000 3750 4010 3760
rect 4140 3750 4150 3760
rect 5290 3750 5300 3760
rect 6020 3750 6330 3760
rect 6350 3750 6360 3760
rect 6370 3750 6440 3760
rect 8320 3750 8360 3760
rect 8370 3750 8380 3760
rect 8530 3750 8540 3760
rect 9710 3750 9730 3760
rect 9750 3750 9760 3760
rect 9780 3750 9790 3760
rect 9850 3750 9860 3760
rect 1640 3740 1710 3750
rect 2560 3740 2600 3750
rect 2670 3740 2850 3750
rect 2860 3740 2890 3750
rect 3120 3740 3190 3750
rect 3300 3740 3310 3750
rect 3880 3740 3890 3750
rect 3990 3740 4000 3750
rect 4090 3740 4100 3750
rect 5290 3740 5300 3750
rect 6040 3740 6350 3750
rect 6360 3740 6440 3750
rect 8180 3740 8210 3750
rect 8310 3740 8350 3750
rect 8380 3740 8390 3750
rect 9680 3740 9690 3750
rect 9780 3740 9800 3750
rect 9850 3740 9870 3750
rect 1630 3730 1700 3740
rect 2570 3730 2600 3740
rect 2680 3730 2710 3740
rect 2740 3730 2890 3740
rect 3150 3730 3180 3740
rect 3280 3730 3290 3740
rect 3300 3730 3310 3740
rect 3880 3730 3890 3740
rect 3980 3730 3990 3740
rect 5290 3730 5300 3740
rect 6070 3730 6440 3740
rect 8310 3730 8350 3740
rect 8380 3730 8390 3740
rect 8540 3730 8570 3740
rect 9690 3730 9700 3740
rect 9780 3730 9800 3740
rect 9810 3730 9830 3740
rect 9930 3730 9960 3740
rect 1610 3720 1690 3730
rect 2580 3720 2590 3730
rect 2770 3720 2880 3730
rect 3280 3720 3290 3730
rect 3300 3720 3310 3730
rect 3870 3720 3890 3730
rect 3970 3720 3990 3730
rect 6070 3720 6450 3730
rect 8170 3720 8180 3730
rect 8330 3720 8360 3730
rect 8370 3720 8410 3730
rect 8540 3720 8590 3730
rect 9910 3720 9920 3730
rect 1620 3710 1680 3720
rect 2860 3710 2880 3720
rect 2970 3710 2990 3720
rect 3120 3710 3130 3720
rect 3280 3710 3290 3720
rect 3870 3710 3880 3720
rect 3960 3710 3980 3720
rect 5300 3710 5310 3720
rect 6070 3710 6450 3720
rect 8180 3710 8190 3720
rect 8390 3710 8410 3720
rect 8550 3710 8580 3720
rect 9950 3710 9960 3720
rect 0 3700 10 3710
rect 1620 3700 1710 3710
rect 2870 3700 2900 3710
rect 2950 3700 3000 3710
rect 3010 3700 3020 3710
rect 3310 3700 3320 3710
rect 3870 3700 3880 3710
rect 3960 3700 3970 3710
rect 4010 3700 4020 3710
rect 5300 3700 5310 3710
rect 6070 3700 6450 3710
rect 7010 3700 7020 3710
rect 8390 3700 8400 3710
rect 8410 3700 8440 3710
rect 8550 3700 8580 3710
rect 0 3690 30 3700
rect 1610 3690 1690 3700
rect 1700 3690 1710 3700
rect 2850 3690 2900 3700
rect 2940 3690 3040 3700
rect 3310 3690 3320 3700
rect 3870 3690 3880 3700
rect 4190 3690 4200 3700
rect 4870 3690 4900 3700
rect 6070 3690 6470 3700
rect 8390 3690 8400 3700
rect 8450 3690 8470 3700
rect 8560 3690 8570 3700
rect 9880 3690 9890 3700
rect 9930 3690 9940 3700
rect 0 3680 30 3690
rect 1610 3680 1690 3690
rect 2860 3680 2870 3690
rect 2910 3680 2920 3690
rect 3030 3680 3060 3690
rect 3320 3680 3330 3690
rect 3870 3680 3880 3690
rect 3940 3680 3960 3690
rect 4160 3680 4180 3690
rect 4880 3680 4940 3690
rect 5310 3680 5320 3690
rect 6070 3680 6470 3690
rect 8400 3680 8410 3690
rect 8450 3680 8460 3690
rect 8470 3680 8490 3690
rect 8560 3680 8570 3690
rect 9870 3680 9880 3690
rect 0 3670 40 3680
rect 1610 3670 1690 3680
rect 1700 3670 1710 3680
rect 3040 3670 3070 3680
rect 3290 3670 3310 3680
rect 3320 3670 3330 3680
rect 3870 3670 3880 3680
rect 3930 3670 3940 3680
rect 4090 3670 4130 3680
rect 4910 3670 4960 3680
rect 5310 3670 5320 3680
rect 6070 3670 6470 3680
rect 8400 3670 8410 3680
rect 8470 3670 8500 3680
rect 8590 3670 8600 3680
rect 9900 3670 9920 3680
rect 0 3660 50 3670
rect 1630 3660 1650 3670
rect 1660 3660 1670 3670
rect 1700 3660 1720 3670
rect 3070 3660 3090 3670
rect 3290 3660 3310 3670
rect 3330 3660 3340 3670
rect 3880 3660 3940 3670
rect 4930 3660 4990 3670
rect 6070 3660 6480 3670
rect 6980 3660 6990 3670
rect 8200 3660 8210 3670
rect 8460 3660 8470 3670
rect 8480 3660 8510 3670
rect 8580 3660 8590 3670
rect 9850 3660 9860 3670
rect 9880 3660 9890 3670
rect 1690 3650 1720 3660
rect 3090 3650 3130 3660
rect 3300 3650 3320 3660
rect 4960 3650 5010 3660
rect 6140 3650 6480 3660
rect 6970 3650 6980 3660
rect 8530 3650 8540 3660
rect 1670 3640 1690 3650
rect 1700 3640 1710 3650
rect 3070 3640 3120 3650
rect 3130 3640 3140 3650
rect 3300 3640 3320 3650
rect 3340 3640 3350 3650
rect 3950 3640 3960 3650
rect 4970 3640 5030 3650
rect 5320 3640 5330 3650
rect 6150 3640 6460 3650
rect 8400 3640 8410 3650
rect 8510 3640 8520 3650
rect 8530 3640 8550 3650
rect 9880 3640 9890 3650
rect 1640 3630 1650 3640
rect 1700 3630 1710 3640
rect 3150 3630 3160 3640
rect 3300 3630 3320 3640
rect 4990 3630 5020 3640
rect 5320 3630 5330 3640
rect 6160 3630 6460 3640
rect 8230 3630 8240 3640
rect 8380 3630 8390 3640
rect 8410 3630 8430 3640
rect 8500 3630 8510 3640
rect 9560 3630 9570 3640
rect 9870 3630 9880 3640
rect 1690 3620 1710 3630
rect 3170 3620 3180 3630
rect 3300 3620 3330 3630
rect 3350 3620 3360 3630
rect 5000 3620 5030 3630
rect 6170 3620 6460 3630
rect 6950 3620 6960 3630
rect 8370 3620 8390 3630
rect 8410 3620 8430 3630
rect 8490 3620 8520 3630
rect 9550 3620 9570 3630
rect 9850 3620 9860 3630
rect 9920 3620 9930 3630
rect 1680 3610 1690 3620
rect 1700 3610 1710 3620
rect 3170 3610 3190 3620
rect 3230 3610 3240 3620
rect 3300 3610 3350 3620
rect 6180 3610 6450 3620
rect 8380 3610 8390 3620
rect 8500 3610 8520 3620
rect 9540 3610 9560 3620
rect 9930 3610 9940 3620
rect 1490 3600 1500 3610
rect 1690 3600 1720 3610
rect 3210 3600 3220 3610
rect 3230 3600 3250 3610
rect 3310 3600 3350 3610
rect 6190 3600 6440 3610
rect 8260 3600 8270 3610
rect 8410 3600 8430 3610
rect 8500 3600 8510 3610
rect 9530 3600 9550 3610
rect 1480 3590 1490 3600
rect 1700 3590 1710 3600
rect 3230 3590 3250 3600
rect 3270 3590 3300 3600
rect 3320 3590 3340 3600
rect 3910 3590 3920 3600
rect 5330 3590 5340 3600
rect 6180 3590 6450 3600
rect 8380 3590 8390 3600
rect 8410 3590 8420 3600
rect 8430 3590 8440 3600
rect 8490 3590 8510 3600
rect 9500 3590 9540 3600
rect 1470 3580 1490 3590
rect 1690 3580 1720 3590
rect 3240 3580 3250 3590
rect 3280 3580 3300 3590
rect 3320 3580 3340 3590
rect 3360 3580 3370 3590
rect 4780 3580 4790 3590
rect 5330 3580 5340 3590
rect 6180 3580 6430 3590
rect 8400 3580 8420 3590
rect 8490 3580 8500 3590
rect 9490 3580 9530 3590
rect 1470 3570 1480 3580
rect 1690 3570 1710 3580
rect 3240 3570 3250 3580
rect 3280 3570 3290 3580
rect 3330 3570 3340 3580
rect 3370 3570 3380 3580
rect 3900 3570 3920 3580
rect 4770 3570 4800 3580
rect 5330 3570 5340 3580
rect 6180 3570 6400 3580
rect 6420 3570 6430 3580
rect 8390 3570 8400 3580
rect 8410 3570 8420 3580
rect 8430 3570 8440 3580
rect 8480 3570 8490 3580
rect 9470 3570 9530 3580
rect 1460 3560 1480 3570
rect 1680 3560 1710 3570
rect 3330 3560 3340 3570
rect 3900 3560 3920 3570
rect 4750 3560 4790 3570
rect 5330 3560 5340 3570
rect 6180 3560 6390 3570
rect 8390 3560 8400 3570
rect 8460 3560 8470 3570
rect 9440 3560 9510 3570
rect 1450 3550 1480 3560
rect 1690 3550 1700 3560
rect 3340 3550 3350 3560
rect 3380 3550 3390 3560
rect 3900 3550 3930 3560
rect 4740 3550 4750 3560
rect 4760 3550 4770 3560
rect 5330 3550 5340 3560
rect 6170 3550 6370 3560
rect 8320 3550 8330 3560
rect 8440 3550 8460 3560
rect 9430 3550 9500 3560
rect 1450 3540 1480 3550
rect 1690 3540 1700 3550
rect 3270 3540 3280 3550
rect 3900 3540 3930 3550
rect 4730 3540 4740 3550
rect 4750 3540 4760 3550
rect 6170 3540 6370 3550
rect 8330 3540 8340 3550
rect 8430 3540 8450 3550
rect 8480 3540 8490 3550
rect 9420 3540 9480 3550
rect 1440 3530 1480 3540
rect 1690 3530 1700 3540
rect 2710 3530 2720 3540
rect 3280 3530 3300 3540
rect 3390 3530 3400 3540
rect 3910 3530 3930 3540
rect 4720 3530 4750 3540
rect 6170 3530 6350 3540
rect 8400 3530 8410 3540
rect 8420 3530 8450 3540
rect 8480 3530 8490 3540
rect 9400 3530 9470 3540
rect 1430 3520 1480 3530
rect 1690 3520 1700 3530
rect 3280 3520 3310 3530
rect 3920 3520 3930 3530
rect 4710 3520 4740 3530
rect 5330 3520 5340 3530
rect 6160 3520 6350 3530
rect 6360 3520 6370 3530
rect 6870 3520 6880 3530
rect 8340 3520 8350 3530
rect 8430 3520 8440 3530
rect 8450 3520 8470 3530
rect 9390 3520 9450 3530
rect 1430 3510 1470 3520
rect 2570 3510 2580 3520
rect 3290 3510 3300 3520
rect 3310 3510 3320 3520
rect 3400 3510 3410 3520
rect 3920 3510 3930 3520
rect 4710 3510 4730 3520
rect 6160 3510 6370 3520
rect 8350 3510 8360 3520
rect 8430 3510 8470 3520
rect 8490 3510 8500 3520
rect 9360 3510 9430 3520
rect 1420 3500 1470 3510
rect 2500 3500 2540 3510
rect 2550 3500 2600 3510
rect 3920 3500 3940 3510
rect 5010 3500 5050 3510
rect 6160 3500 6350 3510
rect 8350 3500 8380 3510
rect 8440 3500 8450 3510
rect 8480 3500 8500 3510
rect 9290 3500 9410 3510
rect 1420 3490 1470 3500
rect 2440 3490 2480 3500
rect 2610 3490 2630 3500
rect 3310 3490 3330 3500
rect 3920 3490 3940 3500
rect 4990 3490 5010 3500
rect 5040 3490 5050 3500
rect 6160 3490 6340 3500
rect 8350 3490 8380 3500
rect 8440 3490 8460 3500
rect 9270 3490 9350 3500
rect 9360 3490 9380 3500
rect 1410 3480 1460 3490
rect 2390 3480 2400 3490
rect 2410 3480 2420 3490
rect 2690 3480 2750 3490
rect 3310 3480 3360 3490
rect 3920 3480 3940 3490
rect 4320 3480 4350 3490
rect 4670 3480 4680 3490
rect 4970 3480 4990 3490
rect 6160 3480 6330 3490
rect 6840 3480 6850 3490
rect 8360 3480 8380 3490
rect 8400 3480 8410 3490
rect 8470 3480 8480 3490
rect 9260 3480 9280 3490
rect 9340 3480 9360 3490
rect 9600 3480 9620 3490
rect 1410 3470 1460 3480
rect 2370 3470 2390 3480
rect 2400 3470 2410 3480
rect 2720 3470 2740 3480
rect 2760 3470 2810 3480
rect 3350 3470 3360 3480
rect 3380 3470 3390 3480
rect 3920 3470 3950 3480
rect 4320 3470 4350 3480
rect 4520 3470 4620 3480
rect 4630 3470 4690 3480
rect 4960 3470 4970 3480
rect 6150 3470 6320 3480
rect 6830 3470 6840 3480
rect 8480 3470 8490 3480
rect 9240 3470 9270 3480
rect 9310 3470 9320 3480
rect 9590 3470 9610 3480
rect 1400 3460 1450 3470
rect 2350 3460 2370 3470
rect 2810 3460 2820 3470
rect 3360 3460 3390 3470
rect 3430 3460 3440 3470
rect 3920 3460 3950 3470
rect 4300 3460 4350 3470
rect 4510 3460 4690 3470
rect 4940 3460 4950 3470
rect 6140 3460 6320 3470
rect 6820 3460 6830 3470
rect 8420 3460 8430 3470
rect 8480 3460 8490 3470
rect 8530 3460 8550 3470
rect 9220 3460 9260 3470
rect 9290 3460 9300 3470
rect 9570 3460 9600 3470
rect 1400 3450 1450 3460
rect 2300 3450 2310 3460
rect 2320 3450 2340 3460
rect 2850 3450 2870 3460
rect 3350 3450 3380 3460
rect 3390 3450 3400 3460
rect 3410 3450 3420 3460
rect 3430 3450 3440 3460
rect 3920 3450 3950 3460
rect 4310 3450 4350 3460
rect 4480 3450 4520 3460
rect 4590 3450 4690 3460
rect 4920 3450 4940 3460
rect 5870 3450 5880 3460
rect 6140 3450 6320 3460
rect 6810 3450 6820 3460
rect 8430 3450 8460 3460
rect 8520 3450 8530 3460
rect 8540 3450 8550 3460
rect 9210 3450 9240 3460
rect 9270 3450 9280 3460
rect 9550 3450 9600 3460
rect 1390 3440 1450 3450
rect 2280 3440 2290 3450
rect 2880 3440 2900 3450
rect 3380 3440 3390 3450
rect 3430 3440 3440 3450
rect 3930 3440 3960 3450
rect 4300 3440 4340 3450
rect 4460 3440 4480 3450
rect 4610 3440 4680 3450
rect 4900 3440 4930 3450
rect 5020 3440 5030 3450
rect 5330 3440 5340 3450
rect 5850 3440 5890 3450
rect 5900 3440 5910 3450
rect 5940 3440 5950 3450
rect 5960 3440 5970 3450
rect 6140 3440 6280 3450
rect 6300 3440 6320 3450
rect 6800 3440 6810 3450
rect 8450 3440 8470 3450
rect 8490 3440 8500 3450
rect 8520 3440 8530 3450
rect 8540 3440 8550 3450
rect 9200 3440 9220 3450
rect 9540 3440 9580 3450
rect 1390 3430 1450 3440
rect 2890 3430 2940 3440
rect 3930 3430 3960 3440
rect 4300 3430 4340 3440
rect 4410 3430 4460 3440
rect 4560 3430 4670 3440
rect 4900 3430 4910 3440
rect 5330 3430 5340 3440
rect 5850 3430 5990 3440
rect 6020 3430 6030 3440
rect 6130 3430 6270 3440
rect 6790 3430 6800 3440
rect 8450 3430 8480 3440
rect 8500 3430 8510 3440
rect 8540 3430 8550 3440
rect 9190 3430 9210 3440
rect 9530 3430 9580 3440
rect 1380 3420 1450 3430
rect 2240 3420 2250 3430
rect 2920 3420 2960 3430
rect 3410 3420 3420 3430
rect 3940 3420 3970 3430
rect 4300 3420 4330 3430
rect 4420 3420 4440 3430
rect 4510 3420 4660 3430
rect 4880 3420 4900 3430
rect 4970 3420 4990 3430
rect 5330 3420 5340 3430
rect 5860 3420 6020 3430
rect 6050 3420 6060 3430
rect 6130 3420 6240 3430
rect 6780 3420 6790 3430
rect 9170 3420 9190 3430
rect 9530 3420 9570 3430
rect 1380 3410 1440 3420
rect 2230 3410 2240 3420
rect 2960 3410 2970 3420
rect 3940 3410 3970 3420
rect 4290 3410 4330 3420
rect 4430 3410 4640 3420
rect 4700 3410 4710 3420
rect 4870 3410 4880 3420
rect 4940 3410 4950 3420
rect 5330 3410 5340 3420
rect 5840 3410 6020 3420
rect 6040 3410 6060 3420
rect 6130 3410 6230 3420
rect 8490 3410 8500 3420
rect 8530 3410 8540 3420
rect 9090 3410 9120 3420
rect 9160 3410 9180 3420
rect 9210 3410 9220 3420
rect 9530 3410 9560 3420
rect 1370 3400 1440 3410
rect 2210 3400 2230 3410
rect 2980 3400 2990 3410
rect 3950 3400 3980 3410
rect 4280 3400 4330 3410
rect 4450 3400 4610 3410
rect 4620 3400 4700 3410
rect 4850 3400 4860 3410
rect 4920 3400 4930 3410
rect 5000 3400 5010 3410
rect 5680 3400 5690 3410
rect 5860 3400 6060 3410
rect 6130 3400 6210 3410
rect 8500 3400 8510 3410
rect 9090 3400 9110 3410
rect 9520 3400 9550 3410
rect 1370 3390 1430 3400
rect 2190 3390 2220 3400
rect 2990 3390 3010 3400
rect 3950 3390 3980 3400
rect 4280 3390 4300 3400
rect 4310 3390 4330 3400
rect 4460 3390 4550 3400
rect 4620 3390 4630 3400
rect 4640 3390 4690 3400
rect 4750 3390 4770 3400
rect 4830 3390 4850 3400
rect 4910 3390 4920 3400
rect 5010 3390 5020 3400
rect 5680 3390 5710 3400
rect 5850 3390 6050 3400
rect 6140 3390 6200 3400
rect 8500 3390 8530 3400
rect 9100 3390 9110 3400
rect 9520 3390 9540 3400
rect 1360 3380 1430 3390
rect 2180 3380 2200 3390
rect 3020 3380 3040 3390
rect 3510 3380 3520 3390
rect 3960 3380 3980 3390
rect 4270 3380 4290 3390
rect 4300 3380 4320 3390
rect 4620 3380 4630 3390
rect 4750 3380 4780 3390
rect 4810 3380 4830 3390
rect 4900 3380 4910 3390
rect 5010 3380 5020 3390
rect 5680 3380 5730 3390
rect 5850 3380 6040 3390
rect 6140 3380 6200 3390
rect 8500 3380 8530 3390
rect 9110 3380 9120 3390
rect 9510 3380 9530 3390
rect 1360 3370 1420 3380
rect 2160 3370 2190 3380
rect 3030 3370 3040 3380
rect 3520 3370 3530 3380
rect 3960 3370 3990 3380
rect 4270 3370 4290 3380
rect 4300 3370 4330 3380
rect 4740 3370 4760 3380
rect 4770 3370 4800 3380
rect 5010 3370 5020 3380
rect 5630 3370 5650 3380
rect 5670 3370 5740 3380
rect 5830 3370 5840 3380
rect 5850 3370 6050 3380
rect 6140 3370 6170 3380
rect 6720 3370 6730 3380
rect 8500 3370 8520 3380
rect 9110 3370 9120 3380
rect 9500 3370 9520 3380
rect 9750 3370 9810 3380
rect 1360 3360 1420 3370
rect 2160 3360 2180 3370
rect 3050 3360 3060 3370
rect 3490 3360 3500 3370
rect 3970 3360 3990 3370
rect 4270 3360 4280 3370
rect 4300 3360 4320 3370
rect 4710 3360 4790 3370
rect 5320 3360 5330 3370
rect 5640 3360 5740 3370
rect 5850 3360 6050 3370
rect 6130 3360 6160 3370
rect 6710 3360 6720 3370
rect 8500 3360 8520 3370
rect 9110 3360 9120 3370
rect 9490 3360 9520 3370
rect 9730 3360 9740 3370
rect 1350 3350 1410 3360
rect 2160 3350 2170 3360
rect 3060 3350 3070 3360
rect 3480 3350 3510 3360
rect 3960 3350 4010 3360
rect 4260 3350 4280 3360
rect 4290 3350 4320 3360
rect 4690 3350 4780 3360
rect 5320 3350 5330 3360
rect 5640 3350 5760 3360
rect 5850 3350 6050 3360
rect 6130 3350 6160 3360
rect 8500 3350 8520 3360
rect 9490 3350 9510 3360
rect 1350 3340 1410 3350
rect 2140 3340 2150 3350
rect 3070 3340 3080 3350
rect 3480 3340 3490 3350
rect 3500 3340 3520 3350
rect 3570 3340 3580 3350
rect 3970 3340 4010 3350
rect 4260 3340 4270 3350
rect 4290 3340 4320 3350
rect 4660 3340 4760 3350
rect 4850 3340 4860 3350
rect 5630 3340 5760 3350
rect 5850 3340 6080 3350
rect 6130 3340 6160 3350
rect 6690 3340 6700 3350
rect 8490 3340 8500 3350
rect 9080 3340 9090 3350
rect 9480 3340 9500 3350
rect 9790 3340 9800 3350
rect 1340 3330 1410 3340
rect 2120 3330 2140 3340
rect 3090 3330 3100 3340
rect 3490 3330 3520 3340
rect 3980 3330 4010 3340
rect 4250 3330 4270 3340
rect 4280 3330 4320 3340
rect 4630 3330 4750 3340
rect 4790 3330 4820 3340
rect 4840 3330 4850 3340
rect 5000 3330 5010 3340
rect 5620 3330 5770 3340
rect 5850 3330 6060 3340
rect 6130 3330 6160 3340
rect 6670 3330 6680 3340
rect 9040 3330 9060 3340
rect 9130 3330 9140 3340
rect 9460 3330 9490 3340
rect 9720 3330 9760 3340
rect 1340 3320 1410 3330
rect 2120 3320 2130 3330
rect 3090 3320 3110 3330
rect 3510 3320 3530 3330
rect 3980 3320 4020 3330
rect 4240 3320 4270 3330
rect 4280 3320 4320 3330
rect 4610 3320 4740 3330
rect 4770 3320 4810 3330
rect 5000 3320 5010 3330
rect 5620 3320 5780 3330
rect 5840 3320 6080 3330
rect 6130 3320 6170 3330
rect 6660 3320 6680 3330
rect 9060 3320 9070 3330
rect 9450 3320 9480 3330
rect 9710 3320 9720 3330
rect 9730 3320 9760 3330
rect 1330 3310 1400 3320
rect 2110 3310 2120 3320
rect 3100 3310 3120 3320
rect 3500 3310 3510 3320
rect 3530 3310 3540 3320
rect 3990 3310 4030 3320
rect 4240 3310 4260 3320
rect 4280 3310 4320 3320
rect 4600 3310 4670 3320
rect 4690 3310 4720 3320
rect 4750 3310 4780 3320
rect 5000 3310 5010 3320
rect 5310 3310 5320 3320
rect 5620 3310 5780 3320
rect 5840 3310 6000 3320
rect 6010 3310 6090 3320
rect 6120 3310 6170 3320
rect 6670 3310 6680 3320
rect 9070 3310 9080 3320
rect 9440 3310 9470 3320
rect 9700 3310 9710 3320
rect 9740 3310 9770 3320
rect 1330 3300 1400 3310
rect 2100 3300 2110 3310
rect 3990 3300 4040 3310
rect 4240 3300 4320 3310
rect 4590 3300 4650 3310
rect 4740 3300 4760 3310
rect 4980 3300 5010 3310
rect 5620 3300 5790 3310
rect 5820 3300 6180 3310
rect 6660 3300 6680 3310
rect 9070 3300 9080 3310
rect 9110 3300 9120 3310
rect 9430 3300 9460 3310
rect 9670 3300 9710 3310
rect 9730 3300 9740 3310
rect 1320 3290 1400 3300
rect 2100 3290 2110 3300
rect 3120 3290 3130 3300
rect 3540 3290 3550 3300
rect 3570 3290 3580 3300
rect 4000 3290 4060 3300
rect 4230 3290 4310 3300
rect 4580 3290 4600 3300
rect 4980 3290 5000 3300
rect 5620 3290 5790 3300
rect 5800 3290 6170 3300
rect 8470 3290 8480 3300
rect 9060 3290 9070 3300
rect 9090 3290 9100 3300
rect 9420 3290 9450 3300
rect 9650 3290 9700 3300
rect 9710 3290 9740 3300
rect 1320 3280 1390 3290
rect 2090 3280 2100 3290
rect 3130 3280 3140 3290
rect 3560 3280 3600 3290
rect 4010 3280 4070 3290
rect 4230 3280 4310 3290
rect 4510 3280 4520 3290
rect 4550 3280 4580 3290
rect 4690 3280 4730 3290
rect 4970 3280 5000 3290
rect 5620 3280 6180 3290
rect 6660 3280 6670 3290
rect 9050 3280 9080 3290
rect 9400 3280 9440 3290
rect 9640 3280 9720 3290
rect 9990 3280 9990 3290
rect 1320 3270 1390 3280
rect 2080 3270 2100 3280
rect 3130 3270 3150 3280
rect 3570 3270 3590 3280
rect 4020 3270 4090 3280
rect 4230 3270 4310 3280
rect 4490 3270 4530 3280
rect 4690 3270 4700 3280
rect 4970 3270 4990 3280
rect 5300 3270 5310 3280
rect 5620 3270 6190 3280
rect 6570 3270 6600 3280
rect 6660 3270 6670 3280
rect 9050 3270 9060 3280
rect 9390 3270 9430 3280
rect 9630 3270 9680 3280
rect 9980 3270 9990 3280
rect 1310 3260 1390 3270
rect 2070 3260 2100 3270
rect 3140 3260 3150 3270
rect 3570 3260 3600 3270
rect 4030 3260 4110 3270
rect 4230 3260 4320 3270
rect 4450 3260 4470 3270
rect 4650 3260 4700 3270
rect 4730 3260 4750 3270
rect 4960 3260 4990 3270
rect 5630 3260 6190 3270
rect 6550 3260 6560 3270
rect 6650 3260 6670 3270
rect 9380 3260 9420 3270
rect 9620 3260 9650 3270
rect 9680 3260 9690 3270
rect 9970 3260 9980 3270
rect 1310 3250 1380 3260
rect 2070 3250 2090 3260
rect 3140 3250 3160 3260
rect 4030 3250 4110 3260
rect 4230 3250 4310 3260
rect 4430 3250 4440 3260
rect 4630 3250 4660 3260
rect 4740 3250 4750 3260
rect 4950 3250 4990 3260
rect 5630 3250 6200 3260
rect 6530 3250 6540 3260
rect 6650 3250 6660 3260
rect 9110 3250 9120 3260
rect 9370 3250 9390 3260
rect 9410 3250 9420 3260
rect 9600 3250 9640 3260
rect 9690 3250 9700 3260
rect 1300 3240 1380 3250
rect 2060 3240 2080 3250
rect 3140 3240 3170 3250
rect 4040 3240 4120 3250
rect 4230 3240 4260 3250
rect 4280 3240 4340 3250
rect 4400 3240 4420 3250
rect 4600 3240 4660 3250
rect 4740 3240 4750 3250
rect 4950 3240 4990 3250
rect 5640 3240 6200 3250
rect 6580 3240 6590 3250
rect 6650 3240 6660 3250
rect 9100 3240 9110 3250
rect 9370 3240 9380 3250
rect 9400 3240 9410 3250
rect 9590 3240 9630 3250
rect 9670 3240 9700 3250
rect 9950 3240 9960 3250
rect 1300 3230 1380 3240
rect 2060 3230 2070 3240
rect 4050 3230 4120 3240
rect 4240 3230 4260 3240
rect 4280 3230 4380 3240
rect 4620 3230 4650 3240
rect 4960 3230 4980 3240
rect 5290 3230 5300 3240
rect 5630 3230 6200 3240
rect 6580 3230 6590 3240
rect 6640 3230 6660 3240
rect 9090 3230 9100 3240
rect 9120 3230 9130 3240
rect 9360 3230 9370 3240
rect 9380 3230 9400 3240
rect 9570 3230 9610 3240
rect 9640 3230 9660 3240
rect 9950 3230 9980 3240
rect 1290 3220 1370 3230
rect 2060 3220 2070 3230
rect 3150 3220 3160 3230
rect 3560 3220 3570 3230
rect 3610 3220 3620 3230
rect 4050 3220 4140 3230
rect 4280 3220 4370 3230
rect 4630 3220 4650 3230
rect 4940 3220 4980 3230
rect 5650 3220 6210 3230
rect 6580 3220 6590 3230
rect 6650 3220 6660 3230
rect 9080 3220 9090 3230
rect 9130 3220 9140 3230
rect 9350 3220 9390 3230
rect 9560 3220 9600 3230
rect 9950 3220 9970 3230
rect 1290 3210 1370 3220
rect 2060 3210 2070 3220
rect 4070 3210 4150 3220
rect 4280 3210 4360 3220
rect 4580 3210 4600 3220
rect 4930 3210 4940 3220
rect 4950 3210 4960 3220
rect 4970 3210 4980 3220
rect 5650 3210 6210 3220
rect 6460 3210 6470 3220
rect 6580 3210 6590 3220
rect 6640 3210 6660 3220
rect 9140 3210 9150 3220
rect 9340 3210 9350 3220
rect 9360 3210 9380 3220
rect 9520 3210 9600 3220
rect 9960 3210 9970 3220
rect 1290 3200 1360 3210
rect 2050 3200 2070 3210
rect 3160 3200 3170 3210
rect 4060 3200 4150 3210
rect 4280 3200 4350 3210
rect 4520 3200 4540 3210
rect 4920 3200 4930 3210
rect 4960 3200 4970 3210
rect 5280 3200 5290 3210
rect 5670 3200 6210 3210
rect 6440 3200 6450 3210
rect 6580 3200 6590 3210
rect 6630 3200 6660 3210
rect 9070 3200 9080 3210
rect 9150 3200 9160 3210
rect 9360 3200 9370 3210
rect 9500 3200 9590 3210
rect 1280 3190 1360 3200
rect 2040 3190 2070 3200
rect 4070 3190 4160 3200
rect 4290 3190 4340 3200
rect 4490 3190 4510 3200
rect 5690 3190 6210 3200
rect 6410 3190 6420 3200
rect 6630 3190 6650 3200
rect 9170 3190 9200 3200
rect 9210 3190 9220 3200
rect 9250 3190 9260 3200
rect 9320 3190 9330 3200
rect 9360 3190 9370 3200
rect 9510 3190 9570 3200
rect 9580 3190 9590 3200
rect 9920 3190 9930 3200
rect 1280 3180 1360 3190
rect 2040 3180 2070 3190
rect 4060 3180 4110 3190
rect 4120 3180 4170 3190
rect 4300 3180 4350 3190
rect 4470 3180 4490 3190
rect 4900 3180 4910 3190
rect 5710 3180 6220 3190
rect 6380 3180 6390 3190
rect 6630 3180 6650 3190
rect 9040 3180 9060 3190
rect 9190 3180 9260 3190
rect 9310 3180 9330 3190
rect 9350 3180 9370 3190
rect 9490 3180 9590 3190
rect 9640 3180 9650 3190
rect 9900 3180 9910 3190
rect 1270 3170 1350 3180
rect 2030 3170 2060 3180
rect 4070 3170 4170 3180
rect 4300 3170 4380 3180
rect 4460 3170 4490 3180
rect 4900 3170 4920 3180
rect 5720 3170 6230 3180
rect 6630 3170 6650 3180
rect 9030 3170 9110 3180
rect 9220 3170 9370 3180
rect 9490 3170 9540 3180
rect 9620 3170 9640 3180
rect 9890 3170 9900 3180
rect 9940 3170 9950 3180
rect 1270 3160 1350 3170
rect 2030 3160 2060 3170
rect 4070 3160 4170 3170
rect 4460 3160 4480 3170
rect 4890 3160 4900 3170
rect 4930 3160 4940 3170
rect 5740 3160 5890 3170
rect 5900 3160 6240 3170
rect 6310 3160 6320 3170
rect 6570 3160 6580 3170
rect 6630 3160 6650 3170
rect 9020 3160 9060 3170
rect 9090 3160 9100 3170
rect 9250 3160 9320 3170
rect 9350 3160 9370 3170
rect 9480 3160 9530 3170
rect 9590 3160 9600 3170
rect 9620 3160 9630 3170
rect 9930 3160 9940 3170
rect 1270 3150 1350 3160
rect 2030 3150 2060 3160
rect 3750 3150 3760 3160
rect 4070 3150 4180 3160
rect 4410 3150 4420 3160
rect 4460 3150 4480 3160
rect 4870 3150 4900 3160
rect 4920 3150 4930 3160
rect 5770 3150 6250 3160
rect 6280 3150 6290 3160
rect 6570 3150 6580 3160
rect 6630 3150 6650 3160
rect 9000 3150 9040 3160
rect 9090 3150 9100 3160
rect 9260 3150 9300 3160
rect 9350 3150 9370 3160
rect 9470 3150 9530 3160
rect 9620 3150 9630 3160
rect 9920 3150 9930 3160
rect 1260 3140 1340 3150
rect 2030 3140 2050 3150
rect 3180 3140 3190 3150
rect 3720 3140 3730 3150
rect 3740 3140 3780 3150
rect 4070 3140 4190 3150
rect 4430 3140 4440 3150
rect 4460 3140 4480 3150
rect 4870 3140 4890 3150
rect 4910 3140 4920 3150
rect 5800 3140 6200 3150
rect 6210 3140 6220 3150
rect 6570 3140 6580 3150
rect 6620 3140 6640 3150
rect 8990 3140 9020 3150
rect 9090 3140 9100 3150
rect 9250 3140 9290 3150
rect 9350 3140 9360 3150
rect 9460 3140 9530 3150
rect 9610 3140 9620 3150
rect 9900 3140 9910 3150
rect 9920 3140 9930 3150
rect 1260 3130 1340 3140
rect 2030 3130 2040 3140
rect 3180 3130 3190 3140
rect 3720 3130 3740 3140
rect 3760 3130 3790 3140
rect 4080 3130 4200 3140
rect 4470 3130 4490 3140
rect 4850 3130 4880 3140
rect 4900 3130 4910 3140
rect 5850 3130 6170 3140
rect 6570 3130 6580 3140
rect 6620 3130 6640 3140
rect 8970 3130 8990 3140
rect 9090 3130 9100 3140
rect 9210 3130 9270 3140
rect 9350 3130 9360 3140
rect 9450 3130 9540 3140
rect 9870 3130 9880 3140
rect 1250 3120 1340 3130
rect 2030 3120 2040 3130
rect 3180 3120 3190 3130
rect 3720 3120 3730 3130
rect 3770 3120 3830 3130
rect 4080 3120 4160 3130
rect 4170 3120 4200 3130
rect 4460 3120 4470 3130
rect 4490 3120 4520 3130
rect 4840 3120 4860 3130
rect 4890 3120 4910 3130
rect 5910 3120 6060 3130
rect 6080 3120 6090 3130
rect 6100 3120 6110 3130
rect 6570 3120 6580 3130
rect 6610 3120 6640 3130
rect 8950 3120 8970 3130
rect 9080 3120 9100 3130
rect 9200 3120 9220 3130
rect 9440 3120 9450 3130
rect 9460 3120 9550 3130
rect 9850 3120 9860 3130
rect 9870 3120 9880 3130
rect 9930 3120 9940 3130
rect 1250 3110 1340 3120
rect 2020 3110 2040 3120
rect 3180 3110 3190 3120
rect 3770 3110 3830 3120
rect 3860 3110 3870 3120
rect 3880 3110 3890 3120
rect 4030 3110 4040 3120
rect 4090 3110 4120 3120
rect 4140 3110 4160 3120
rect 4170 3110 4210 3120
rect 4470 3110 4480 3120
rect 4500 3110 4540 3120
rect 4830 3110 4850 3120
rect 4880 3110 4910 3120
rect 5250 3110 5260 3120
rect 6570 3110 6580 3120
rect 6610 3110 6630 3120
rect 8380 3110 8390 3120
rect 8940 3110 8950 3120
rect 9070 3110 9100 3120
rect 9200 3110 9220 3120
rect 9340 3110 9350 3120
rect 9420 3110 9440 3120
rect 9460 3110 9540 3120
rect 9850 3110 9860 3120
rect 9940 3110 9950 3120
rect 1250 3100 1340 3110
rect 2020 3100 2040 3110
rect 3180 3100 3190 3110
rect 3790 3100 3830 3110
rect 3850 3100 3860 3110
rect 3890 3100 3900 3110
rect 4100 3100 4130 3110
rect 4150 3100 4170 3110
rect 4180 3100 4220 3110
rect 4480 3100 4490 3110
rect 4520 3100 4560 3110
rect 4810 3100 4840 3110
rect 4870 3100 4900 3110
rect 6560 3100 6580 3110
rect 6620 3100 6630 3110
rect 8920 3100 8930 3110
rect 9060 3100 9100 3110
rect 9200 3100 9220 3110
rect 9330 3100 9340 3110
rect 9400 3100 9440 3110
rect 9460 3100 9530 3110
rect 9870 3100 9880 3110
rect 9940 3100 9960 3110
rect 1240 3090 1330 3100
rect 2020 3090 2040 3100
rect 3180 3090 3190 3100
rect 3780 3090 3820 3100
rect 3850 3090 3860 3100
rect 3930 3090 3940 3100
rect 4040 3090 4050 3100
rect 4100 3090 4130 3100
rect 4160 3090 4190 3100
rect 4200 3090 4230 3100
rect 4550 3090 4590 3100
rect 4790 3090 4820 3100
rect 4870 3090 4890 3100
rect 5240 3090 5250 3100
rect 6560 3090 6570 3100
rect 6610 3090 6630 3100
rect 8430 3090 8440 3100
rect 9060 3090 9100 3100
rect 9200 3090 9230 3100
rect 9390 3090 9440 3100
rect 9460 3090 9520 3100
rect 9820 3090 9830 3100
rect 9870 3090 9890 3100
rect 9940 3090 9990 3100
rect 1240 3080 1330 3090
rect 2020 3080 2030 3090
rect 3180 3080 3200 3090
rect 3660 3080 3670 3090
rect 3780 3080 3870 3090
rect 4110 3080 4140 3090
rect 4170 3080 4240 3090
rect 4510 3080 4520 3090
rect 4570 3080 4620 3090
rect 4750 3080 4810 3090
rect 4850 3080 4880 3090
rect 6560 3080 6570 3090
rect 6610 3080 6630 3090
rect 9060 3080 9090 3090
rect 9210 3080 9240 3090
rect 9370 3080 9440 3090
rect 9460 3080 9510 3090
rect 9940 3080 9950 3090
rect 9960 3080 9990 3090
rect 1230 3070 1320 3080
rect 2010 3070 2030 3080
rect 3180 3070 3200 3080
rect 3780 3070 3880 3080
rect 4120 3070 4150 3080
rect 4180 3070 4200 3080
rect 4220 3070 4250 3080
rect 4520 3070 4530 3080
rect 4610 3070 4760 3080
rect 4830 3070 4880 3080
rect 6560 3070 6570 3080
rect 6610 3070 6630 3080
rect 8420 3070 8430 3080
rect 9050 3070 9080 3080
rect 9220 3070 9260 3080
rect 9360 3070 9450 3080
rect 9470 3070 9500 3080
rect 9970 3070 9990 3080
rect 1230 3060 1320 3070
rect 2010 3060 2020 3070
rect 3170 3060 3190 3070
rect 3760 3060 3770 3070
rect 3800 3060 3810 3070
rect 3830 3060 3880 3070
rect 4010 3060 4030 3070
rect 4060 3060 4070 3070
rect 4130 3060 4150 3070
rect 4190 3060 4220 3070
rect 4230 3060 4260 3070
rect 4540 3060 4550 3070
rect 4690 3060 4700 3070
rect 4710 3060 4720 3070
rect 4810 3060 4870 3070
rect 6560 3060 6570 3070
rect 6610 3060 6630 3070
rect 8390 3060 8400 3070
rect 8410 3060 8420 3070
rect 9050 3060 9090 3070
rect 9230 3060 9290 3070
rect 9330 3060 9460 3070
rect 9480 3060 9500 3070
rect 9790 3060 9800 3070
rect 9980 3060 9990 3070
rect 1230 3050 1320 3060
rect 2010 3050 2020 3060
rect 3170 3050 3190 3060
rect 3740 3050 3760 3060
rect 3830 3050 3870 3060
rect 4020 3050 4030 3060
rect 4140 3050 4160 3060
rect 4200 3050 4220 3060
rect 4240 3050 4280 3060
rect 4550 3050 4570 3060
rect 4800 3050 4860 3060
rect 6560 3050 6570 3060
rect 6600 3050 6620 3060
rect 8360 3050 8370 3060
rect 8390 3050 8410 3060
rect 9040 3050 9090 3060
rect 9250 3050 9500 3060
rect 9780 3050 9790 3060
rect 9890 3050 9900 3060
rect 1220 3040 1310 3050
rect 2010 3040 2020 3050
rect 3170 3040 3190 3050
rect 3740 3040 3750 3050
rect 3830 3040 3850 3050
rect 4040 3040 4050 3050
rect 4140 3040 4160 3050
rect 4210 3040 4290 3050
rect 4570 3040 4590 3050
rect 4780 3040 4850 3050
rect 5220 3040 5230 3050
rect 6550 3040 6570 3050
rect 6600 3040 6610 3050
rect 9040 3040 9080 3050
rect 9240 3040 9500 3050
rect 9770 3040 9780 3050
rect 9830 3040 9840 3050
rect 9890 3040 9900 3050
rect 1220 3030 1310 3040
rect 2010 3030 2020 3040
rect 3170 3030 3190 3040
rect 3740 3030 3750 3040
rect 4160 3030 4180 3040
rect 4220 3030 4300 3040
rect 4590 3030 4630 3040
rect 4750 3030 4820 3040
rect 6550 3030 6570 3040
rect 6590 3030 6610 3040
rect 9040 3030 9080 3040
rect 9230 3030 9490 3040
rect 9770 3030 9780 3040
rect 1210 3020 1310 3030
rect 2010 3020 2020 3030
rect 3170 3020 3200 3030
rect 3740 3020 3750 3030
rect 3760 3020 3770 3030
rect 3800 3020 3830 3030
rect 3840 3020 3850 3030
rect 3910 3020 3920 3030
rect 4090 3020 4100 3030
rect 4160 3020 4190 3030
rect 4230 3020 4310 3030
rect 4600 3020 4800 3030
rect 5210 3020 5220 3030
rect 6550 3020 6570 3030
rect 6590 3020 6620 3030
rect 8400 3020 8420 3030
rect 9040 3020 9080 3030
rect 9140 3020 9150 3030
rect 9220 3020 9430 3030
rect 9460 3020 9480 3030
rect 9900 3020 9910 3030
rect 1210 3010 1300 3020
rect 2010 3010 2020 3020
rect 3160 3010 3200 3020
rect 3730 3010 3780 3020
rect 3790 3010 3800 3020
rect 3820 3010 3830 3020
rect 3840 3010 3850 3020
rect 3860 3010 3870 3020
rect 3890 3010 3910 3020
rect 4100 3010 4110 3020
rect 4180 3010 4200 3020
rect 4240 3010 4320 3020
rect 4620 3010 4780 3020
rect 6550 3010 6560 3020
rect 6590 3010 6610 3020
rect 8430 3010 8440 3020
rect 9040 3010 9080 3020
rect 9130 3010 9170 3020
rect 9210 3010 9420 3020
rect 9790 3010 9800 3020
rect 9820 3010 9890 3020
rect 9900 3010 9910 3020
rect 1200 3000 1300 3010
rect 3160 3000 3200 3010
rect 3740 3000 3790 3010
rect 3810 3000 3850 3010
rect 3890 3000 3900 3010
rect 4050 3000 4070 3010
rect 4190 3000 4220 3010
rect 4240 3000 4330 3010
rect 4660 3000 4770 3010
rect 5200 3000 5210 3010
rect 6550 3000 6560 3010
rect 6590 3000 6610 3010
rect 8400 3000 8410 3010
rect 9030 3000 9080 3010
rect 9130 3000 9180 3010
rect 9200 3000 9420 3010
rect 9840 3000 9860 3010
rect 9890 3000 9900 3010
rect 1200 2990 1300 3000
rect 2010 2990 2020 3000
rect 3160 2990 3200 3000
rect 3770 2990 3780 3000
rect 3790 2990 3800 3000
rect 3820 2990 3840 3000
rect 3860 2990 3870 3000
rect 4200 2990 4330 3000
rect 4510 2990 4520 3000
rect 4620 2990 4630 3000
rect 4660 2990 4760 3000
rect 6550 2990 6560 3000
rect 6590 2990 6610 3000
rect 8440 2990 8450 3000
rect 9020 2990 9090 3000
rect 9120 2990 9180 3000
rect 9200 2990 9380 3000
rect 9400 2990 9410 3000
rect 1200 2980 1300 2990
rect 2000 2980 2010 2990
rect 3160 2980 3200 2990
rect 3860 2980 3880 2990
rect 4210 2980 4350 2990
rect 4510 2980 4520 2990
rect 4660 2980 4670 2990
rect 5190 2980 5200 2990
rect 6550 2980 6560 2990
rect 6580 2980 6610 2990
rect 8440 2980 8450 2990
rect 9000 2980 9080 2990
rect 9120 2980 9360 2990
rect 1190 2970 1290 2980
rect 2000 2970 2020 2980
rect 3160 2970 3200 2980
rect 3860 2970 3870 2980
rect 4040 2970 4050 2980
rect 4140 2970 4150 2980
rect 4230 2970 4350 2980
rect 4510 2970 4520 2980
rect 6550 2970 6560 2980
rect 6580 2970 6600 2980
rect 8440 2970 8450 2980
rect 8990 2970 9080 2980
rect 9110 2970 9150 2980
rect 9190 2970 9330 2980
rect 1190 2960 1290 2970
rect 2000 2960 2020 2970
rect 3160 2960 3190 2970
rect 3790 2960 3800 2970
rect 3880 2960 3890 2970
rect 4040 2960 4050 2970
rect 4150 2960 4160 2970
rect 4250 2960 4360 2970
rect 4510 2960 4520 2970
rect 4530 2960 4540 2970
rect 5180 2960 5190 2970
rect 6550 2960 6560 2970
rect 6580 2960 6600 2970
rect 8970 2960 9070 2970
rect 9110 2960 9130 2970
rect 9190 2960 9290 2970
rect 9300 2960 9320 2970
rect 1180 2950 1280 2960
rect 2000 2950 2010 2960
rect 3160 2950 3170 2960
rect 3780 2950 3810 2960
rect 3850 2950 3860 2960
rect 3990 2950 4000 2960
rect 4250 2950 4370 2960
rect 4530 2950 4560 2960
rect 6540 2950 6560 2960
rect 6580 2950 6600 2960
rect 8420 2950 8440 2960
rect 8960 2950 9070 2960
rect 9100 2950 9130 2960
rect 9190 2950 9280 2960
rect 9300 2950 9310 2960
rect 1180 2940 1280 2950
rect 2000 2940 2010 2950
rect 3160 2940 3170 2950
rect 3820 2940 3830 2950
rect 3860 2940 3880 2950
rect 3890 2940 3900 2950
rect 4270 2940 4380 2950
rect 4540 2940 4560 2950
rect 5170 2940 5180 2950
rect 6540 2940 6570 2950
rect 6580 2940 6600 2950
rect 8940 2940 9070 2950
rect 9100 2940 9120 2950
rect 9200 2940 9270 2950
rect 9710 2940 9730 2950
rect 1180 2930 1280 2940
rect 2000 2930 2010 2940
rect 3160 2930 3170 2940
rect 3850 2930 3880 2940
rect 4010 2930 4020 2940
rect 4040 2930 4050 2940
rect 4280 2930 4400 2940
rect 4550 2930 4560 2940
rect 5170 2930 5180 2940
rect 6540 2930 6560 2940
rect 6580 2930 6590 2940
rect 8930 2930 9060 2940
rect 9090 2930 9110 2940
rect 9210 2930 9270 2940
rect 9380 2930 9420 2940
rect 9700 2930 9710 2940
rect 9730 2930 9740 2940
rect 1170 2920 1270 2930
rect 2000 2920 2010 2930
rect 3810 2920 3830 2930
rect 3850 2920 3860 2930
rect 3930 2920 3950 2930
rect 4200 2920 4210 2930
rect 4290 2920 4410 2930
rect 5160 2920 5170 2930
rect 6540 2920 6550 2930
rect 6580 2920 6590 2930
rect 8980 2920 9060 2930
rect 9090 2920 9110 2930
rect 9210 2920 9250 2930
rect 9370 2920 9410 2930
rect 9710 2920 9720 2930
rect 1170 2910 1260 2920
rect 2000 2910 2010 2920
rect 3150 2910 3160 2920
rect 3810 2910 3850 2920
rect 3880 2910 3890 2920
rect 4210 2910 4220 2920
rect 4310 2910 4420 2920
rect 5160 2910 5170 2920
rect 6540 2910 6550 2920
rect 6570 2910 6590 2920
rect 8770 2910 8780 2920
rect 8960 2910 9060 2920
rect 9080 2910 9100 2920
rect 9220 2910 9250 2920
rect 9270 2910 9290 2920
rect 9370 2910 9410 2920
rect 1160 2900 1260 2910
rect 2000 2900 2010 2910
rect 3150 2900 3160 2910
rect 3780 2900 3790 2910
rect 3880 2900 3910 2910
rect 3920 2900 3950 2910
rect 4010 2900 4020 2910
rect 4330 2900 4430 2910
rect 5150 2900 5160 2910
rect 6540 2900 6560 2910
rect 6570 2900 6590 2910
rect 8270 2900 8280 2910
rect 8750 2900 8770 2910
rect 8940 2900 9060 2910
rect 9070 2900 9100 2910
rect 9220 2900 9250 2910
rect 9270 2900 9290 2910
rect 9370 2900 9410 2910
rect 1160 2890 1250 2900
rect 1990 2890 2010 2900
rect 3150 2890 3160 2900
rect 3890 2890 3900 2900
rect 3920 2890 3940 2900
rect 4350 2890 4440 2900
rect 5150 2890 5170 2900
rect 6540 2890 6590 2900
rect 8920 2890 8990 2900
rect 9000 2890 9090 2900
rect 9230 2890 9250 2900
rect 9360 2890 9400 2900
rect 1160 2880 1250 2890
rect 1990 2880 2000 2890
rect 3150 2880 3160 2890
rect 3590 2880 3600 2890
rect 3890 2880 3900 2890
rect 4360 2880 4450 2890
rect 5140 2880 5170 2890
rect 6540 2880 6580 2890
rect 8900 2880 8960 2890
rect 8990 2880 9080 2890
rect 9230 2880 9240 2890
rect 9370 2880 9390 2890
rect 9990 2880 9990 2890
rect 1150 2870 1250 2880
rect 1990 2870 2000 2880
rect 3150 2870 3160 2880
rect 3600 2870 3610 2880
rect 3850 2870 3870 2880
rect 3890 2870 3900 2880
rect 4250 2870 4260 2880
rect 4380 2870 4470 2880
rect 5140 2870 5170 2880
rect 6540 2870 6590 2880
rect 8880 2870 8940 2880
rect 8990 2870 9070 2880
rect 9990 2870 9990 2880
rect 1150 2860 1240 2870
rect 1990 2860 2000 2870
rect 3150 2860 3160 2870
rect 3860 2860 3900 2870
rect 3910 2860 3920 2870
rect 4400 2860 4480 2870
rect 5130 2860 5170 2870
rect 6530 2860 6580 2870
rect 8820 2860 8900 2870
rect 8990 2860 9060 2870
rect 9970 2860 9990 2870
rect 1140 2850 1230 2860
rect 1990 2850 2010 2860
rect 3150 2850 3160 2860
rect 3810 2850 3830 2860
rect 3860 2850 3880 2860
rect 3900 2850 3910 2860
rect 3930 2850 3940 2860
rect 4410 2850 4490 2860
rect 5120 2850 5170 2860
rect 6530 2850 6550 2860
rect 6560 2850 6570 2860
rect 8780 2850 8870 2860
rect 8980 2850 9050 2860
rect 9970 2850 9990 2860
rect 1140 2840 1230 2850
rect 1990 2840 2000 2850
rect 3150 2840 3160 2850
rect 3860 2840 3870 2850
rect 3900 2840 3940 2850
rect 4430 2840 4510 2850
rect 4630 2840 4660 2850
rect 5110 2840 5170 2850
rect 6530 2840 6570 2850
rect 8710 2840 8820 2850
rect 8960 2840 9040 2850
rect 1130 2830 1230 2840
rect 1990 2830 2000 2840
rect 3150 2830 3160 2840
rect 3890 2830 3900 2840
rect 3920 2830 3930 2840
rect 3980 2830 3990 2840
rect 4250 2830 4260 2840
rect 4450 2830 4530 2840
rect 4620 2830 4680 2840
rect 5090 2830 5170 2840
rect 6530 2830 6570 2840
rect 8670 2830 8790 2840
rect 8940 2830 9030 2840
rect 9360 2830 9370 2840
rect 9380 2830 9390 2840
rect 1130 2820 1230 2830
rect 1990 2820 2000 2830
rect 3150 2820 3160 2830
rect 3910 2820 3930 2830
rect 3960 2820 3970 2830
rect 3980 2820 3990 2830
rect 4460 2820 4550 2830
rect 4600 2820 4730 2830
rect 5080 2820 5170 2830
rect 6530 2820 6570 2830
rect 8210 2820 8220 2830
rect 8680 2820 8750 2830
rect 8920 2820 9020 2830
rect 9360 2820 9370 2830
rect 9640 2820 9650 2830
rect 9990 2820 9990 2830
rect 1120 2810 1220 2820
rect 1990 2810 2000 2820
rect 3150 2810 3160 2820
rect 4480 2810 4750 2820
rect 5070 2810 5170 2820
rect 5840 2810 5850 2820
rect 5870 2810 5880 2820
rect 5910 2810 6080 2820
rect 6530 2810 6570 2820
rect 8910 2810 9010 2820
rect 9420 2810 9430 2820
rect 9630 2810 9650 2820
rect 1120 2800 1210 2810
rect 1980 2800 2000 2810
rect 3130 2800 3150 2810
rect 3960 2800 3970 2810
rect 4490 2800 4770 2810
rect 5050 2800 5170 2810
rect 5790 2800 5820 2810
rect 5830 2800 6110 2810
rect 6520 2800 6570 2810
rect 8870 2800 9000 2810
rect 9580 2800 9590 2810
rect 9630 2800 9640 2810
rect 9920 2800 9930 2810
rect 1120 2790 1210 2800
rect 1980 2790 2000 2800
rect 3140 2790 3150 2800
rect 4260 2790 4270 2800
rect 4500 2790 4790 2800
rect 5020 2790 5070 2800
rect 5100 2790 5170 2800
rect 5740 2790 6120 2800
rect 6530 2790 6560 2800
rect 8840 2790 8990 2800
rect 9590 2790 9600 2800
rect 9630 2790 9650 2800
rect 9940 2790 9950 2800
rect 1110 2780 1210 2790
rect 1980 2780 2000 2790
rect 3130 2780 3150 2790
rect 3950 2780 3960 2790
rect 4520 2780 4790 2790
rect 4980 2780 5060 2790
rect 5100 2780 5180 2790
rect 5560 2780 5680 2790
rect 5700 2780 5760 2790
rect 5770 2780 6130 2790
rect 6520 2780 6560 2790
rect 8800 2780 8850 2790
rect 8870 2780 8980 2790
rect 9480 2780 9490 2790
rect 9640 2780 9660 2790
rect 9960 2780 9970 2790
rect 1110 2770 1200 2780
rect 3130 2770 3150 2780
rect 3860 2770 3870 2780
rect 3900 2770 3910 2780
rect 4540 2770 4810 2780
rect 4950 2770 5050 2780
rect 5100 2770 5170 2780
rect 5550 2770 6130 2780
rect 6520 2770 6550 2780
rect 8170 2770 8180 2780
rect 8750 2770 8780 2780
rect 8860 2770 8960 2780
rect 9450 2770 9460 2780
rect 9630 2770 9640 2780
rect 9670 2770 9680 2780
rect 1100 2760 1190 2770
rect 1980 2760 1990 2770
rect 3150 2760 3160 2770
rect 3860 2760 3880 2770
rect 3890 2760 3940 2770
rect 4160 2760 4180 2770
rect 4560 2760 4820 2770
rect 4940 2760 5030 2770
rect 5090 2760 5100 2770
rect 5120 2760 5180 2770
rect 5540 2760 6050 2770
rect 6120 2760 6130 2770
rect 6530 2760 6560 2770
rect 8730 2760 8750 2770
rect 8850 2760 8940 2770
rect 9680 2760 9690 2770
rect 9920 2760 9930 2770
rect 1100 2750 1190 2760
rect 1980 2750 2000 2760
rect 3150 2750 3160 2760
rect 3920 2750 3930 2760
rect 4190 2750 4200 2760
rect 4590 2750 4840 2760
rect 4860 2750 4880 2760
rect 4910 2750 5020 2760
rect 5090 2750 5100 2760
rect 5110 2750 5180 2760
rect 5530 2750 6040 2760
rect 6520 2750 6550 2760
rect 8710 2750 8740 2760
rect 8840 2750 8930 2760
rect 9400 2750 9410 2760
rect 9490 2750 9500 2760
rect 9530 2750 9540 2760
rect 9690 2750 9700 2760
rect 9910 2750 9920 2760
rect 1090 2740 1180 2750
rect 1980 2740 2010 2750
rect 3150 2740 3160 2750
rect 3920 2740 3930 2750
rect 4620 2740 5020 2750
rect 5100 2740 5180 2750
rect 5520 2740 5990 2750
rect 6520 2740 6550 2750
rect 7070 2740 7080 2750
rect 7630 2740 7640 2750
rect 8690 2740 8730 2750
rect 8800 2740 8930 2750
rect 9400 2740 9410 2750
rect 9520 2740 9530 2750
rect 9630 2740 9640 2750
rect 9710 2740 9720 2750
rect 9910 2740 9920 2750
rect 1090 2730 1180 2740
rect 1980 2730 2000 2740
rect 3150 2730 3160 2740
rect 3880 2730 3900 2740
rect 3910 2730 3920 2740
rect 4670 2730 5040 2740
rect 5120 2730 5180 2740
rect 5510 2730 5960 2740
rect 5970 2730 5990 2740
rect 6130 2730 6140 2740
rect 6520 2730 6550 2740
rect 8140 2730 8150 2740
rect 8680 2730 8740 2740
rect 8770 2730 8860 2740
rect 8890 2730 8930 2740
rect 9410 2730 9420 2740
rect 9540 2730 9550 2740
rect 9630 2730 9640 2740
rect 9690 2730 9700 2740
rect 9910 2730 9920 2740
rect 1080 2720 1170 2730
rect 1970 2720 2000 2730
rect 3150 2720 3160 2730
rect 3880 2720 3910 2730
rect 4690 2720 4700 2730
rect 4710 2720 5030 2730
rect 5120 2720 5190 2730
rect 5310 2720 5340 2730
rect 5500 2720 5950 2730
rect 6140 2720 6150 2730
rect 6520 2720 6550 2730
rect 8680 2720 8740 2730
rect 8750 2720 8940 2730
rect 9390 2720 9400 2730
rect 9560 2720 9570 2730
rect 9910 2720 9920 2730
rect 1080 2710 1150 2720
rect 1980 2710 2000 2720
rect 3150 2710 3160 2720
rect 3890 2710 3900 2720
rect 4730 2710 5010 2720
rect 5120 2710 5190 2720
rect 5240 2710 5370 2720
rect 5490 2710 5940 2720
rect 6150 2710 6160 2720
rect 6510 2710 6540 2720
rect 7650 2710 7660 2720
rect 8690 2710 8830 2720
rect 8900 2710 8940 2720
rect 9260 2710 9280 2720
rect 9370 2710 9380 2720
rect 9580 2710 9590 2720
rect 9620 2710 9630 2720
rect 9670 2710 9690 2720
rect 9920 2710 9940 2720
rect 1070 2700 1140 2710
rect 1980 2700 2000 2710
rect 3150 2700 3160 2710
rect 3890 2700 3910 2710
rect 4270 2700 4280 2710
rect 4770 2700 5010 2710
rect 5120 2700 5180 2710
rect 5220 2700 5380 2710
rect 5470 2700 5930 2710
rect 6510 2700 6540 2710
rect 8690 2700 8700 2710
rect 8710 2700 8740 2710
rect 8750 2700 8820 2710
rect 8930 2700 8940 2710
rect 9240 2700 9280 2710
rect 9600 2700 9610 2710
rect 9640 2700 9650 2710
rect 9940 2700 9980 2710
rect 1070 2690 1130 2700
rect 1980 2690 2000 2700
rect 3890 2690 3900 2700
rect 3910 2690 3920 2700
rect 4270 2690 4280 2700
rect 4860 2690 4990 2700
rect 5000 2690 5010 2700
rect 5120 2690 5170 2700
rect 5220 2690 5380 2700
rect 5460 2690 5890 2700
rect 6510 2690 6540 2700
rect 8760 2690 8810 2700
rect 8930 2690 9020 2700
rect 9220 2690 9270 2700
rect 9620 2690 9630 2700
rect 9660 2690 9670 2700
rect 9940 2690 9990 2700
rect 1070 2680 1130 2690
rect 1980 2680 1990 2690
rect 3890 2680 3900 2690
rect 4270 2680 4280 2690
rect 4840 2680 5000 2690
rect 5120 2680 5160 2690
rect 5210 2680 5380 2690
rect 5450 2680 5880 2690
rect 6510 2680 6540 2690
rect 6960 2680 6970 2690
rect 8780 2680 8800 2690
rect 8950 2680 9080 2690
rect 9170 2680 9260 2690
rect 9640 2680 9650 2690
rect 9680 2680 9690 2690
rect 9960 2680 9990 2690
rect 1060 2670 1120 2680
rect 3890 2670 3900 2680
rect 4220 2670 4230 2680
rect 4240 2670 4250 2680
rect 4840 2670 5000 2680
rect 5110 2670 5150 2680
rect 5190 2670 5370 2680
rect 5440 2670 5880 2680
rect 6190 2670 6200 2680
rect 6510 2670 6540 2680
rect 8980 2670 9250 2680
rect 9660 2670 9670 2680
rect 9700 2670 9710 2680
rect 9970 2670 9990 2680
rect 1060 2660 1110 2670
rect 1970 2660 1980 2670
rect 2260 2660 2330 2670
rect 2930 2660 2950 2670
rect 3020 2660 3050 2670
rect 3140 2660 3150 2670
rect 3890 2660 3910 2670
rect 4210 2660 4220 2670
rect 4830 2660 4900 2670
rect 4910 2660 4990 2670
rect 5090 2660 5100 2670
rect 5110 2660 5140 2670
rect 5180 2660 5370 2670
rect 5430 2660 5850 2670
rect 6200 2660 6210 2670
rect 6510 2660 6540 2670
rect 9000 2660 9240 2670
rect 9680 2660 9690 2670
rect 9720 2660 9730 2670
rect 9980 2660 9990 2670
rect 1050 2650 1100 2660
rect 1960 2650 1970 2660
rect 2200 2650 2220 2660
rect 2330 2650 2370 2660
rect 2890 2650 2910 2660
rect 3090 2650 3110 2660
rect 3120 2650 3130 2660
rect 3140 2650 3150 2660
rect 3890 2650 3900 2660
rect 4200 2650 4210 2660
rect 4820 2650 4870 2660
rect 4900 2650 4980 2660
rect 5090 2650 5120 2660
rect 5160 2650 5370 2660
rect 5420 2650 5820 2660
rect 5830 2650 5850 2660
rect 6210 2650 6220 2660
rect 6510 2650 6530 2660
rect 6920 2650 6930 2660
rect 8070 2650 8080 2660
rect 9010 2650 9230 2660
rect 9700 2650 9710 2660
rect 9740 2650 9750 2660
rect 9990 2650 9990 2660
rect 1050 2640 1100 2650
rect 1960 2640 1970 2650
rect 2160 2640 2170 2650
rect 2350 2640 2390 2650
rect 2870 2640 2880 2650
rect 2950 2640 2970 2650
rect 3050 2640 3060 2650
rect 3120 2640 3150 2650
rect 3890 2640 3900 2650
rect 4810 2640 4820 2650
rect 4830 2640 4840 2650
rect 4880 2640 4980 2650
rect 5070 2640 5100 2650
rect 5130 2640 5360 2650
rect 5410 2640 5830 2650
rect 6510 2640 6530 2650
rect 9020 2640 9080 2650
rect 9190 2640 9210 2650
rect 9720 2640 9730 2650
rect 9760 2640 9770 2650
rect 1040 2630 1090 2640
rect 1960 2630 1970 2640
rect 2140 2630 2150 2640
rect 2190 2630 2200 2640
rect 2370 2630 2390 2640
rect 2860 2630 2870 2640
rect 4730 2630 4740 2640
rect 4800 2630 4810 2640
rect 4860 2630 4950 2640
rect 5060 2630 5080 2640
rect 5110 2630 5360 2640
rect 5400 2630 5830 2640
rect 6230 2630 6240 2640
rect 6510 2630 6530 2640
rect 8050 2630 8060 2640
rect 9030 2630 9080 2640
rect 9180 2630 9200 2640
rect 9740 2630 9750 2640
rect 9780 2630 9790 2640
rect 1040 2620 1090 2630
rect 1950 2620 1960 2630
rect 2110 2620 2120 2630
rect 2160 2620 2180 2630
rect 2280 2620 2310 2630
rect 2380 2620 2400 2630
rect 2850 2620 2860 2630
rect 2950 2620 2960 2630
rect 3090 2620 3110 2630
rect 3230 2620 3240 2630
rect 3900 2620 3920 2630
rect 4830 2620 4950 2630
rect 5040 2620 5060 2630
rect 5090 2620 5350 2630
rect 5380 2620 5830 2630
rect 5850 2620 5860 2630
rect 6230 2620 6240 2630
rect 6510 2620 6520 2630
rect 9040 2620 9080 2630
rect 9170 2620 9190 2630
rect 9760 2620 9770 2630
rect 9800 2620 9810 2630
rect 9850 2620 9860 2630
rect 1030 2610 1090 2620
rect 2090 2610 2100 2620
rect 2130 2610 2140 2620
rect 2260 2610 2270 2620
rect 2290 2610 2340 2620
rect 2390 2610 2400 2620
rect 2840 2610 2860 2620
rect 2930 2610 2940 2620
rect 3090 2610 3120 2620
rect 3890 2610 3930 2620
rect 4800 2610 4950 2620
rect 4970 2610 5000 2620
rect 5010 2610 5040 2620
rect 5080 2610 5340 2620
rect 5360 2610 5820 2620
rect 5830 2610 5840 2620
rect 6240 2610 6250 2620
rect 6510 2610 6520 2620
rect 6880 2610 6890 2620
rect 8030 2610 8040 2620
rect 9050 2610 9080 2620
rect 9160 2610 9190 2620
rect 9780 2610 9790 2620
rect 9820 2610 9830 2620
rect 1030 2600 1080 2610
rect 1940 2600 1950 2610
rect 2120 2600 2130 2610
rect 2170 2600 2190 2610
rect 2320 2600 2360 2610
rect 2390 2600 2410 2610
rect 2830 2600 2860 2610
rect 3110 2600 3130 2610
rect 3250 2600 3260 2610
rect 3890 2600 3930 2610
rect 4260 2600 4270 2610
rect 4780 2600 5010 2610
rect 5050 2600 5810 2610
rect 5820 2600 5830 2610
rect 5900 2600 5910 2610
rect 6510 2600 6520 2610
rect 6870 2600 6880 2610
rect 9050 2600 9080 2610
rect 9160 2600 9190 2610
rect 9840 2600 9850 2610
rect 1020 2590 1080 2600
rect 1940 2590 1950 2600
rect 2060 2590 2070 2600
rect 2090 2590 2160 2600
rect 2390 2590 2410 2600
rect 2830 2590 2860 2600
rect 3130 2590 3160 2600
rect 3900 2590 3920 2600
rect 4740 2590 4970 2600
rect 5030 2590 5790 2600
rect 5830 2590 5840 2600
rect 5860 2590 5880 2600
rect 6250 2590 6260 2600
rect 6510 2590 6520 2600
rect 6860 2590 6870 2600
rect 9050 2590 9080 2600
rect 9160 2590 9170 2600
rect 9820 2590 9830 2600
rect 1020 2580 1060 2590
rect 2050 2580 2060 2590
rect 2080 2580 2090 2590
rect 2120 2580 2130 2590
rect 2390 2580 2410 2590
rect 2840 2580 2850 2590
rect 3900 2580 3920 2590
rect 3940 2580 3950 2590
rect 4220 2580 4230 2590
rect 4690 2580 4920 2590
rect 5010 2580 5800 2590
rect 5810 2580 5840 2590
rect 5880 2580 5890 2590
rect 6260 2580 6270 2590
rect 6510 2580 6520 2590
rect 8000 2580 8010 2590
rect 9010 2580 9020 2590
rect 9030 2580 9100 2590
rect 9110 2580 9160 2590
rect 1010 2570 1060 2580
rect 2040 2570 2050 2580
rect 2070 2570 2100 2580
rect 2110 2570 2120 2580
rect 2400 2570 2410 2580
rect 2970 2570 2980 2580
rect 3270 2570 3280 2580
rect 4050 2570 4060 2580
rect 4540 2570 4870 2580
rect 4990 2570 5780 2580
rect 5790 2570 5840 2580
rect 9020 2570 9150 2580
rect 9860 2570 9870 2580
rect 1010 2560 1060 2570
rect 2030 2560 2040 2570
rect 2330 2560 2350 2570
rect 2830 2560 2840 2570
rect 2900 2560 2910 2570
rect 3270 2560 3280 2570
rect 3910 2560 3930 2570
rect 4060 2560 4070 2570
rect 4200 2560 4220 2570
rect 4500 2560 4800 2570
rect 4950 2560 4960 2570
rect 4970 2560 4980 2570
rect 4990 2560 5770 2570
rect 5810 2560 5820 2570
rect 6270 2560 6280 2570
rect 9040 2560 9150 2570
rect 9480 2560 9490 2570
rect 9960 2560 9970 2570
rect 1000 2550 1060 2560
rect 2410 2550 2420 2560
rect 2880 2550 2890 2560
rect 3960 2550 3980 2560
rect 3990 2550 4000 2560
rect 4170 2550 4180 2560
rect 4500 2550 4690 2560
rect 4730 2550 4740 2560
rect 4920 2550 4930 2560
rect 4940 2550 5790 2560
rect 7150 2550 7160 2560
rect 7250 2550 7270 2560
rect 9050 2550 9160 2560
rect 9380 2550 9390 2560
rect 9410 2550 9420 2560
rect 9430 2550 9440 2560
rect 9560 2550 9570 2560
rect 9990 2550 9990 2560
rect 1000 2540 1060 2550
rect 2000 2540 2030 2550
rect 2370 2540 2390 2550
rect 2870 2540 2880 2550
rect 3920 2540 3930 2550
rect 4160 2540 4170 2550
rect 4230 2540 4240 2550
rect 4260 2540 4300 2550
rect 4510 2540 4600 2550
rect 4850 2540 4870 2550
rect 4880 2540 5770 2550
rect 6280 2540 6290 2550
rect 7160 2540 7170 2550
rect 7230 2540 7280 2550
rect 7770 2540 7780 2550
rect 9060 2540 9160 2550
rect 9420 2540 9430 2550
rect 9460 2540 9470 2550
rect 9500 2540 9520 2550
rect 990 2530 1040 2540
rect 1920 2530 1930 2540
rect 1990 2530 2020 2540
rect 2350 2530 2390 2540
rect 2830 2530 2840 2540
rect 2860 2530 2870 2540
rect 2880 2530 2890 2540
rect 2920 2530 2940 2540
rect 3140 2530 3150 2540
rect 3920 2530 3930 2540
rect 3950 2530 3960 2540
rect 4090 2530 4100 2540
rect 4840 2530 5770 2540
rect 6290 2530 6300 2540
rect 7250 2530 7280 2540
rect 7940 2530 7950 2540
rect 9060 2530 9150 2540
rect 9340 2530 9350 2540
rect 9370 2530 9390 2540
rect 9420 2530 9430 2540
rect 9560 2530 9580 2540
rect 9590 2530 9600 2540
rect 9980 2530 9990 2540
rect 990 2520 1040 2530
rect 1920 2520 1930 2530
rect 1990 2520 2010 2530
rect 2330 2520 2390 2530
rect 3180 2520 3190 2530
rect 3920 2520 3970 2530
rect 4100 2520 4110 2530
rect 4150 2520 4160 2530
rect 4720 2520 5770 2530
rect 7260 2520 7300 2530
rect 9060 2520 9150 2530
rect 9330 2520 9340 2530
rect 9420 2520 9430 2530
rect 9480 2520 9490 2530
rect 9510 2520 9520 2530
rect 9610 2520 9620 2530
rect 980 2510 1050 2520
rect 1920 2510 1930 2520
rect 1980 2510 2030 2520
rect 3920 2510 3940 2520
rect 3950 2510 3960 2520
rect 4110 2510 4120 2520
rect 4130 2510 4160 2520
rect 4670 2510 4690 2520
rect 4700 2510 5750 2520
rect 5760 2510 5770 2520
rect 6300 2510 6310 2520
rect 6790 2510 6800 2520
rect 7270 2510 7280 2520
rect 9050 2510 9150 2520
rect 9300 2510 9330 2520
rect 9470 2510 9480 2520
rect 9490 2510 9500 2520
rect 9610 2510 9620 2520
rect 9640 2510 9650 2520
rect 9970 2510 9980 2520
rect 980 2500 1040 2510
rect 1920 2500 1930 2510
rect 1970 2500 2000 2510
rect 3940 2500 3960 2510
rect 3970 2500 3980 2510
rect 4030 2500 4050 2510
rect 4090 2500 4100 2510
rect 4110 2500 4120 2510
rect 4150 2500 4160 2510
rect 4650 2500 4800 2510
rect 4830 2500 5770 2510
rect 7280 2500 7290 2510
rect 7310 2500 7320 2510
rect 9080 2500 9140 2510
rect 9470 2500 9480 2510
rect 9570 2500 9580 2510
rect 970 2490 1040 2500
rect 1910 2490 1930 2500
rect 3940 2490 3960 2500
rect 3990 2490 4010 2500
rect 4020 2490 4060 2500
rect 4090 2490 4130 2500
rect 4650 2490 5640 2500
rect 5660 2490 5760 2500
rect 6310 2490 6320 2500
rect 7290 2490 7300 2500
rect 9090 2490 9130 2500
rect 9560 2490 9580 2500
rect 970 2480 1040 2490
rect 1910 2480 1930 2490
rect 3980 2480 4010 2490
rect 4020 2480 4130 2490
rect 4600 2480 4610 2490
rect 4650 2480 5640 2490
rect 5660 2480 5760 2490
rect 6770 2480 6780 2490
rect 7290 2480 7300 2490
rect 9100 2480 9110 2490
rect 960 2470 1040 2480
rect 1910 2470 1920 2480
rect 3910 2470 3920 2480
rect 3940 2470 3950 2480
rect 3990 2470 4080 2480
rect 4100 2470 4110 2480
rect 4590 2470 4630 2480
rect 4650 2470 5610 2480
rect 5660 2470 5750 2480
rect 6320 2470 6330 2480
rect 7260 2470 7270 2480
rect 7300 2470 7310 2480
rect 7840 2470 7850 2480
rect 9450 2470 9460 2480
rect 960 2460 1030 2470
rect 3940 2460 3950 2470
rect 3980 2460 3990 2470
rect 4020 2460 4080 2470
rect 4590 2460 5590 2470
rect 5650 2460 5740 2470
rect 6760 2460 6770 2470
rect 7270 2460 7310 2470
rect 7340 2460 7350 2470
rect 9450 2460 9490 2470
rect 9730 2460 9740 2470
rect 950 2450 1030 2460
rect 1900 2450 1920 2460
rect 3910 2450 3920 2460
rect 3950 2450 3960 2460
rect 3980 2450 4010 2460
rect 4020 2450 4090 2460
rect 4580 2450 5560 2460
rect 5650 2450 5740 2460
rect 7280 2450 7290 2460
rect 7350 2450 7360 2460
rect 9290 2450 9300 2460
rect 9460 2450 9470 2460
rect 9490 2450 9500 2460
rect 9730 2450 9740 2460
rect 950 2440 1040 2450
rect 1900 2440 1910 2450
rect 3240 2440 3250 2450
rect 3950 2440 3960 2450
rect 3980 2440 4040 2450
rect 4060 2440 4080 2450
rect 4560 2440 4570 2450
rect 4600 2440 4610 2450
rect 4620 2440 5560 2450
rect 5610 2440 5630 2450
rect 5660 2440 5720 2450
rect 5730 2440 5750 2450
rect 6340 2440 6350 2450
rect 6750 2440 6760 2450
rect 9440 2440 9450 2450
rect 9470 2440 9480 2450
rect 9490 2440 9520 2450
rect 9750 2440 9760 2450
rect 940 2430 1040 2440
rect 1900 2430 1910 2440
rect 3920 2430 3930 2440
rect 3980 2430 4010 2440
rect 4030 2430 4040 2440
rect 4580 2430 4590 2440
rect 4610 2430 4890 2440
rect 4900 2430 5570 2440
rect 5650 2430 5710 2440
rect 7370 2430 7380 2440
rect 9260 2430 9270 2440
rect 9290 2430 9300 2440
rect 9430 2430 9440 2440
rect 9480 2430 9500 2440
rect 940 2420 1030 2430
rect 1900 2420 1910 2430
rect 3980 2420 4000 2430
rect 4010 2420 4040 2430
rect 4570 2420 4590 2430
rect 4600 2420 5550 2430
rect 5640 2420 5700 2430
rect 6350 2420 6360 2430
rect 7380 2420 7390 2430
rect 9230 2420 9240 2430
rect 9380 2420 9400 2430
rect 9470 2420 9490 2430
rect 9520 2420 9530 2430
rect 9790 2420 9800 2430
rect 930 2410 1030 2420
rect 1900 2410 1910 2420
rect 3260 2410 3270 2420
rect 4580 2410 4680 2420
rect 4690 2410 4820 2420
rect 4840 2410 5550 2420
rect 5560 2410 5570 2420
rect 5640 2410 5690 2420
rect 6740 2410 6750 2420
rect 7340 2410 7350 2420
rect 9250 2410 9260 2420
rect 9300 2410 9310 2420
rect 9430 2410 9440 2420
rect 9460 2410 9470 2420
rect 9480 2410 9490 2420
rect 9700 2410 9710 2420
rect 930 2400 1020 2410
rect 1900 2400 1910 2410
rect 3260 2400 3280 2410
rect 4530 2400 4560 2410
rect 4590 2400 4650 2410
rect 4660 2400 4670 2410
rect 4700 2400 4790 2410
rect 4800 2400 5560 2410
rect 5620 2400 5690 2410
rect 6360 2400 6370 2410
rect 7400 2400 7420 2410
rect 9290 2400 9300 2410
rect 9320 2400 9330 2410
rect 9580 2400 9590 2410
rect 920 2390 1020 2400
rect 1890 2390 1910 2400
rect 3250 2390 3290 2400
rect 4560 2390 4570 2400
rect 4600 2390 4680 2400
rect 4700 2390 4710 2400
rect 4720 2390 5570 2400
rect 5580 2390 5690 2400
rect 7410 2390 7430 2400
rect 9180 2390 9190 2400
rect 9280 2390 9290 2400
rect 9400 2390 9430 2400
rect 920 2380 1010 2390
rect 1890 2380 1900 2390
rect 3260 2380 3290 2390
rect 4590 2380 5690 2390
rect 6370 2380 6380 2390
rect 7390 2380 7400 2390
rect 8390 2380 8400 2390
rect 9310 2380 9320 2390
rect 9530 2380 9550 2390
rect 9580 2380 9590 2390
rect 9610 2380 9630 2390
rect 9690 2380 9700 2390
rect 9710 2380 9720 2390
rect 910 2370 1010 2380
rect 1880 2370 1900 2380
rect 3270 2370 3290 2380
rect 4540 2370 4710 2380
rect 4720 2370 5700 2380
rect 6730 2370 6740 2380
rect 9410 2370 9420 2380
rect 9540 2370 9570 2380
rect 9620 2370 9630 2380
rect 9680 2370 9690 2380
rect 9800 2370 9810 2380
rect 910 2360 1010 2370
rect 1880 2360 1890 2370
rect 3280 2360 3290 2370
rect 4480 2360 4580 2370
rect 4690 2360 5670 2370
rect 6380 2360 6390 2370
rect 6730 2360 6740 2370
rect 7420 2360 7430 2370
rect 7440 2360 7450 2370
rect 8400 2360 8410 2370
rect 9380 2360 9390 2370
rect 9400 2360 9410 2370
rect 9630 2360 9640 2370
rect 9670 2360 9680 2370
rect 9800 2360 9810 2370
rect 900 2350 1000 2360
rect 1880 2350 1890 2360
rect 3280 2350 3300 2360
rect 4590 2350 4600 2360
rect 4610 2350 4640 2360
rect 4650 2350 5660 2360
rect 6730 2350 6740 2360
rect 6840 2350 6850 2360
rect 6870 2350 6880 2360
rect 7440 2350 7460 2360
rect 8400 2350 8420 2360
rect 9150 2350 9160 2360
rect 9260 2350 9270 2360
rect 9350 2350 9360 2360
rect 9380 2350 9390 2360
rect 9460 2350 9480 2360
rect 9840 2350 9850 2360
rect 900 2340 1000 2350
rect 1880 2340 1890 2350
rect 3280 2340 3300 2350
rect 4500 2340 5670 2350
rect 6390 2340 6400 2350
rect 6730 2340 6740 2350
rect 6830 2340 6900 2350
rect 7450 2340 7460 2350
rect 7470 2340 7480 2350
rect 8420 2340 8430 2350
rect 9150 2340 9160 2350
rect 9260 2340 9270 2350
rect 9320 2340 9330 2350
rect 9340 2340 9360 2350
rect 9430 2340 9480 2350
rect 9620 2340 9640 2350
rect 9710 2340 9720 2350
rect 9830 2340 9850 2350
rect 890 2330 1000 2340
rect 1870 2330 1880 2340
rect 3290 2330 3310 2340
rect 4510 2330 4520 2340
rect 4530 2330 5650 2340
rect 6730 2330 6740 2340
rect 6830 2330 6910 2340
rect 7470 2330 7490 2340
rect 8440 2330 8460 2340
rect 8470 2330 8480 2340
rect 8490 2330 8500 2340
rect 9150 2330 9160 2340
rect 9210 2330 9220 2340
rect 9250 2330 9260 2340
rect 9270 2330 9280 2340
rect 9340 2330 9360 2340
rect 9400 2330 9410 2340
rect 9720 2330 9730 2340
rect 9810 2330 9840 2340
rect 880 2320 990 2330
rect 1870 2320 1880 2330
rect 3290 2320 3310 2330
rect 4510 2320 5480 2330
rect 5520 2320 5660 2330
rect 6840 2320 6930 2330
rect 8410 2320 8420 2330
rect 8490 2320 8520 2330
rect 9230 2320 9250 2330
rect 9360 2320 9370 2330
rect 9390 2320 9410 2330
rect 9440 2320 9450 2330
rect 9550 2320 9560 2330
rect 9710 2320 9730 2330
rect 9790 2320 9800 2330
rect 9810 2320 9830 2330
rect 880 2310 990 2320
rect 1870 2310 1880 2320
rect 3290 2310 3310 2320
rect 4500 2310 5660 2320
rect 6410 2310 6420 2320
rect 6730 2310 6740 2320
rect 6840 2310 6950 2320
rect 8520 2310 8540 2320
rect 9150 2310 9160 2320
rect 9380 2310 9390 2320
rect 9470 2310 9490 2320
rect 9820 2310 9830 2320
rect 870 2300 990 2310
rect 1870 2300 1880 2310
rect 3290 2300 3310 2310
rect 4470 2300 5480 2310
rect 5510 2300 5540 2310
rect 5560 2300 5660 2310
rect 6730 2300 6740 2310
rect 6830 2300 6950 2310
rect 7050 2300 7060 2310
rect 7490 2300 7500 2310
rect 7530 2300 7540 2310
rect 8540 2300 8560 2310
rect 9220 2300 9230 2310
rect 9370 2300 9380 2310
rect 9420 2300 9440 2310
rect 9620 2300 9640 2310
rect 870 2290 990 2300
rect 1860 2290 1880 2300
rect 3300 2290 3320 2300
rect 4440 2290 5480 2300
rect 5500 2290 5520 2300
rect 5530 2290 5640 2300
rect 6420 2290 6430 2300
rect 6730 2290 6740 2300
rect 6830 2290 6950 2300
rect 7040 2290 7070 2300
rect 7540 2290 7560 2300
rect 8550 2290 8560 2300
rect 9150 2290 9160 2300
rect 9210 2290 9220 2300
rect 9250 2290 9260 2300
rect 9610 2290 9620 2300
rect 9630 2290 9640 2300
rect 9720 2290 9730 2300
rect 860 2280 980 2290
rect 1860 2280 1870 2290
rect 3300 2280 3320 2290
rect 4070 2280 4180 2290
rect 4330 2280 5470 2290
rect 5480 2280 5520 2290
rect 5530 2280 5630 2290
rect 5920 2280 5940 2290
rect 6000 2280 6010 2290
rect 6730 2280 6740 2290
rect 6830 2280 6960 2290
rect 7040 2280 7100 2290
rect 7500 2280 7510 2290
rect 7560 2280 7570 2290
rect 8560 2280 8570 2290
rect 9190 2280 9210 2290
rect 9250 2280 9260 2290
rect 9580 2280 9590 2290
rect 9730 2280 9740 2290
rect 9790 2280 9800 2290
rect 860 2270 980 2280
rect 1860 2270 1870 2280
rect 3300 2270 3320 2280
rect 4070 2270 4150 2280
rect 4210 2270 4220 2280
rect 4230 2270 4240 2280
rect 4250 2270 5430 2280
rect 5440 2270 5460 2280
rect 5490 2270 5510 2280
rect 5530 2270 5650 2280
rect 6000 2270 6010 2280
rect 6430 2270 6440 2280
rect 6730 2270 6740 2280
rect 6820 2270 6970 2280
rect 7050 2270 7170 2280
rect 7570 2270 7580 2280
rect 8570 2270 8580 2280
rect 9180 2270 9190 2280
rect 9260 2270 9270 2280
rect 9500 2270 9510 2280
rect 850 2260 980 2270
rect 1850 2260 1870 2270
rect 3300 2260 3320 2270
rect 4130 2260 5410 2270
rect 5480 2260 5510 2270
rect 5520 2260 5530 2270
rect 5540 2260 5640 2270
rect 6730 2260 6740 2270
rect 6820 2260 6890 2270
rect 6900 2260 6990 2270
rect 7070 2260 7090 2270
rect 7120 2260 7200 2270
rect 7510 2260 7520 2270
rect 7580 2260 7590 2270
rect 8580 2260 8590 2270
rect 9340 2260 9350 2270
rect 9360 2260 9370 2270
rect 9520 2260 9530 2270
rect 9790 2260 9800 2270
rect 850 2250 980 2260
rect 1850 2250 1860 2260
rect 3300 2250 3320 2260
rect 4260 2250 4270 2260
rect 4290 2250 4310 2260
rect 4330 2250 5420 2260
rect 5530 2250 5540 2260
rect 5550 2250 5640 2260
rect 6820 2250 6900 2260
rect 6910 2250 6920 2260
rect 6940 2250 7000 2260
rect 7040 2250 7050 2260
rect 7080 2250 7110 2260
rect 7150 2250 7170 2260
rect 7180 2250 7240 2260
rect 7250 2250 7260 2260
rect 7590 2250 7600 2260
rect 8600 2250 8610 2260
rect 9130 2250 9140 2260
rect 9590 2250 9600 2260
rect 840 2240 980 2250
rect 1850 2240 1860 2250
rect 3300 2240 3330 2250
rect 4340 2240 5420 2250
rect 5430 2240 5440 2250
rect 5540 2240 5590 2250
rect 6830 2240 6940 2250
rect 6950 2240 7020 2250
rect 7040 2240 7130 2250
rect 7220 2240 7270 2250
rect 7600 2240 7610 2250
rect 8630 2240 8640 2250
rect 9100 2240 9110 2250
rect 9590 2240 9600 2250
rect 840 2230 980 2240
rect 1850 2230 1860 2240
rect 3310 2230 3330 2240
rect 4350 2230 5410 2240
rect 5540 2230 5600 2240
rect 6450 2230 6460 2240
rect 6860 2230 6930 2240
rect 6980 2230 6990 2240
rect 7000 2230 7140 2240
rect 7240 2230 7280 2240
rect 7610 2230 7620 2240
rect 8730 2230 8740 2240
rect 8760 2230 8780 2240
rect 9070 2230 9090 2240
rect 9580 2230 9590 2240
rect 830 2220 980 2230
rect 1850 2220 1860 2230
rect 3310 2220 3340 2230
rect 4360 2220 5400 2230
rect 5460 2220 5470 2230
rect 5500 2220 5520 2230
rect 5530 2220 5570 2230
rect 5580 2220 5590 2230
rect 6880 2220 6960 2230
rect 7040 2220 7090 2230
rect 7100 2220 7140 2230
rect 7260 2220 7300 2230
rect 7360 2220 7370 2230
rect 7520 2220 7530 2230
rect 7620 2220 7640 2230
rect 8690 2220 8710 2230
rect 9050 2220 9060 2230
rect 9550 2220 9560 2230
rect 9810 2220 9820 2230
rect 830 2210 980 2220
rect 1850 2210 1860 2220
rect 3300 2210 3340 2220
rect 4340 2210 5390 2220
rect 5470 2210 5490 2220
rect 5510 2210 5520 2220
rect 5530 2210 5580 2220
rect 5600 2210 5610 2220
rect 6460 2210 6470 2220
rect 6900 2210 6970 2220
rect 7290 2210 7330 2220
rect 7340 2210 7380 2220
rect 7520 2210 7530 2220
rect 7630 2210 7650 2220
rect 8830 2210 8840 2220
rect 9000 2210 9010 2220
rect 9330 2210 9340 2220
rect 9560 2210 9570 2220
rect 820 2200 980 2210
rect 1850 2200 1860 2210
rect 3300 2200 3340 2210
rect 4350 2200 5370 2210
rect 5470 2200 5500 2210
rect 5510 2200 5530 2210
rect 5580 2200 5590 2210
rect 6740 2200 6750 2210
rect 6910 2200 6990 2210
rect 7300 2200 7380 2210
rect 7520 2200 7530 2210
rect 7640 2200 7660 2210
rect 8850 2200 8860 2210
rect 8920 2200 8940 2210
rect 9580 2200 9590 2210
rect 9670 2200 9680 2210
rect 9710 2200 9720 2210
rect 9980 2200 9990 2210
rect 820 2190 980 2200
rect 1850 2190 1860 2200
rect 2710 2190 2720 2200
rect 3310 2190 3340 2200
rect 4360 2190 5360 2200
rect 5470 2190 5490 2200
rect 5510 2190 5520 2200
rect 5530 2190 5550 2200
rect 6740 2190 6750 2200
rect 6920 2190 7010 2200
rect 7320 2190 7380 2200
rect 7510 2190 7530 2200
rect 7650 2190 7680 2200
rect 9370 2190 9380 2200
rect 9720 2190 9730 2200
rect 9960 2190 9990 2200
rect 810 2180 980 2190
rect 1840 2180 1860 2190
rect 2670 2180 2680 2190
rect 2750 2180 2760 2190
rect 3300 2180 3340 2190
rect 4350 2180 5330 2190
rect 5470 2180 5490 2190
rect 5520 2180 5540 2190
rect 6470 2180 6480 2190
rect 6740 2180 6750 2190
rect 6940 2180 7030 2190
rect 7330 2180 7350 2190
rect 7380 2180 7390 2190
rect 7510 2180 7520 2190
rect 7650 2180 7680 2190
rect 9390 2180 9400 2190
rect 9720 2180 9730 2190
rect 9960 2180 9970 2190
rect 800 2170 980 2180
rect 1840 2170 1850 2180
rect 2440 2170 2450 2180
rect 2750 2170 2760 2180
rect 3300 2170 3330 2180
rect 4360 2170 5320 2180
rect 5480 2170 5510 2180
rect 6960 2170 7050 2180
rect 7380 2170 7390 2180
rect 7510 2170 7520 2180
rect 7670 2170 7690 2180
rect 9240 2170 9250 2180
rect 9410 2170 9420 2180
rect 800 2160 980 2170
rect 1840 2160 1850 2170
rect 2430 2160 2440 2170
rect 2640 2160 2650 2170
rect 2740 2160 2750 2170
rect 3300 2160 3330 2170
rect 4360 2160 5150 2170
rect 5160 2160 5310 2170
rect 6970 2160 7060 2170
rect 7310 2160 7320 2170
rect 7380 2160 7390 2170
rect 7500 2160 7510 2170
rect 7670 2160 7710 2170
rect 9240 2160 9250 2170
rect 9560 2160 9570 2170
rect 790 2150 980 2160
rect 1840 2150 1850 2160
rect 2420 2150 2440 2160
rect 2630 2150 2640 2160
rect 2730 2150 2740 2160
rect 3300 2150 3330 2160
rect 4360 2150 5310 2160
rect 6950 2150 7080 2160
rect 7290 2150 7300 2160
rect 7420 2150 7440 2160
rect 7480 2150 7520 2160
rect 7670 2150 7730 2160
rect 9450 2150 9460 2160
rect 790 2140 970 2150
rect 1840 2140 1850 2150
rect 2430 2140 2450 2150
rect 2630 2140 2640 2150
rect 2710 2140 2730 2150
rect 3300 2140 3340 2150
rect 4360 2140 5170 2150
rect 5180 2140 5290 2150
rect 6750 2140 6760 2150
rect 6970 2140 6990 2150
rect 7000 2140 7090 2150
rect 7250 2140 7290 2150
rect 7420 2140 7440 2150
rect 7460 2140 7510 2150
rect 7670 2140 7680 2150
rect 7700 2140 7740 2150
rect 780 2130 970 2140
rect 2450 2130 2460 2140
rect 2530 2130 2540 2140
rect 2640 2130 2660 2140
rect 3300 2130 3340 2140
rect 4360 2130 5170 2140
rect 5180 2130 5280 2140
rect 6500 2130 6510 2140
rect 6750 2130 6760 2140
rect 6990 2130 7070 2140
rect 7240 2130 7290 2140
rect 7420 2130 7510 2140
rect 7710 2130 7800 2140
rect 7820 2130 7850 2140
rect 780 2120 970 2130
rect 1840 2120 1850 2130
rect 3300 2120 3340 2130
rect 4370 2120 5270 2130
rect 5400 2120 5410 2130
rect 6750 2120 6760 2130
rect 7000 2120 7090 2130
rect 7220 2120 7290 2130
rect 7430 2120 7490 2130
rect 7730 2120 7850 2130
rect 770 2110 970 2120
rect 3300 2110 3340 2120
rect 4360 2110 5300 2120
rect 7020 2110 7290 2120
rect 7420 2110 7480 2120
rect 7750 2110 7850 2120
rect 8390 2110 8400 2120
rect 9740 2110 9760 2120
rect 770 2100 970 2110
rect 1840 2100 1850 2110
rect 3300 2100 3340 2110
rect 4350 2100 5250 2110
rect 5260 2100 5290 2110
rect 6140 2100 6150 2110
rect 7030 2100 7280 2110
rect 7830 2100 7850 2110
rect 8400 2100 8410 2110
rect 760 2090 960 2100
rect 1840 2090 1850 2100
rect 3300 2090 3340 2100
rect 4340 2090 5290 2100
rect 6520 2090 6530 2100
rect 6760 2090 6770 2100
rect 7040 2090 7240 2100
rect 7250 2090 7270 2100
rect 7830 2090 7870 2100
rect 8410 2090 8420 2100
rect 9540 2090 9560 2100
rect 760 2080 950 2090
rect 1840 2080 1850 2090
rect 3300 2080 3340 2090
rect 4340 2080 5190 2090
rect 5200 2080 5280 2090
rect 6520 2080 6530 2090
rect 6760 2080 6770 2090
rect 7060 2080 7260 2090
rect 7830 2080 7870 2090
rect 8420 2080 8430 2090
rect 9230 2080 9240 2090
rect 9260 2080 9270 2090
rect 9330 2080 9340 2090
rect 9470 2080 9480 2090
rect 750 2070 950 2080
rect 1840 2070 1850 2080
rect 3290 2070 3340 2080
rect 4350 2070 5260 2080
rect 6150 2070 6160 2080
rect 6510 2070 6530 2080
rect 6760 2070 6770 2080
rect 7050 2070 7180 2080
rect 7210 2070 7250 2080
rect 7830 2070 7870 2080
rect 8430 2070 8460 2080
rect 9220 2070 9230 2080
rect 9270 2070 9280 2080
rect 9380 2070 9400 2080
rect 9670 2070 9680 2080
rect 750 2060 950 2070
rect 1840 2060 1850 2070
rect 3300 2060 3350 2070
rect 4350 2060 5110 2070
rect 5130 2060 5160 2070
rect 5170 2060 5260 2070
rect 6510 2060 6540 2070
rect 6760 2060 6770 2070
rect 7070 2060 7220 2070
rect 7320 2060 7330 2070
rect 7730 2060 7760 2070
rect 7830 2060 7880 2070
rect 8440 2060 8480 2070
rect 9180 2060 9200 2070
rect 9310 2060 9320 2070
rect 9560 2060 9570 2070
rect 9580 2060 9590 2070
rect 9640 2060 9670 2070
rect 740 2050 950 2060
rect 3290 2050 3350 2060
rect 4370 2050 5060 2060
rect 5070 2050 5080 2060
rect 5120 2050 5130 2060
rect 5140 2050 5150 2060
rect 5160 2050 5240 2060
rect 5250 2050 5260 2060
rect 6510 2050 6540 2060
rect 6770 2050 6780 2060
rect 7100 2050 7130 2060
rect 7150 2050 7170 2060
rect 7210 2050 7250 2060
rect 7730 2050 7740 2060
rect 7750 2050 7760 2060
rect 7830 2050 7880 2060
rect 8470 2050 8480 2060
rect 8500 2050 8510 2060
rect 9240 2050 9250 2060
rect 9490 2050 9510 2060
rect 9630 2050 9660 2060
rect 740 2040 950 2050
rect 3300 2040 3350 2050
rect 4370 2040 5110 2050
rect 5150 2040 5240 2050
rect 6510 2040 6540 2050
rect 7160 2040 7180 2050
rect 7220 2040 7230 2050
rect 7730 2040 7780 2050
rect 7850 2040 7890 2050
rect 8520 2040 8530 2050
rect 9160 2040 9170 2050
rect 730 2030 960 2040
rect 1840 2030 1850 2040
rect 3300 2030 3350 2040
rect 4370 2030 5120 2040
rect 5150 2030 5230 2040
rect 5260 2030 5270 2040
rect 6520 2030 6540 2040
rect 6770 2030 6780 2040
rect 7730 2030 7790 2040
rect 7850 2030 7910 2040
rect 7930 2030 7960 2040
rect 7980 2030 8000 2040
rect 8530 2030 8550 2040
rect 9110 2030 9120 2040
rect 9320 2030 9390 2040
rect 9460 2030 9470 2040
rect 730 2020 950 2030
rect 1840 2020 1850 2030
rect 3300 2020 3350 2030
rect 4350 2020 4360 2030
rect 4370 2020 5130 2030
rect 5140 2020 5150 2030
rect 5170 2020 5230 2030
rect 5250 2020 5260 2030
rect 6520 2020 6540 2030
rect 6770 2020 6780 2030
rect 7740 2020 7790 2030
rect 7860 2020 7870 2030
rect 7890 2020 8000 2030
rect 8530 2020 8570 2030
rect 9220 2020 9320 2030
rect 9390 2020 9400 2030
rect 9410 2020 9420 2030
rect 9460 2020 9470 2030
rect 720 2010 940 2020
rect 1840 2010 1850 2020
rect 3310 2010 3350 2020
rect 4370 2010 5150 2020
rect 5210 2010 5230 2020
rect 6520 2010 6540 2020
rect 6770 2010 6780 2020
rect 7760 2010 7790 2020
rect 7850 2010 7860 2020
rect 7940 2010 7990 2020
rect 8550 2010 8600 2020
rect 9150 2010 9180 2020
rect 720 2000 930 2010
rect 1840 2000 1850 2010
rect 3310 2000 3350 2010
rect 4340 2000 4350 2010
rect 4360 2000 5160 2010
rect 5210 2000 5220 2010
rect 6520 2000 6540 2010
rect 6770 2000 6780 2010
rect 7850 2000 7890 2010
rect 7950 2000 7970 2010
rect 8570 2000 8620 2010
rect 710 1990 930 2000
rect 1840 1990 1850 2000
rect 3310 1990 3350 2000
rect 4340 1990 5010 2000
rect 5030 1990 5140 2000
rect 5150 1990 5160 2000
rect 6160 1990 6180 2000
rect 6200 1990 6210 2000
rect 6230 1990 6240 2000
rect 6520 1990 6540 2000
rect 6770 1990 6790 2000
rect 7720 1990 7760 2000
rect 7820 1990 7830 2000
rect 7860 1990 7970 2000
rect 8590 1990 8680 2000
rect 9060 1990 9070 2000
rect 710 1980 930 1990
rect 3310 1980 3350 1990
rect 4330 1980 4820 1990
rect 4840 1980 5060 1990
rect 5140 1980 5150 1990
rect 6160 1980 6180 1990
rect 6190 1980 6240 1990
rect 6520 1980 6550 1990
rect 6770 1980 6790 1990
rect 7720 1980 7780 1990
rect 7840 1980 7850 1990
rect 7870 1980 7980 1990
rect 8610 1980 8710 1990
rect 700 1970 930 1980
rect 1840 1970 1850 1980
rect 3320 1970 3350 1980
rect 4350 1970 4830 1980
rect 4840 1970 4850 1980
rect 4870 1970 4910 1980
rect 4920 1970 4930 1980
rect 4940 1970 5030 1980
rect 6140 1970 6150 1980
rect 6220 1970 6230 1980
rect 6530 1970 6550 1980
rect 6780 1970 6790 1980
rect 7720 1970 7770 1980
rect 7850 1970 7860 1980
rect 7880 1970 7980 1980
rect 8680 1970 8730 1980
rect 700 1960 940 1970
rect 3320 1960 3350 1970
rect 4360 1960 4860 1970
rect 4880 1960 4910 1970
rect 4920 1960 4990 1970
rect 5000 1960 5030 1970
rect 6190 1960 6200 1970
rect 6210 1960 6270 1970
rect 6530 1960 6550 1970
rect 6780 1960 6790 1970
rect 7730 1960 7770 1970
rect 7860 1960 7870 1970
rect 7890 1960 7970 1970
rect 8710 1960 8720 1970
rect 8730 1960 8770 1970
rect 8810 1960 8860 1970
rect 8880 1960 8950 1970
rect 9010 1960 9020 1970
rect 690 1950 940 1960
rect 1840 1950 1850 1960
rect 3320 1950 3350 1960
rect 4360 1950 5030 1960
rect 6170 1950 6190 1960
rect 6200 1950 6310 1960
rect 6540 1950 6550 1960
rect 6780 1950 6800 1960
rect 7730 1950 7780 1960
rect 7950 1950 7960 1960
rect 8760 1950 8810 1960
rect 9880 1950 9890 1960
rect 9900 1950 9910 1960
rect 9920 1950 9960 1960
rect 690 1940 930 1950
rect 1840 1940 1850 1950
rect 3320 1940 3350 1950
rect 4360 1940 5020 1950
rect 6170 1940 6310 1950
rect 6520 1940 6530 1950
rect 6540 1940 6560 1950
rect 6780 1940 6790 1950
rect 7330 1940 7340 1950
rect 7730 1940 7780 1950
rect 7900 1940 7940 1950
rect 680 1930 930 1940
rect 1840 1930 1850 1940
rect 3320 1930 3350 1940
rect 4380 1930 4540 1940
rect 4620 1930 4780 1940
rect 4860 1930 4980 1940
rect 6170 1930 6340 1940
rect 6520 1930 6560 1940
rect 6780 1930 6800 1940
rect 7730 1930 7780 1940
rect 9650 1930 9660 1940
rect 9860 1930 9870 1940
rect 9900 1930 9910 1940
rect 680 1920 920 1930
rect 1840 1920 1850 1930
rect 3320 1920 3350 1930
rect 4380 1920 4490 1930
rect 4600 1920 4610 1930
rect 4640 1920 4780 1930
rect 4870 1920 4980 1930
rect 6180 1920 6340 1930
rect 6520 1920 6570 1930
rect 6780 1920 6800 1930
rect 7730 1920 7770 1930
rect 670 1910 920 1920
rect 1840 1910 1850 1920
rect 3320 1910 3350 1920
rect 4410 1910 4480 1920
rect 4570 1910 4590 1920
rect 4610 1910 4620 1920
rect 4650 1910 4770 1920
rect 4880 1910 4970 1920
rect 6180 1910 6340 1920
rect 6530 1910 6570 1920
rect 6780 1910 6800 1920
rect 7730 1910 7790 1920
rect 9690 1910 9710 1920
rect 9900 1910 9910 1920
rect 9970 1910 9980 1920
rect 670 1900 920 1910
rect 1840 1900 1850 1910
rect 2660 1900 2680 1910
rect 3320 1900 3350 1910
rect 4390 1900 4400 1910
rect 4410 1900 4420 1910
rect 4430 1900 4480 1910
rect 4500 1900 4520 1910
rect 4540 1900 4630 1910
rect 4650 1900 4770 1910
rect 4800 1900 4850 1910
rect 4870 1900 4970 1910
rect 5010 1900 5020 1910
rect 5030 1900 5040 1910
rect 6150 1900 6160 1910
rect 6180 1900 6340 1910
rect 6540 1900 6580 1910
rect 6780 1900 6800 1910
rect 7730 1900 7780 1910
rect 9720 1900 9730 1910
rect 9950 1900 9960 1910
rect 9970 1900 9980 1910
rect 660 1890 920 1900
rect 1840 1890 1850 1900
rect 2550 1890 2560 1900
rect 2570 1890 2700 1900
rect 3320 1890 3350 1900
rect 4350 1890 4360 1900
rect 4420 1890 4480 1900
rect 4500 1890 4540 1900
rect 4550 1890 4560 1900
rect 4570 1890 4630 1900
rect 4650 1890 4770 1900
rect 4800 1890 4810 1900
rect 4820 1890 4850 1900
rect 4870 1890 4880 1900
rect 4890 1890 4960 1900
rect 5000 1890 5020 1900
rect 5030 1890 5050 1900
rect 6150 1890 6160 1900
rect 6180 1890 6340 1900
rect 6550 1890 6590 1900
rect 6780 1890 6790 1900
rect 7740 1890 7790 1900
rect 9740 1890 9750 1900
rect 660 1880 910 1890
rect 1840 1880 1850 1890
rect 2480 1880 2720 1890
rect 3320 1880 3350 1890
rect 4330 1880 4340 1890
rect 4400 1880 4410 1890
rect 4420 1880 4480 1890
rect 4500 1880 4550 1890
rect 4580 1880 4630 1890
rect 4650 1880 4760 1890
rect 4800 1880 4810 1890
rect 4820 1880 4850 1890
rect 4870 1880 4880 1890
rect 4900 1880 4910 1890
rect 4920 1880 4950 1890
rect 5020 1880 5040 1890
rect 6150 1880 6160 1890
rect 6180 1880 6350 1890
rect 6480 1880 6490 1890
rect 6500 1880 6540 1890
rect 6560 1880 6570 1890
rect 6790 1880 6800 1890
rect 7740 1880 7780 1890
rect 9680 1880 9690 1890
rect 650 1870 920 1880
rect 1840 1870 1860 1880
rect 2470 1870 2600 1880
rect 2620 1870 2750 1880
rect 3320 1870 3340 1880
rect 4310 1870 4320 1880
rect 4350 1870 4360 1880
rect 4390 1870 4400 1880
rect 4420 1870 4470 1880
rect 4500 1870 4540 1880
rect 4610 1870 4630 1880
rect 4650 1870 4760 1880
rect 4790 1870 4800 1880
rect 4810 1870 4850 1880
rect 4870 1870 4880 1880
rect 4900 1870 4910 1880
rect 4930 1870 4960 1880
rect 5090 1870 5100 1880
rect 5110 1870 5120 1880
rect 6170 1870 6350 1880
rect 6460 1870 6550 1880
rect 6570 1870 6580 1880
rect 6790 1870 6800 1880
rect 7740 1870 7790 1880
rect 9990 1870 9990 1880
rect 650 1860 920 1870
rect 1850 1860 1860 1870
rect 2440 1860 2800 1870
rect 3310 1860 3340 1870
rect 4280 1860 4290 1870
rect 4330 1860 4340 1870
rect 4410 1860 4420 1870
rect 4430 1860 4470 1870
rect 4510 1860 4540 1870
rect 4580 1860 4590 1870
rect 4600 1860 4630 1870
rect 4650 1860 4760 1870
rect 4790 1860 4800 1870
rect 4810 1860 4850 1870
rect 4870 1860 4880 1870
rect 4900 1860 4910 1870
rect 4920 1860 4950 1870
rect 5000 1860 5010 1870
rect 5140 1860 5150 1870
rect 6140 1860 6170 1870
rect 6180 1860 6350 1870
rect 6460 1860 6560 1870
rect 6570 1860 6590 1870
rect 6790 1860 6800 1870
rect 7740 1860 7790 1870
rect 9190 1860 9200 1870
rect 9270 1860 9280 1870
rect 9320 1860 9340 1870
rect 640 1850 910 1860
rect 1840 1850 1850 1860
rect 2420 1850 2530 1860
rect 2560 1850 2780 1860
rect 2790 1850 2830 1860
rect 3310 1850 3340 1860
rect 4280 1850 4290 1860
rect 4310 1850 4320 1860
rect 4350 1850 4360 1860
rect 4390 1850 4400 1860
rect 4430 1850 4470 1860
rect 4510 1850 4530 1860
rect 4550 1850 4580 1860
rect 4610 1850 4630 1860
rect 4650 1850 4750 1860
rect 4780 1850 4850 1860
rect 4870 1850 4890 1860
rect 4920 1850 4950 1860
rect 5040 1850 5050 1860
rect 6130 1850 6290 1860
rect 6320 1850 6330 1860
rect 6450 1850 6600 1860
rect 6790 1850 6800 1860
rect 7740 1850 7790 1860
rect 8380 1850 8390 1860
rect 9190 1850 9200 1860
rect 9330 1850 9340 1860
rect 9730 1850 9750 1860
rect 9760 1850 9770 1860
rect 640 1840 910 1850
rect 1850 1840 1860 1850
rect 2390 1840 2520 1850
rect 2580 1840 2760 1850
rect 2820 1840 2850 1850
rect 3310 1840 3340 1850
rect 4420 1840 4480 1850
rect 4510 1840 4530 1850
rect 4550 1840 4580 1850
rect 4610 1840 4630 1850
rect 4650 1840 4750 1850
rect 4780 1840 4790 1850
rect 4810 1840 4850 1850
rect 4870 1840 4900 1850
rect 4930 1840 4940 1850
rect 5140 1840 5150 1850
rect 6110 1840 6280 1850
rect 6460 1840 6610 1850
rect 6790 1840 6810 1850
rect 7740 1840 7790 1850
rect 8370 1840 8380 1850
rect 8400 1840 8410 1850
rect 9180 1840 9190 1850
rect 9200 1840 9210 1850
rect 9310 1840 9320 1850
rect 9690 1840 9700 1850
rect 9760 1840 9770 1850
rect 9970 1840 9980 1850
rect 630 1830 910 1840
rect 2380 1830 2530 1840
rect 2550 1830 2710 1840
rect 2850 1830 2880 1840
rect 3310 1830 3340 1840
rect 4270 1830 4280 1840
rect 4430 1830 4480 1840
rect 4510 1830 4530 1840
rect 4550 1830 4580 1840
rect 4600 1830 4630 1840
rect 4650 1830 4740 1840
rect 4780 1830 4790 1840
rect 4810 1830 4850 1840
rect 4880 1830 4890 1840
rect 4930 1830 4940 1840
rect 5100 1830 5110 1840
rect 5120 1830 5140 1840
rect 5260 1830 5270 1840
rect 6080 1830 6270 1840
rect 6460 1830 6560 1840
rect 6590 1830 6620 1840
rect 6790 1830 6810 1840
rect 7750 1830 7790 1840
rect 8370 1830 8380 1840
rect 8400 1830 8410 1840
rect 9110 1830 9120 1840
rect 9200 1830 9210 1840
rect 9320 1830 9330 1840
rect 9760 1830 9770 1840
rect 630 1820 910 1830
rect 2350 1820 2430 1830
rect 2440 1820 2500 1830
rect 2540 1820 2560 1830
rect 2860 1820 2880 1830
rect 3310 1820 3330 1830
rect 4420 1820 4470 1830
rect 4510 1820 4530 1830
rect 4550 1820 4580 1830
rect 4600 1820 4630 1830
rect 4650 1820 4740 1830
rect 4770 1820 4790 1830
rect 4820 1820 4850 1830
rect 4900 1820 4910 1830
rect 5090 1820 5100 1830
rect 5190 1820 5200 1830
rect 6080 1820 6280 1830
rect 6470 1820 6570 1830
rect 6610 1820 6630 1830
rect 6790 1820 6800 1830
rect 7340 1820 7350 1830
rect 7740 1820 7780 1830
rect 9190 1820 9200 1830
rect 9290 1820 9310 1830
rect 9380 1820 9390 1830
rect 9760 1820 9770 1830
rect 9980 1820 9990 1830
rect 630 1810 900 1820
rect 1850 1810 1860 1820
rect 2330 1810 2360 1820
rect 2410 1810 2430 1820
rect 2820 1810 2840 1820
rect 3300 1810 3330 1820
rect 4340 1810 4350 1820
rect 4420 1810 4480 1820
rect 4510 1810 4530 1820
rect 4540 1810 4560 1820
rect 4610 1810 4630 1820
rect 4650 1810 4740 1820
rect 4770 1810 4790 1820
rect 4830 1810 4840 1820
rect 4850 1810 4860 1820
rect 4880 1810 4890 1820
rect 4900 1810 4910 1820
rect 4970 1810 5000 1820
rect 5030 1810 5040 1820
rect 5190 1810 5200 1820
rect 5300 1810 5310 1820
rect 6080 1810 6280 1820
rect 6500 1810 6560 1820
rect 6790 1810 6800 1820
rect 7340 1810 7350 1820
rect 7750 1810 7790 1820
rect 8370 1810 8390 1820
rect 9270 1810 9280 1820
rect 9760 1810 9770 1820
rect 620 1800 900 1810
rect 2310 1800 2330 1810
rect 2460 1800 2500 1810
rect 2790 1800 2800 1810
rect 3300 1800 3330 1810
rect 4270 1800 4280 1810
rect 4290 1800 4300 1810
rect 4420 1800 4440 1810
rect 4450 1800 4480 1810
rect 4510 1800 4540 1810
rect 4590 1800 4620 1810
rect 4640 1800 4740 1810
rect 4770 1800 4780 1810
rect 4840 1800 4850 1810
rect 4880 1800 4890 1810
rect 4900 1800 4910 1810
rect 4920 1800 4930 1810
rect 4980 1800 5000 1810
rect 5030 1800 5040 1810
rect 5080 1800 5090 1810
rect 5180 1800 5190 1810
rect 5230 1800 5240 1810
rect 6070 1800 6280 1810
rect 6510 1800 6580 1810
rect 6790 1800 6800 1810
rect 7750 1800 7790 1810
rect 8370 1800 8380 1810
rect 8390 1800 8400 1810
rect 9250 1800 9270 1810
rect 9400 1800 9410 1810
rect 9450 1800 9460 1810
rect 9950 1800 9960 1810
rect 9970 1800 9980 1810
rect 620 1790 900 1800
rect 1850 1790 1860 1800
rect 2300 1790 2330 1800
rect 2390 1790 2460 1800
rect 2520 1790 2550 1800
rect 2570 1790 2710 1800
rect 3300 1790 3320 1800
rect 4290 1790 4300 1800
rect 4360 1790 4370 1800
rect 4390 1790 4400 1800
rect 4420 1790 4430 1800
rect 4440 1790 4480 1800
rect 4510 1790 4540 1800
rect 4550 1790 4560 1800
rect 4570 1790 4610 1800
rect 4650 1790 4730 1800
rect 4760 1790 4780 1800
rect 4840 1790 4850 1800
rect 4880 1790 4890 1800
rect 4950 1790 4980 1800
rect 5220 1790 5230 1800
rect 5250 1790 5260 1800
rect 6040 1790 6050 1800
rect 6070 1790 6290 1800
rect 6520 1790 6590 1800
rect 6790 1790 6810 1800
rect 7750 1790 7790 1800
rect 8370 1790 8400 1800
rect 9240 1790 9260 1800
rect 9760 1790 9770 1800
rect 610 1780 890 1790
rect 1850 1780 1870 1790
rect 2340 1780 2420 1790
rect 3290 1780 3320 1790
rect 4290 1780 4300 1790
rect 4400 1780 4410 1790
rect 4420 1780 4480 1790
rect 4510 1780 4610 1790
rect 4650 1780 4730 1790
rect 4760 1780 4780 1790
rect 4880 1780 4890 1790
rect 5070 1780 5080 1790
rect 5170 1780 5180 1790
rect 5220 1780 5230 1790
rect 6050 1780 6290 1790
rect 6550 1780 6600 1790
rect 6790 1780 6810 1790
rect 7750 1780 7800 1790
rect 8360 1780 8400 1790
rect 9740 1780 9770 1790
rect 9910 1780 9920 1790
rect 9960 1780 9970 1790
rect 610 1770 900 1780
rect 1860 1770 1870 1780
rect 3290 1770 3320 1780
rect 4360 1770 4370 1780
rect 4380 1770 4390 1780
rect 4430 1770 4480 1780
rect 4510 1770 4610 1780
rect 4650 1770 4720 1780
rect 4840 1770 4850 1780
rect 5020 1770 5030 1780
rect 5170 1770 5180 1780
rect 5210 1770 5240 1780
rect 5340 1770 5350 1780
rect 6050 1770 6300 1780
rect 6550 1770 6620 1780
rect 6800 1770 6810 1780
rect 7760 1770 7810 1780
rect 8360 1770 8400 1780
rect 9220 1770 9230 1780
rect 9740 1770 9780 1780
rect 9930 1770 9940 1780
rect 610 1760 890 1770
rect 1860 1760 1880 1770
rect 3290 1760 3320 1770
rect 4340 1760 4360 1770
rect 4400 1760 4410 1770
rect 4420 1760 4450 1770
rect 4460 1760 4480 1770
rect 4500 1760 4610 1770
rect 4640 1760 4690 1770
rect 4710 1760 4720 1770
rect 4750 1760 4760 1770
rect 4800 1760 4810 1770
rect 4830 1760 4860 1770
rect 4950 1760 4960 1770
rect 5200 1760 5210 1770
rect 5230 1760 5240 1770
rect 5340 1760 5350 1770
rect 6040 1760 6310 1770
rect 6550 1760 6620 1770
rect 6800 1760 6810 1770
rect 7760 1760 7810 1770
rect 8360 1760 8370 1770
rect 9210 1760 9220 1770
rect 9700 1760 9710 1770
rect 9740 1760 9780 1770
rect 9950 1760 9960 1770
rect 600 1750 890 1760
rect 1870 1750 1880 1760
rect 3280 1750 3310 1760
rect 4280 1750 4290 1760
rect 4380 1750 4390 1760
rect 4400 1750 4410 1760
rect 4430 1750 4450 1760
rect 4460 1750 4480 1760
rect 4510 1750 4540 1760
rect 4570 1750 4620 1760
rect 4640 1750 4700 1760
rect 4750 1750 4760 1760
rect 4820 1750 4840 1760
rect 4920 1750 4930 1760
rect 4950 1750 4960 1760
rect 5060 1750 5070 1760
rect 5160 1750 5170 1760
rect 5200 1750 5210 1760
rect 5220 1750 5230 1760
rect 5340 1750 5350 1760
rect 6050 1750 6320 1760
rect 6550 1750 6620 1760
rect 6800 1750 6810 1760
rect 7760 1750 7800 1760
rect 8360 1750 8390 1760
rect 9740 1750 9760 1760
rect 600 1740 890 1750
rect 1870 1740 1880 1750
rect 3280 1740 3310 1750
rect 4280 1740 4290 1750
rect 4360 1740 4370 1750
rect 4400 1740 4410 1750
rect 4430 1740 4480 1750
rect 4500 1740 4530 1750
rect 4580 1740 4620 1750
rect 4650 1740 4710 1750
rect 4750 1740 4760 1750
rect 4770 1740 4780 1750
rect 4940 1740 4960 1750
rect 5060 1740 5070 1750
rect 5150 1740 5160 1750
rect 5190 1740 5200 1750
rect 5430 1740 5440 1750
rect 6030 1740 6310 1750
rect 6550 1740 6640 1750
rect 6800 1740 6810 1750
rect 7770 1740 7810 1750
rect 8360 1740 8390 1750
rect 9110 1740 9120 1750
rect 9740 1740 9760 1750
rect 9840 1740 9850 1750
rect 9920 1740 9930 1750
rect 9940 1740 9950 1750
rect 590 1730 880 1740
rect 1870 1730 1880 1740
rect 3280 1730 3310 1740
rect 4280 1730 4290 1740
rect 4300 1730 4310 1740
rect 4430 1730 4480 1740
rect 4500 1730 4530 1740
rect 4580 1730 4620 1740
rect 4650 1730 4700 1740
rect 4740 1730 4750 1740
rect 4800 1730 4830 1740
rect 4950 1730 4960 1740
rect 5060 1730 5070 1740
rect 5190 1730 5200 1740
rect 5210 1730 5220 1740
rect 5330 1730 5340 1740
rect 5420 1730 5430 1740
rect 6030 1730 6310 1740
rect 6510 1730 6530 1740
rect 6550 1730 6660 1740
rect 6800 1730 6810 1740
rect 7770 1730 7800 1740
rect 8370 1730 8390 1740
rect 9110 1730 9120 1740
rect 9740 1730 9760 1740
rect 9840 1730 9860 1740
rect 590 1720 880 1730
rect 1880 1720 1890 1730
rect 3280 1720 3300 1730
rect 4280 1720 4290 1730
rect 4300 1720 4310 1730
rect 4430 1720 4480 1730
rect 4510 1720 4530 1730
rect 4590 1720 4630 1730
rect 4660 1720 4700 1730
rect 4740 1720 4760 1730
rect 4830 1720 4840 1730
rect 4950 1720 4970 1730
rect 5050 1720 5060 1730
rect 5180 1720 5190 1730
rect 5310 1720 5320 1730
rect 5400 1720 5410 1730
rect 5990 1720 6000 1730
rect 6030 1720 6320 1730
rect 6490 1720 6510 1730
rect 6540 1720 6670 1730
rect 6800 1720 6810 1730
rect 7770 1720 7810 1730
rect 8370 1720 8390 1730
rect 9110 1720 9120 1730
rect 9190 1720 9200 1730
rect 9740 1720 9760 1730
rect 9780 1720 9790 1730
rect 9830 1720 9840 1730
rect 9920 1720 9930 1730
rect 590 1710 880 1720
rect 1880 1710 1900 1720
rect 3270 1710 3300 1720
rect 4430 1710 4480 1720
rect 4500 1710 4530 1720
rect 4550 1710 4570 1720
rect 4590 1710 4630 1720
rect 4660 1710 4700 1720
rect 4730 1710 4760 1720
rect 4920 1710 4930 1720
rect 5000 1710 5010 1720
rect 5050 1710 5060 1720
rect 5180 1710 5190 1720
rect 5260 1710 5270 1720
rect 5990 1710 6020 1720
rect 6050 1710 6200 1720
rect 6230 1710 6320 1720
rect 6490 1710 6500 1720
rect 6540 1710 6670 1720
rect 6800 1710 6810 1720
rect 7350 1710 7360 1720
rect 7760 1710 7810 1720
rect 8370 1710 8390 1720
rect 9110 1710 9120 1720
rect 9740 1710 9750 1720
rect 9900 1710 9910 1720
rect 580 1700 870 1710
rect 1880 1700 1890 1710
rect 3260 1700 3290 1710
rect 4400 1700 4480 1710
rect 4500 1700 4530 1710
rect 4550 1700 4570 1710
rect 4600 1700 4640 1710
rect 4660 1700 4700 1710
rect 4730 1700 4750 1710
rect 5030 1700 5040 1710
rect 5170 1700 5180 1710
rect 5190 1700 5200 1710
rect 5300 1700 5320 1710
rect 6010 1700 6210 1710
rect 6230 1700 6330 1710
rect 6540 1700 6670 1710
rect 6800 1700 6810 1710
rect 7760 1700 7820 1710
rect 8360 1700 8380 1710
rect 9110 1700 9120 1710
rect 9200 1700 9210 1710
rect 9740 1700 9760 1710
rect 9780 1700 9790 1710
rect 9910 1700 9920 1710
rect 580 1690 870 1700
rect 1880 1690 1900 1700
rect 3260 1690 3290 1700
rect 4340 1690 4350 1700
rect 4400 1690 4480 1700
rect 4510 1690 4530 1700
rect 4550 1690 4580 1700
rect 4600 1690 4640 1700
rect 4670 1690 4690 1700
rect 4730 1690 4750 1700
rect 4790 1690 4810 1700
rect 4840 1690 4850 1700
rect 4890 1690 4900 1700
rect 4990 1690 5000 1700
rect 5170 1690 5180 1700
rect 5250 1690 5260 1700
rect 5450 1690 5460 1700
rect 6000 1690 6210 1700
rect 6240 1690 6330 1700
rect 6530 1690 6660 1700
rect 6800 1690 6810 1700
rect 7770 1690 7810 1700
rect 8360 1690 8390 1700
rect 9740 1690 9760 1700
rect 9780 1690 9790 1700
rect 9890 1690 9900 1700
rect 9910 1690 9920 1700
rect 570 1680 870 1690
rect 1880 1680 1900 1690
rect 3260 1680 3280 1690
rect 4340 1680 4350 1690
rect 4390 1680 4420 1690
rect 4440 1680 4480 1690
rect 4510 1680 4580 1690
rect 4610 1680 4640 1690
rect 4670 1680 4690 1690
rect 4720 1680 4750 1690
rect 4770 1680 4790 1690
rect 4840 1680 4850 1690
rect 4890 1680 4900 1690
rect 5040 1680 5050 1690
rect 5160 1680 5170 1690
rect 5180 1680 5190 1690
rect 5290 1680 5300 1690
rect 5980 1680 6000 1690
rect 6020 1680 6200 1690
rect 6250 1680 6330 1690
rect 6480 1680 6490 1690
rect 6520 1680 6660 1690
rect 6800 1680 6810 1690
rect 7770 1680 7810 1690
rect 8360 1680 8390 1690
rect 9200 1680 9210 1690
rect 9740 1680 9760 1690
rect 9780 1680 9790 1690
rect 570 1670 870 1680
rect 1890 1670 1900 1680
rect 3250 1670 3280 1680
rect 4070 1670 4080 1680
rect 4290 1670 4300 1680
rect 4340 1670 4360 1680
rect 4450 1670 4480 1680
rect 4510 1670 4530 1680
rect 4560 1670 4590 1680
rect 4610 1670 4650 1680
rect 4670 1670 4690 1680
rect 4720 1670 4740 1680
rect 4770 1670 4790 1680
rect 4840 1670 4870 1680
rect 5240 1670 5250 1680
rect 5300 1670 5310 1680
rect 5370 1670 5380 1680
rect 6010 1670 6020 1680
rect 6040 1670 6200 1680
rect 6250 1670 6330 1680
rect 6510 1670 6650 1680
rect 6800 1670 6810 1680
rect 7770 1670 7810 1680
rect 8340 1670 8390 1680
rect 9750 1670 9770 1680
rect 9790 1670 9800 1680
rect 570 1660 870 1670
rect 1890 1660 1910 1670
rect 3240 1660 3270 1670
rect 4290 1660 4300 1670
rect 4410 1660 4430 1670
rect 4460 1660 4480 1670
rect 4550 1660 4590 1670
rect 4640 1660 4650 1670
rect 4670 1660 4690 1670
rect 4720 1660 4730 1670
rect 4760 1660 4790 1670
rect 4890 1660 4900 1670
rect 4910 1660 4930 1670
rect 5030 1660 5040 1670
rect 5280 1660 5300 1670
rect 5430 1660 5450 1670
rect 5960 1660 5970 1670
rect 5980 1660 5990 1670
rect 6010 1660 6030 1670
rect 6040 1660 6200 1670
rect 6260 1660 6330 1670
rect 6500 1660 6650 1670
rect 6800 1660 6810 1670
rect 7770 1660 7810 1670
rect 8340 1660 8390 1670
rect 9740 1660 9780 1670
rect 9890 1660 9900 1670
rect 560 1650 870 1660
rect 1890 1650 1910 1660
rect 3240 1650 3260 1660
rect 4290 1650 4300 1660
rect 4310 1650 4320 1660
rect 4380 1650 4400 1660
rect 4430 1650 4440 1660
rect 4450 1650 4460 1660
rect 4470 1650 4480 1660
rect 4530 1650 4540 1660
rect 4550 1650 4600 1660
rect 4650 1650 4660 1660
rect 4670 1650 4690 1660
rect 4770 1650 4780 1660
rect 4890 1650 4940 1660
rect 4980 1650 4990 1660
rect 5030 1650 5040 1660
rect 5230 1650 5240 1660
rect 5430 1650 5440 1660
rect 5980 1650 6000 1660
rect 6010 1650 6200 1660
rect 6260 1650 6340 1660
rect 6500 1650 6650 1660
rect 6800 1650 6820 1660
rect 7770 1650 7810 1660
rect 8340 1650 8400 1660
rect 9880 1650 9890 1660
rect 560 1640 870 1650
rect 1900 1640 1920 1650
rect 3240 1640 3260 1650
rect 4080 1640 4090 1650
rect 4310 1640 4320 1650
rect 4450 1640 4460 1650
rect 4470 1640 4480 1650
rect 4550 1640 4620 1650
rect 4670 1640 4680 1650
rect 4760 1640 4770 1650
rect 4800 1640 4810 1650
rect 4920 1640 4930 1650
rect 5020 1640 5040 1650
rect 5230 1640 5240 1650
rect 5270 1640 5280 1650
rect 5940 1640 5960 1650
rect 5980 1640 6200 1650
rect 6270 1640 6340 1650
rect 6490 1640 6500 1650
rect 6510 1640 6650 1650
rect 6800 1640 6810 1650
rect 7770 1640 7820 1650
rect 8340 1640 8370 1650
rect 9880 1640 9890 1650
rect 560 1630 870 1640
rect 1910 1630 1920 1640
rect 3230 1630 3260 1640
rect 4270 1630 4280 1640
rect 4310 1630 4320 1640
rect 4390 1630 4420 1640
rect 4470 1630 4500 1640
rect 4550 1630 4620 1640
rect 4660 1630 4700 1640
rect 4750 1630 4760 1640
rect 4780 1630 4810 1640
rect 4840 1630 4850 1640
rect 4880 1630 4900 1640
rect 5020 1630 5030 1640
rect 5210 1630 5230 1640
rect 5280 1630 5290 1640
rect 5950 1630 5960 1640
rect 6000 1630 6200 1640
rect 6270 1630 6340 1640
rect 6500 1630 6660 1640
rect 6800 1630 6820 1640
rect 7770 1630 7820 1640
rect 8330 1630 8370 1640
rect 550 1620 860 1630
rect 1910 1620 1920 1630
rect 3220 1620 3250 1630
rect 4370 1620 4380 1630
rect 4470 1620 4500 1630
rect 4540 1620 4660 1630
rect 4670 1620 4720 1630
rect 4760 1620 4800 1630
rect 4970 1620 4990 1630
rect 5010 1620 5030 1630
rect 5190 1620 5210 1630
rect 5540 1620 5550 1630
rect 5990 1620 6200 1630
rect 6280 1620 6330 1630
rect 6490 1620 6680 1630
rect 6800 1620 6810 1630
rect 7770 1620 7820 1630
rect 8330 1620 8380 1630
rect 9240 1620 9250 1630
rect 9870 1620 9880 1630
rect 550 1610 860 1620
rect 1920 1610 1930 1620
rect 3220 1610 3250 1620
rect 4090 1610 4100 1620
rect 4280 1610 4290 1620
rect 4400 1610 4410 1620
rect 4470 1610 4720 1620
rect 4750 1610 4800 1620
rect 4810 1610 4820 1620
rect 4980 1610 4990 1620
rect 5020 1610 5030 1620
rect 5270 1610 5280 1620
rect 5430 1610 5440 1620
rect 5970 1610 6210 1620
rect 6280 1610 6330 1620
rect 6480 1610 6700 1620
rect 6800 1610 6810 1620
rect 7780 1610 7820 1620
rect 8350 1610 8390 1620
rect 9120 1610 9130 1620
rect 9180 1610 9210 1620
rect 540 1600 860 1610
rect 1920 1600 1930 1610
rect 3210 1600 3240 1610
rect 4350 1600 4360 1610
rect 4460 1600 4810 1610
rect 5170 1600 5190 1610
rect 5530 1600 5540 1610
rect 5970 1600 6210 1610
rect 6280 1600 6330 1610
rect 6440 1600 6710 1610
rect 6800 1600 6820 1610
rect 7360 1600 7370 1610
rect 7780 1600 7830 1610
rect 8330 1600 8380 1610
rect 9150 1600 9160 1610
rect 540 1590 860 1600
rect 1920 1590 1930 1600
rect 3200 1590 3230 1600
rect 4320 1590 4330 1600
rect 4450 1590 4570 1600
rect 4840 1590 4900 1600
rect 5140 1590 5150 1600
rect 5240 1590 5250 1600
rect 5510 1590 5530 1600
rect 5960 1590 6210 1600
rect 6280 1590 6340 1600
rect 6440 1590 6720 1600
rect 6800 1590 6810 1600
rect 7360 1590 7370 1600
rect 7780 1590 7820 1600
rect 8330 1590 8390 1600
rect 9860 1590 9870 1600
rect 540 1580 850 1590
rect 1930 1580 1940 1590
rect 3200 1580 3220 1590
rect 4100 1580 4110 1590
rect 4300 1580 4310 1590
rect 4420 1580 4500 1590
rect 4610 1580 4660 1590
rect 4700 1580 4730 1590
rect 4800 1580 4850 1590
rect 4940 1580 4960 1590
rect 5220 1580 5230 1590
rect 5300 1580 5310 1590
rect 5380 1580 5400 1590
rect 5960 1580 6210 1590
rect 6280 1580 6330 1590
rect 6430 1580 6730 1590
rect 6800 1580 6810 1590
rect 7790 1580 7820 1590
rect 8320 1580 8380 1590
rect 530 1570 850 1580
rect 1940 1570 1950 1580
rect 3190 1570 3220 1580
rect 4390 1570 4440 1580
rect 4520 1570 4700 1580
rect 4740 1570 4790 1580
rect 4930 1570 4960 1580
rect 4990 1570 5000 1580
rect 5160 1570 5200 1580
rect 5230 1570 5240 1580
rect 5370 1570 5380 1580
rect 5410 1570 5420 1580
rect 5430 1570 5460 1580
rect 5480 1570 5500 1580
rect 5970 1570 6220 1580
rect 6280 1570 6340 1580
rect 6420 1570 6730 1580
rect 6800 1570 6810 1580
rect 7780 1570 7820 1580
rect 8320 1570 8390 1580
rect 9840 1570 9850 1580
rect 9920 1570 9940 1580
rect 9980 1570 9990 1580
rect 530 1560 850 1570
rect 1940 1560 1950 1570
rect 3180 1560 3210 1570
rect 4490 1560 4710 1570
rect 4730 1560 4780 1570
rect 4790 1560 4800 1570
rect 4830 1560 4840 1570
rect 4980 1560 4990 1570
rect 5030 1560 5060 1570
rect 5350 1560 5370 1570
rect 5430 1560 5480 1570
rect 5960 1560 6220 1570
rect 6290 1560 6340 1570
rect 6400 1560 6730 1570
rect 6790 1560 6800 1570
rect 7780 1560 7830 1570
rect 8320 1560 8390 1570
rect 9740 1560 9800 1570
rect 9910 1560 9930 1570
rect 530 1550 840 1560
rect 1950 1550 1960 1560
rect 3180 1550 3210 1560
rect 4460 1550 4810 1560
rect 4830 1550 4850 1560
rect 4990 1550 5000 1560
rect 5030 1550 5050 1560
rect 5080 1550 5100 1560
rect 5300 1550 5310 1560
rect 5330 1550 5340 1560
rect 5350 1550 5360 1560
rect 5630 1550 5640 1560
rect 5810 1550 5820 1560
rect 5980 1550 6220 1560
rect 6290 1550 6330 1560
rect 6400 1550 6730 1560
rect 6790 1550 6810 1560
rect 7790 1550 7840 1560
rect 8320 1550 8390 1560
rect 9810 1550 9820 1560
rect 9830 1550 9840 1560
rect 9910 1550 9930 1560
rect 520 1540 840 1550
rect 1960 1540 1970 1550
rect 3170 1540 3200 1550
rect 4430 1540 4440 1550
rect 4460 1540 4820 1550
rect 4980 1540 5000 1550
rect 5070 1540 5100 1550
rect 5110 1540 5120 1550
rect 5340 1540 5350 1550
rect 5680 1540 5700 1550
rect 5960 1540 6230 1550
rect 6290 1540 6340 1550
rect 6410 1540 6730 1550
rect 6790 1540 6800 1550
rect 7790 1540 7840 1550
rect 8310 1540 8370 1550
rect 9790 1540 9800 1550
rect 9830 1540 9840 1550
rect 520 1530 840 1540
rect 1960 1530 1970 1540
rect 3160 1530 3190 1540
rect 4410 1530 4440 1540
rect 4470 1530 4870 1540
rect 4890 1530 4910 1540
rect 4920 1530 4940 1540
rect 4980 1530 5000 1540
rect 5120 1530 5150 1540
rect 5580 1530 5590 1540
rect 5640 1530 5660 1540
rect 5680 1530 5700 1540
rect 5920 1530 5930 1540
rect 5960 1530 5970 1540
rect 5980 1530 6230 1540
rect 6300 1530 6340 1540
rect 6410 1530 6730 1540
rect 6790 1530 6800 1540
rect 7790 1530 7830 1540
rect 8310 1530 8380 1540
rect 9800 1530 9810 1540
rect 9820 1530 9830 1540
rect 9930 1530 9940 1540
rect 9950 1530 9960 1540
rect 520 1520 830 1530
rect 1970 1520 1980 1530
rect 3150 1520 3180 1530
rect 4130 1520 4140 1530
rect 4400 1520 4440 1530
rect 4470 1520 4910 1530
rect 4920 1520 4950 1530
rect 4970 1520 5000 1530
rect 5140 1520 5180 1530
rect 5330 1520 5340 1530
rect 5580 1520 5600 1530
rect 5630 1520 5640 1530
rect 5680 1520 5700 1530
rect 5880 1520 5890 1530
rect 5960 1520 5970 1530
rect 5980 1520 5990 1530
rect 6010 1520 6200 1530
rect 6220 1520 6230 1530
rect 6300 1520 6340 1530
rect 6400 1520 6730 1530
rect 6790 1520 6800 1530
rect 7370 1520 7380 1530
rect 7790 1520 7840 1530
rect 8310 1520 8370 1530
rect 9780 1520 9790 1530
rect 9940 1520 9950 1530
rect 510 1510 840 1520
rect 1980 1510 1990 1520
rect 3140 1510 3170 1520
rect 4340 1510 4350 1520
rect 4390 1510 4450 1520
rect 4470 1510 4960 1520
rect 4980 1510 5000 1520
rect 5170 1510 5200 1520
rect 5310 1510 5330 1520
rect 5580 1510 5600 1520
rect 5680 1510 5690 1520
rect 5940 1510 5950 1520
rect 5960 1510 6200 1520
rect 6220 1510 6240 1520
rect 6300 1510 6340 1520
rect 6380 1510 6760 1520
rect 6790 1510 6800 1520
rect 7370 1510 7380 1520
rect 7800 1510 7830 1520
rect 8310 1510 8380 1520
rect 9820 1510 9830 1520
rect 510 1500 830 1510
rect 3120 1500 3160 1510
rect 4130 1500 4140 1510
rect 4360 1500 4380 1510
rect 4390 1500 4450 1510
rect 4470 1500 4930 1510
rect 4980 1500 5000 1510
rect 5190 1500 5230 1510
rect 5580 1500 5600 1510
rect 5720 1500 5730 1510
rect 5940 1500 6200 1510
rect 6300 1500 6340 1510
rect 6380 1500 6760 1510
rect 6790 1500 6800 1510
rect 7800 1500 7840 1510
rect 8310 1500 8360 1510
rect 9130 1500 9140 1510
rect 9710 1500 9720 1510
rect 9770 1500 9790 1510
rect 9900 1500 9910 1510
rect 9980 1500 9990 1510
rect 510 1490 830 1500
rect 1990 1490 2000 1500
rect 3110 1490 3150 1500
rect 4370 1490 4450 1500
rect 4470 1490 4940 1500
rect 4950 1490 4960 1500
rect 4980 1490 5000 1500
rect 5010 1490 5020 1500
rect 5220 1490 5230 1500
rect 5240 1490 5250 1500
rect 5720 1490 5730 1500
rect 5960 1490 6200 1500
rect 6300 1490 6340 1500
rect 6380 1490 6770 1500
rect 6790 1490 6800 1500
rect 7800 1490 7830 1500
rect 8300 1490 8360 1500
rect 9350 1490 9370 1500
rect 9900 1490 9910 1500
rect 9920 1490 9930 1500
rect 500 1480 830 1490
rect 2000 1480 2010 1490
rect 3110 1480 3140 1490
rect 4380 1480 4440 1490
rect 4470 1480 4940 1490
rect 4950 1480 4960 1490
rect 4970 1480 4990 1490
rect 5010 1480 5020 1490
rect 5030 1480 5040 1490
rect 5070 1480 5090 1490
rect 5110 1480 5120 1490
rect 5240 1480 5250 1490
rect 5260 1480 5270 1490
rect 5580 1480 5590 1490
rect 5720 1480 5730 1490
rect 5850 1480 5880 1490
rect 5890 1480 5940 1490
rect 5960 1480 6200 1490
rect 6310 1480 6330 1490
rect 6370 1480 6770 1490
rect 6790 1480 6800 1490
rect 7800 1480 7830 1490
rect 8300 1480 8360 1490
rect 9180 1480 9190 1490
rect 9360 1480 9370 1490
rect 9760 1480 9780 1490
rect 9800 1480 9810 1490
rect 9910 1480 9920 1490
rect 500 1470 840 1480
rect 2010 1470 2020 1480
rect 3100 1470 3130 1480
rect 4380 1470 4440 1480
rect 4560 1470 4960 1480
rect 4970 1470 4980 1480
rect 5260 1470 5290 1480
rect 5470 1470 5490 1480
rect 5690 1470 5720 1480
rect 5870 1470 5880 1480
rect 5890 1470 6190 1480
rect 6310 1470 6330 1480
rect 6370 1470 6760 1480
rect 6790 1470 6800 1480
rect 7800 1470 7850 1480
rect 8310 1470 8370 1480
rect 9710 1470 9720 1480
rect 500 1460 840 1470
rect 900 1460 910 1470
rect 980 1460 990 1470
rect 2020 1460 2030 1470
rect 3090 1460 3120 1470
rect 4360 1460 4370 1470
rect 4380 1460 4390 1470
rect 4680 1460 4960 1470
rect 4970 1460 4980 1470
rect 5010 1460 5030 1470
rect 5280 1460 5300 1470
rect 5480 1460 5490 1470
rect 5700 1460 5720 1470
rect 5880 1460 6190 1470
rect 6300 1460 6330 1470
rect 6360 1460 6760 1470
rect 6790 1460 6800 1470
rect 7810 1460 7840 1470
rect 8300 1460 8370 1470
rect 9590 1460 9640 1470
rect 9750 1460 9760 1470
rect 490 1450 840 1460
rect 880 1450 890 1460
rect 990 1450 1000 1460
rect 2020 1450 2040 1460
rect 3070 1450 3110 1460
rect 4480 1450 4500 1460
rect 4520 1450 4540 1460
rect 4560 1450 4580 1460
rect 4600 1450 4620 1460
rect 4640 1450 4650 1460
rect 4680 1450 4690 1460
rect 4740 1450 4780 1460
rect 4830 1450 4840 1460
rect 4890 1450 4960 1460
rect 4970 1450 4990 1460
rect 5010 1450 5060 1460
rect 5080 1450 5100 1460
rect 5110 1450 5120 1460
rect 5290 1450 5300 1460
rect 5480 1450 5490 1460
rect 5890 1450 6200 1460
rect 6310 1450 6340 1460
rect 6360 1450 6780 1460
rect 7810 1450 7850 1460
rect 8300 1450 8370 1460
rect 9580 1450 9590 1460
rect 9630 1450 9640 1460
rect 9750 1450 9760 1460
rect 9780 1450 9790 1460
rect 490 1440 840 1450
rect 860 1440 870 1450
rect 1000 1440 1010 1450
rect 2030 1440 2040 1450
rect 3060 1440 3100 1450
rect 4430 1440 4450 1450
rect 4480 1440 4500 1450
rect 4520 1440 4540 1450
rect 4560 1440 4580 1450
rect 4600 1440 4620 1450
rect 4640 1440 4660 1450
rect 4670 1440 4690 1450
rect 4710 1440 4730 1450
rect 4790 1440 4830 1450
rect 4840 1440 4850 1450
rect 4880 1440 4890 1450
rect 4900 1440 4950 1450
rect 4980 1440 4990 1450
rect 5010 1440 5020 1450
rect 5030 1440 5050 1450
rect 5140 1440 5170 1450
rect 5220 1440 5230 1450
rect 5300 1440 5310 1450
rect 5580 1440 5600 1450
rect 5900 1440 6200 1450
rect 6310 1440 6330 1450
rect 6350 1440 6780 1450
rect 7380 1440 7390 1450
rect 7810 1440 7840 1450
rect 8300 1440 8360 1450
rect 9130 1440 9140 1450
rect 9630 1440 9640 1450
rect 490 1430 840 1440
rect 1010 1430 1020 1440
rect 2040 1430 2050 1440
rect 3050 1430 3090 1440
rect 4430 1430 4460 1440
rect 4470 1430 4500 1440
rect 4520 1430 4540 1440
rect 4560 1430 4580 1440
rect 4600 1430 4620 1440
rect 4630 1430 4650 1440
rect 4670 1430 4690 1440
rect 4710 1430 4730 1440
rect 4740 1430 4760 1440
rect 4830 1430 4840 1440
rect 4880 1430 4890 1440
rect 4900 1430 4950 1440
rect 4980 1430 4990 1440
rect 5000 1430 5070 1440
rect 5140 1430 5170 1440
rect 5310 1430 5320 1440
rect 5570 1430 5600 1440
rect 5890 1430 6200 1440
rect 6310 1430 6780 1440
rect 7380 1430 7390 1440
rect 7820 1430 7850 1440
rect 8300 1430 8360 1440
rect 9630 1430 9640 1440
rect 9730 1430 9740 1440
rect 480 1420 840 1430
rect 1010 1420 1020 1430
rect 2050 1420 2060 1430
rect 3040 1420 3080 1430
rect 4370 1420 4380 1430
rect 4400 1420 4410 1430
rect 4440 1420 4460 1430
rect 4470 1420 4500 1430
rect 4520 1420 4540 1430
rect 4560 1420 4580 1430
rect 4600 1420 4620 1430
rect 4630 1420 4640 1430
rect 4650 1420 4660 1430
rect 4670 1420 4690 1430
rect 4710 1420 4720 1430
rect 4740 1420 4760 1430
rect 4780 1420 4800 1430
rect 4810 1420 4820 1430
rect 4900 1420 4970 1430
rect 4990 1420 5100 1430
rect 5120 1420 5130 1430
rect 5150 1420 5160 1430
rect 5320 1420 5330 1430
rect 5340 1420 5350 1430
rect 5570 1420 5580 1430
rect 5890 1420 6200 1430
rect 6310 1420 6780 1430
rect 7820 1420 7860 1430
rect 8290 1420 8360 1430
rect 9520 1420 9550 1430
rect 9620 1420 9640 1430
rect 9760 1420 9770 1430
rect 480 1410 850 1420
rect 1000 1410 1030 1420
rect 2060 1410 2070 1420
rect 3030 1410 3070 1420
rect 4440 1410 4460 1420
rect 4480 1410 4500 1420
rect 4520 1410 4540 1420
rect 4560 1410 4580 1420
rect 4640 1410 4650 1420
rect 4680 1410 4690 1420
rect 4710 1410 4720 1420
rect 4740 1410 4760 1420
rect 4770 1410 4800 1420
rect 4830 1410 4840 1420
rect 4850 1410 4870 1420
rect 4890 1410 4900 1420
rect 4910 1410 4950 1420
rect 4960 1410 4980 1420
rect 5000 1410 5080 1420
rect 5090 1410 5110 1420
rect 5120 1410 5150 1420
rect 5340 1410 5350 1420
rect 5560 1410 5580 1420
rect 5620 1410 5630 1420
rect 5930 1410 6200 1420
rect 6310 1410 6790 1420
rect 7820 1410 7850 1420
rect 8290 1410 8360 1420
rect 9720 1410 9740 1420
rect 480 1400 850 1410
rect 990 1400 1030 1410
rect 2060 1400 2080 1410
rect 3020 1400 3060 1410
rect 4380 1400 4390 1410
rect 4440 1400 4460 1410
rect 4480 1400 4500 1410
rect 4520 1400 4530 1410
rect 4740 1400 4760 1410
rect 4770 1400 4790 1410
rect 4800 1400 4810 1410
rect 4830 1400 4850 1410
rect 4860 1400 4870 1410
rect 4890 1400 4950 1410
rect 4960 1400 4980 1410
rect 4990 1400 5070 1410
rect 5080 1400 5100 1410
rect 5180 1400 5190 1410
rect 5340 1400 5350 1410
rect 5360 1400 5370 1410
rect 5500 1400 5510 1410
rect 5550 1400 5570 1410
rect 5620 1400 5630 1410
rect 5890 1400 5900 1410
rect 5910 1400 6200 1410
rect 6310 1400 6790 1410
rect 6800 1400 6810 1410
rect 7820 1400 7860 1410
rect 8290 1400 8360 1410
rect 9240 1400 9250 1410
rect 9690 1400 9700 1410
rect 470 1390 840 1400
rect 990 1390 1030 1400
rect 2070 1390 2090 1400
rect 3000 1390 3050 1400
rect 4440 1390 4460 1400
rect 4550 1390 4680 1400
rect 4710 1390 4740 1400
rect 4780 1390 4790 1400
rect 4800 1390 4810 1400
rect 4820 1390 4830 1400
rect 4840 1390 4850 1400
rect 4860 1390 4870 1400
rect 4880 1390 4890 1400
rect 4900 1390 4930 1400
rect 4940 1390 4980 1400
rect 4990 1390 5090 1400
rect 5110 1390 5120 1400
rect 5170 1390 5190 1400
rect 5350 1390 5380 1400
rect 5510 1390 5560 1400
rect 5610 1390 5620 1400
rect 5890 1390 6200 1400
rect 6310 1390 6790 1400
rect 6800 1390 6810 1400
rect 7820 1390 7860 1400
rect 8280 1390 8360 1400
rect 9720 1390 9730 1400
rect 470 1380 840 1390
rect 990 1380 1020 1390
rect 2080 1380 2100 1390
rect 2990 1380 3030 1390
rect 4390 1380 4400 1390
rect 4500 1380 4780 1390
rect 4870 1380 4890 1390
rect 4900 1380 4920 1390
rect 4940 1380 4960 1390
rect 4970 1380 4980 1390
rect 4990 1380 5140 1390
rect 5150 1380 5160 1390
rect 5370 1380 5390 1390
rect 5520 1380 5540 1390
rect 5600 1380 5620 1390
rect 5890 1380 6200 1390
rect 6310 1380 6790 1390
rect 6800 1380 6810 1390
rect 7820 1380 7860 1390
rect 8290 1380 8320 1390
rect 8330 1380 8340 1390
rect 9260 1380 9270 1390
rect 9280 1380 9290 1390
rect 9950 1380 9990 1390
rect 470 1370 840 1380
rect 980 1370 1020 1380
rect 2080 1370 2110 1380
rect 2890 1370 2910 1380
rect 2970 1370 3020 1380
rect 4170 1370 4180 1380
rect 4460 1370 4480 1380
rect 4500 1370 4790 1380
rect 4810 1370 4820 1380
rect 4840 1370 4860 1380
rect 4870 1370 4920 1380
rect 4950 1370 4960 1380
rect 4970 1370 4980 1380
rect 4990 1370 5120 1380
rect 5150 1370 5160 1380
rect 5190 1370 5200 1380
rect 5270 1370 5280 1380
rect 5380 1370 5400 1380
rect 5610 1370 5620 1380
rect 5920 1370 6200 1380
rect 6310 1370 6790 1380
rect 7390 1370 7400 1380
rect 7830 1370 7860 1380
rect 8290 1370 8320 1380
rect 9250 1370 9260 1380
rect 9990 1370 9990 1380
rect 470 1360 840 1370
rect 960 1360 1020 1370
rect 2080 1360 2120 1370
rect 2860 1360 2900 1370
rect 2950 1360 3010 1370
rect 4430 1360 4480 1370
rect 4510 1360 4820 1370
rect 4840 1360 4860 1370
rect 4890 1360 4910 1370
rect 4920 1360 4930 1370
rect 4940 1360 4950 1370
rect 4970 1360 4980 1370
rect 4990 1360 5120 1370
rect 5250 1360 5260 1370
rect 5270 1360 5290 1370
rect 5410 1360 5420 1370
rect 5490 1360 5500 1370
rect 5600 1360 5610 1370
rect 5920 1360 6200 1370
rect 6310 1360 6790 1370
rect 7390 1360 7400 1370
rect 7830 1360 7860 1370
rect 8280 1360 8340 1370
rect 9690 1360 9700 1370
rect 9810 1360 9820 1370
rect 460 1350 840 1360
rect 940 1350 1020 1360
rect 2080 1350 2130 1360
rect 2850 1350 2910 1360
rect 2940 1350 2990 1360
rect 4400 1350 4410 1360
rect 4420 1350 4480 1360
rect 4510 1350 4820 1360
rect 4840 1350 4860 1360
rect 4870 1350 4920 1360
rect 4950 1350 4960 1360
rect 4970 1350 5110 1360
rect 5120 1350 5130 1360
rect 5180 1350 5220 1360
rect 5420 1350 5430 1360
rect 5500 1350 5510 1360
rect 5580 1350 5600 1360
rect 5930 1350 5950 1360
rect 5960 1350 6200 1360
rect 6310 1350 6790 1360
rect 7830 1350 7860 1360
rect 8270 1350 8340 1360
rect 9820 1350 9830 1360
rect 9960 1350 9970 1360
rect 460 1340 820 1350
rect 830 1340 840 1350
rect 940 1340 1020 1350
rect 2090 1340 2140 1350
rect 2840 1340 2980 1350
rect 4180 1340 4190 1350
rect 4410 1340 4490 1350
rect 4510 1340 4830 1350
rect 4850 1340 4940 1350
rect 4950 1340 4970 1350
rect 4980 1340 5080 1350
rect 5090 1340 5100 1350
rect 5140 1340 5210 1350
rect 5430 1340 5440 1350
rect 5520 1340 5540 1350
rect 5570 1340 5590 1350
rect 5930 1340 6200 1350
rect 6310 1340 6790 1350
rect 6810 1340 6820 1350
rect 7830 1340 7860 1350
rect 8280 1340 8310 1350
rect 9800 1340 9810 1350
rect 460 1330 840 1340
rect 930 1330 1020 1340
rect 2080 1330 2150 1340
rect 2820 1330 2970 1340
rect 4410 1330 4490 1340
rect 4510 1330 4970 1340
rect 4980 1330 5100 1340
rect 5200 1330 5210 1340
rect 5220 1330 5250 1340
rect 5380 1330 5390 1340
rect 5440 1330 5450 1340
rect 5530 1330 5570 1340
rect 5930 1330 6200 1340
rect 6310 1330 6800 1340
rect 6810 1330 6820 1340
rect 7830 1330 7860 1340
rect 9260 1330 9270 1340
rect 9640 1330 9650 1340
rect 9780 1330 9800 1340
rect 9830 1330 9840 1340
rect 450 1320 830 1330
rect 930 1320 1020 1330
rect 2080 1320 2150 1330
rect 2810 1320 2960 1330
rect 4410 1320 4490 1330
rect 4510 1320 4850 1330
rect 4860 1320 4940 1330
rect 4950 1320 4970 1330
rect 4990 1320 5070 1330
rect 5180 1320 5190 1330
rect 5200 1320 5240 1330
rect 5450 1320 5460 1330
rect 5930 1320 6200 1330
rect 6310 1320 6800 1330
rect 7830 1320 7860 1330
rect 9260 1320 9270 1330
rect 9640 1320 9650 1330
rect 9680 1320 9690 1330
rect 9710 1320 9720 1330
rect 9760 1320 9770 1330
rect 9830 1320 9840 1330
rect 450 1310 810 1320
rect 820 1310 830 1320
rect 920 1310 1020 1320
rect 2080 1310 2160 1320
rect 2790 1310 2930 1320
rect 3510 1310 3520 1320
rect 4190 1310 4200 1320
rect 4420 1310 4500 1320
rect 4510 1310 4970 1320
rect 4990 1310 5050 1320
rect 5120 1310 5140 1320
rect 5210 1310 5230 1320
rect 5240 1310 5250 1320
rect 5300 1310 5320 1320
rect 5440 1310 5450 1320
rect 5460 1310 5470 1320
rect 5930 1310 6200 1320
rect 6320 1310 6810 1320
rect 7840 1310 7860 1320
rect 9760 1310 9770 1320
rect 9830 1310 9840 1320
rect 450 1300 810 1310
rect 820 1300 830 1310
rect 920 1300 1020 1310
rect 2080 1300 2170 1310
rect 2790 1300 2920 1310
rect 4420 1300 4500 1310
rect 4520 1300 4970 1310
rect 4980 1300 5030 1310
rect 5110 1300 5160 1310
rect 5210 1300 5260 1310
rect 5300 1300 5310 1310
rect 5520 1300 5600 1310
rect 5920 1300 6200 1310
rect 6320 1300 6800 1310
rect 6810 1300 6820 1310
rect 7830 1300 7870 1310
rect 9700 1300 9710 1310
rect 9760 1300 9770 1310
rect 9780 1300 9800 1310
rect 9810 1300 9820 1310
rect 440 1290 820 1300
rect 920 1290 1010 1300
rect 2070 1290 2180 1300
rect 2760 1290 2910 1300
rect 4420 1290 4500 1300
rect 4520 1290 4940 1300
rect 4950 1290 4970 1300
rect 4980 1290 5010 1300
rect 5090 1290 5170 1300
rect 5370 1290 5450 1300
rect 5480 1290 5490 1300
rect 5510 1290 5550 1300
rect 5560 1290 5590 1300
rect 5920 1290 6210 1300
rect 6320 1290 6790 1300
rect 7400 1290 7410 1300
rect 7840 1290 7870 1300
rect 9760 1290 9770 1300
rect 9780 1290 9800 1300
rect 9990 1290 9990 1300
rect 440 1280 820 1290
rect 920 1280 1010 1290
rect 2040 1280 2190 1290
rect 2740 1280 2890 1290
rect 3500 1280 3510 1290
rect 4430 1280 4500 1290
rect 4520 1280 4930 1290
rect 4940 1280 4950 1290
rect 4990 1280 5000 1290
rect 5130 1280 5150 1290
rect 5200 1280 5300 1290
rect 5370 1280 5440 1290
rect 5670 1280 5690 1290
rect 5920 1280 6210 1290
rect 6310 1280 6790 1290
rect 7840 1280 7880 1290
rect 9260 1280 9270 1290
rect 9790 1280 9800 1290
rect 9820 1280 9830 1290
rect 9970 1280 9990 1290
rect 440 1270 820 1280
rect 920 1270 1010 1280
rect 2040 1270 2200 1280
rect 2720 1270 2880 1280
rect 4430 1270 4500 1280
rect 4520 1270 4930 1280
rect 4940 1270 4950 1280
rect 5120 1270 5160 1280
rect 5200 1270 5230 1280
rect 5250 1270 5290 1280
rect 5680 1270 5690 1280
rect 5930 1270 6210 1280
rect 6310 1270 6790 1280
rect 7400 1270 7410 1280
rect 7850 1270 7880 1280
rect 9130 1270 9140 1280
rect 9760 1270 9770 1280
rect 9820 1270 9830 1280
rect 9950 1270 9960 1280
rect 9980 1270 9990 1280
rect 430 1260 820 1270
rect 920 1260 1010 1270
rect 2040 1260 2200 1270
rect 2700 1260 2860 1270
rect 4430 1260 4510 1270
rect 4530 1260 4930 1270
rect 4940 1260 4960 1270
rect 5040 1260 5090 1270
rect 5120 1260 5170 1270
rect 5680 1260 5690 1270
rect 5930 1260 6210 1270
rect 6310 1260 6790 1270
rect 7850 1260 7880 1270
rect 9650 1260 9660 1270
rect 9740 1260 9750 1270
rect 9760 1260 9770 1270
rect 9960 1260 9970 1270
rect 430 1250 820 1260
rect 920 1250 1010 1260
rect 2040 1250 2210 1260
rect 2680 1250 2840 1260
rect 3500 1250 3510 1260
rect 4440 1250 4510 1260
rect 4530 1250 4930 1260
rect 4950 1250 5020 1260
rect 5070 1250 5130 1260
rect 5680 1250 5690 1260
rect 5920 1250 6220 1260
rect 6310 1250 6790 1260
rect 7850 1250 7880 1260
rect 9500 1250 9510 1260
rect 9670 1250 9680 1260
rect 9740 1250 9760 1260
rect 9990 1250 9990 1260
rect 430 1240 810 1250
rect 910 1240 1010 1250
rect 2030 1240 2200 1250
rect 2210 1240 2220 1250
rect 2650 1240 2820 1250
rect 4440 1240 4510 1250
rect 4530 1240 4940 1250
rect 5010 1240 5050 1250
rect 5680 1240 5690 1250
rect 5910 1240 5930 1250
rect 5940 1240 6230 1250
rect 6310 1240 6770 1250
rect 6790 1240 6800 1250
rect 7850 1240 7880 1250
rect 9280 1240 9290 1250
rect 9730 1240 9770 1250
rect 9820 1240 9830 1250
rect 420 1230 810 1240
rect 910 1230 1010 1240
rect 2030 1230 2250 1240
rect 2640 1230 2800 1240
rect 4200 1230 4210 1240
rect 4440 1230 4520 1240
rect 4530 1230 4760 1240
rect 4810 1230 4930 1240
rect 4950 1230 5000 1240
rect 5910 1230 5930 1240
rect 5940 1230 6230 1240
rect 6310 1230 6750 1240
rect 6790 1230 6800 1240
rect 7860 1230 7890 1240
rect 9500 1230 9510 1240
rect 9630 1230 9640 1240
rect 9660 1230 9670 1240
rect 9750 1230 9780 1240
rect 9960 1230 9970 1240
rect 420 1220 810 1230
rect 900 1220 1000 1230
rect 2030 1220 2270 1230
rect 2630 1220 2780 1230
rect 4440 1220 4520 1230
rect 4530 1220 4790 1230
rect 4870 1220 4910 1230
rect 5090 1220 5100 1230
rect 5910 1220 6240 1230
rect 6310 1220 6360 1230
rect 6370 1220 6740 1230
rect 7860 1220 7890 1230
rect 9520 1220 9530 1230
rect 9720 1220 9730 1230
rect 9760 1220 9800 1230
rect 9960 1220 9970 1230
rect 420 1210 790 1220
rect 800 1210 810 1220
rect 900 1210 1000 1220
rect 2020 1210 2140 1220
rect 2160 1210 2230 1220
rect 2240 1210 2300 1220
rect 2630 1210 2760 1220
rect 3800 1210 3810 1220
rect 4440 1210 4520 1220
rect 4540 1210 4680 1220
rect 4790 1210 4830 1220
rect 4840 1210 4850 1220
rect 4880 1210 4900 1220
rect 4950 1210 4970 1220
rect 4980 1210 4990 1220
rect 5080 1210 5100 1220
rect 5680 1210 5690 1220
rect 5890 1210 6240 1220
rect 6360 1210 6730 1220
rect 7860 1210 7890 1220
rect 9500 1210 9510 1220
rect 9620 1210 9630 1220
rect 9760 1210 9820 1220
rect 9960 1210 9970 1220
rect 410 1200 800 1210
rect 890 1200 980 1210
rect 990 1200 1000 1210
rect 2020 1200 2110 1210
rect 2180 1200 2190 1210
rect 2250 1200 2330 1210
rect 2600 1200 2610 1210
rect 2620 1200 2750 1210
rect 4450 1200 4520 1210
rect 4540 1200 4570 1210
rect 4700 1200 4760 1210
rect 4900 1200 4920 1210
rect 4930 1200 4980 1210
rect 5090 1200 5100 1210
rect 5170 1200 5180 1210
rect 5680 1200 5700 1210
rect 5910 1200 6250 1210
rect 6380 1200 6720 1210
rect 7410 1200 7420 1210
rect 7860 1200 7900 1210
rect 9140 1200 9150 1210
rect 9770 1200 9820 1210
rect 9960 1200 9970 1210
rect 410 1190 800 1200
rect 890 1190 980 1200
rect 2010 1190 2100 1200
rect 2250 1190 2420 1200
rect 2430 1190 2450 1200
rect 2490 1190 2500 1200
rect 2510 1190 2740 1200
rect 3830 1190 3840 1200
rect 4470 1190 4480 1200
rect 4610 1190 4710 1200
rect 4900 1190 4980 1200
rect 5090 1190 5100 1200
rect 5160 1190 5180 1200
rect 5680 1190 5690 1200
rect 5910 1190 6250 1200
rect 6390 1190 6700 1200
rect 6820 1190 6830 1200
rect 7410 1190 7420 1200
rect 7870 1190 7900 1200
rect 9610 1190 9620 1200
rect 9640 1190 9650 1200
rect 9770 1190 9780 1200
rect 9810 1190 9820 1200
rect 9940 1190 9990 1200
rect 410 1180 790 1190
rect 870 1180 960 1190
rect 2010 1180 2100 1190
rect 2250 1180 2730 1190
rect 4540 1180 4670 1190
rect 4690 1180 4700 1190
rect 4720 1180 4730 1190
rect 4900 1180 4980 1190
rect 5090 1180 5110 1190
rect 5170 1180 5180 1190
rect 5210 1180 5300 1190
rect 5880 1180 6250 1190
rect 6390 1180 6690 1190
rect 6800 1180 6810 1190
rect 6820 1180 6830 1190
rect 7870 1180 7900 1190
rect 9350 1180 9360 1190
rect 9500 1180 9510 1190
rect 9700 1180 9710 1190
rect 9760 1180 9780 1190
rect 9810 1180 9820 1190
rect 400 1170 790 1180
rect 870 1170 960 1180
rect 980 1170 990 1180
rect 2010 1170 2080 1180
rect 2270 1170 2740 1180
rect 2750 1170 2830 1180
rect 3550 1170 3560 1180
rect 4450 1170 4570 1180
rect 4580 1170 4590 1180
rect 4720 1170 4730 1180
rect 4900 1170 4980 1180
rect 5090 1170 5110 1180
rect 5130 1170 5330 1180
rect 5370 1170 5380 1180
rect 5680 1170 5700 1180
rect 5880 1170 6250 1180
rect 6370 1170 6670 1180
rect 6800 1170 6810 1180
rect 6820 1170 6830 1180
rect 7870 1170 7910 1180
rect 9630 1170 9640 1180
rect 9700 1170 9710 1180
rect 9760 1170 9770 1180
rect 400 1160 780 1170
rect 870 1160 990 1170
rect 2010 1160 2070 1170
rect 2280 1160 2850 1170
rect 3560 1160 3570 1170
rect 3870 1160 3880 1170
rect 4210 1160 4220 1170
rect 4460 1160 4560 1170
rect 4650 1160 4670 1170
rect 4720 1160 4730 1170
rect 4750 1160 4760 1170
rect 4910 1160 4980 1170
rect 5050 1160 5390 1170
rect 5420 1160 5430 1170
rect 5680 1160 5690 1170
rect 5880 1160 5890 1170
rect 5900 1160 6250 1170
rect 6380 1160 6660 1170
rect 6800 1160 6810 1170
rect 6820 1160 6830 1170
rect 7880 1160 7910 1170
rect 9360 1160 9370 1170
rect 9510 1160 9520 1170
rect 9700 1160 9710 1170
rect 9800 1160 9820 1170
rect 390 1150 640 1160
rect 660 1150 670 1160
rect 680 1150 780 1160
rect 870 1150 990 1160
rect 2010 1150 2070 1160
rect 2290 1150 2850 1160
rect 4460 1150 4560 1160
rect 4580 1150 4590 1160
rect 4650 1150 4670 1160
rect 4910 1150 5380 1160
rect 5420 1150 5430 1160
rect 5450 1150 5460 1160
rect 5680 1150 5690 1160
rect 5840 1150 5860 1160
rect 5920 1150 6250 1160
rect 6380 1150 6640 1160
rect 6820 1150 6830 1160
rect 7870 1150 7910 1160
rect 9150 1150 9160 1160
rect 9710 1150 9720 1160
rect 9820 1150 9830 1160
rect 390 1140 610 1150
rect 680 1140 760 1150
rect 880 1140 980 1150
rect 2010 1140 2050 1150
rect 2330 1140 2870 1150
rect 4460 1140 4560 1150
rect 4580 1140 4590 1150
rect 4660 1140 4670 1150
rect 4900 1140 5400 1150
rect 5430 1140 5440 1150
rect 5450 1140 5460 1150
rect 5620 1140 5670 1150
rect 5680 1140 5690 1150
rect 5890 1140 5900 1150
rect 5920 1140 6260 1150
rect 6380 1140 6630 1150
rect 6820 1140 6830 1150
rect 7880 1140 7910 1150
rect 9530 1140 9540 1150
rect 9610 1140 9620 1150
rect 9820 1140 9830 1150
rect 390 1130 620 1140
rect 750 1130 770 1140
rect 880 1130 990 1140
rect 2000 1130 2040 1140
rect 2330 1130 2880 1140
rect 3910 1130 3920 1140
rect 4460 1130 4560 1140
rect 4580 1130 4590 1140
rect 4650 1130 4670 1140
rect 4830 1130 5400 1140
rect 5680 1130 5690 1140
rect 5730 1130 5740 1140
rect 5900 1130 5910 1140
rect 5940 1130 6260 1140
rect 6410 1130 6610 1140
rect 7880 1130 7910 1140
rect 9340 1130 9350 1140
rect 9380 1130 9390 1140
rect 380 1120 630 1130
rect 760 1120 770 1130
rect 880 1120 990 1130
rect 2000 1120 2040 1130
rect 2350 1120 2890 1130
rect 4460 1120 4560 1130
rect 4660 1120 4670 1130
rect 4690 1120 4700 1130
rect 4710 1120 4720 1130
rect 4730 1120 5400 1130
rect 5680 1120 5690 1130
rect 5730 1120 5740 1130
rect 5900 1120 5910 1130
rect 5920 1120 5930 1130
rect 5940 1120 6260 1130
rect 6400 1120 6600 1130
rect 7880 1120 7910 1130
rect 9600 1120 9610 1130
rect 9720 1120 9730 1130
rect 380 1110 610 1120
rect 750 1110 770 1120
rect 880 1110 990 1120
rect 1990 1110 2030 1120
rect 2350 1110 2890 1120
rect 4470 1110 4560 1120
rect 4590 1110 4600 1120
rect 4610 1110 4620 1120
rect 4630 1110 5400 1120
rect 5410 1110 5440 1120
rect 5520 1110 5530 1120
rect 5620 1110 5630 1120
rect 5680 1110 5690 1120
rect 5800 1110 5810 1120
rect 5900 1110 6260 1120
rect 6400 1110 6580 1120
rect 7880 1110 7910 1120
rect 9360 1110 9370 1120
rect 9540 1110 9550 1120
rect 9600 1110 9610 1120
rect 9720 1110 9730 1120
rect 9810 1110 9820 1120
rect 380 1100 610 1110
rect 750 1100 760 1110
rect 870 1100 980 1110
rect 1600 1100 1610 1110
rect 1990 1100 2030 1110
rect 2380 1100 2650 1110
rect 2800 1100 2890 1110
rect 3620 1100 3630 1110
rect 4110 1100 4120 1110
rect 4470 1100 5440 1110
rect 5450 1100 5470 1110
rect 5480 1100 5500 1110
rect 5660 1100 5670 1110
rect 5680 1100 5690 1110
rect 5720 1100 5820 1110
rect 5830 1100 5890 1110
rect 5900 1100 6270 1110
rect 6400 1100 6560 1110
rect 6810 1100 6820 1110
rect 7880 1100 7910 1110
rect 9390 1100 9400 1110
rect 9540 1100 9550 1110
rect 9590 1100 9600 1110
rect 9720 1100 9730 1110
rect 9820 1100 9830 1110
rect 9880 1100 9900 1110
rect 370 1090 620 1100
rect 750 1090 760 1100
rect 870 1090 980 1100
rect 1540 1090 1550 1100
rect 1990 1090 2020 1100
rect 2400 1090 2410 1100
rect 2420 1090 2500 1100
rect 2520 1090 2530 1100
rect 2810 1090 2890 1100
rect 3630 1090 3640 1100
rect 3970 1090 3980 1100
rect 4100 1090 4130 1100
rect 4480 1090 5470 1100
rect 5650 1090 5700 1100
rect 5720 1090 5890 1100
rect 5910 1090 6270 1100
rect 6420 1090 6540 1100
rect 7880 1090 7910 1100
rect 9230 1090 9240 1100
rect 9360 1090 9370 1100
rect 9580 1090 9590 1100
rect 9720 1090 9730 1100
rect 9820 1090 9830 1100
rect 9870 1090 9920 1100
rect 370 1080 620 1090
rect 870 1080 980 1090
rect 1990 1080 2020 1090
rect 2820 1080 2900 1090
rect 4090 1080 4110 1090
rect 4220 1080 4230 1090
rect 4480 1080 5220 1090
rect 5230 1080 5480 1090
rect 5520 1080 5530 1090
rect 5590 1080 5600 1090
rect 5650 1080 5690 1090
rect 5700 1080 5870 1090
rect 5950 1080 6270 1090
rect 6430 1080 6520 1090
rect 6810 1080 6820 1090
rect 7420 1080 7430 1090
rect 7890 1080 7910 1090
rect 9290 1080 9300 1090
rect 9570 1080 9580 1090
rect 9720 1080 9730 1090
rect 9880 1080 9920 1090
rect 9940 1080 9960 1090
rect 9970 1080 9980 1090
rect 360 1070 620 1080
rect 860 1070 980 1080
rect 1510 1070 1520 1080
rect 1640 1070 1650 1080
rect 1980 1070 2020 1080
rect 2840 1070 2910 1080
rect 4010 1070 4020 1080
rect 4100 1070 4110 1080
rect 4220 1070 4230 1080
rect 4480 1070 5200 1080
rect 5210 1070 5440 1080
rect 5450 1070 5470 1080
rect 5490 1070 5520 1080
rect 5590 1070 5670 1080
rect 5710 1070 5850 1080
rect 5870 1070 5880 1080
rect 5990 1070 6010 1080
rect 6030 1070 6270 1080
rect 6460 1070 6470 1080
rect 6480 1070 6500 1080
rect 6810 1070 6820 1080
rect 7420 1070 7430 1080
rect 7890 1070 7920 1080
rect 9560 1070 9580 1080
rect 9720 1070 9730 1080
rect 9850 1070 9860 1080
rect 9880 1070 9890 1080
rect 9990 1070 9990 1080
rect 360 1060 630 1070
rect 740 1060 750 1070
rect 860 1060 980 1070
rect 1980 1060 2020 1070
rect 2840 1060 2900 1070
rect 4020 1060 4030 1070
rect 4070 1060 4080 1070
rect 4100 1060 4130 1070
rect 4480 1060 5440 1070
rect 5450 1060 5470 1070
rect 5480 1060 5510 1070
rect 5520 1060 5560 1070
rect 5570 1060 5600 1070
rect 5620 1060 5670 1070
rect 5680 1060 5690 1070
rect 5710 1060 5800 1070
rect 5810 1060 5840 1070
rect 5850 1060 5890 1070
rect 5910 1060 5920 1070
rect 5960 1060 6270 1070
rect 6450 1060 6480 1070
rect 6810 1060 6820 1070
rect 7420 1060 7430 1070
rect 7900 1060 7920 1070
rect 9070 1060 9080 1070
rect 9360 1060 9370 1070
rect 9560 1060 9570 1070
rect 9840 1060 9850 1070
rect 9990 1060 9990 1070
rect 350 1050 630 1060
rect 740 1050 750 1060
rect 860 1050 970 1060
rect 1990 1050 2020 1060
rect 2840 1050 2900 1060
rect 4070 1050 4080 1060
rect 4090 1050 4130 1060
rect 4220 1050 4230 1060
rect 4480 1050 5370 1060
rect 5380 1050 5510 1060
rect 5520 1050 5600 1060
rect 5610 1050 5630 1060
rect 5640 1050 5670 1060
rect 5680 1050 5690 1060
rect 5700 1050 5770 1060
rect 5790 1050 5830 1060
rect 5850 1050 5860 1060
rect 5880 1050 5930 1060
rect 5960 1050 6280 1060
rect 6440 1050 6460 1060
rect 6810 1050 6820 1060
rect 7420 1050 7430 1060
rect 7900 1050 7920 1060
rect 9070 1050 9080 1060
rect 9130 1050 9140 1060
rect 9300 1050 9310 1060
rect 9530 1050 9540 1060
rect 9550 1050 9570 1060
rect 9800 1050 9820 1060
rect 9950 1050 9970 1060
rect 9980 1050 9990 1060
rect 350 1040 630 1050
rect 860 1040 970 1050
rect 1650 1040 1660 1050
rect 1980 1040 2010 1050
rect 2840 1040 2900 1050
rect 3680 1040 3690 1050
rect 4060 1040 4080 1050
rect 4110 1040 4120 1050
rect 4200 1040 4220 1050
rect 4570 1040 5470 1050
rect 5500 1040 5630 1050
rect 5640 1040 5670 1050
rect 5680 1040 5690 1050
rect 5720 1040 5770 1050
rect 5780 1040 5820 1050
rect 5880 1040 5940 1050
rect 5950 1040 6280 1050
rect 6410 1040 6440 1050
rect 6810 1040 6820 1050
rect 7420 1040 7430 1050
rect 7900 1040 7920 1050
rect 8170 1040 8180 1050
rect 9120 1040 9130 1050
rect 9300 1040 9310 1050
rect 9720 1040 9730 1050
rect 9820 1040 9830 1050
rect 9910 1040 9930 1050
rect 9950 1040 9970 1050
rect 9990 1040 9990 1050
rect 340 1030 630 1040
rect 730 1030 740 1040
rect 850 1030 970 1040
rect 1980 1030 2010 1040
rect 2840 1030 2900 1040
rect 3690 1030 3700 1040
rect 4200 1030 4210 1040
rect 4600 1030 5420 1040
rect 5430 1030 5490 1040
rect 5510 1030 5520 1040
rect 5550 1030 5590 1040
rect 5600 1030 5670 1040
rect 5680 1030 5690 1040
rect 5710 1030 5820 1040
rect 5840 1030 5860 1040
rect 5880 1030 6290 1040
rect 6400 1030 6430 1040
rect 6810 1030 6820 1040
rect 7900 1030 7920 1040
rect 8160 1030 8180 1040
rect 9290 1030 9310 1040
rect 9420 1030 9430 1040
rect 9520 1030 9530 1040
rect 9730 1030 9740 1040
rect 9820 1030 9830 1040
rect 9950 1030 9970 1040
rect 340 1020 650 1030
rect 730 1020 740 1030
rect 840 1020 960 1030
rect 1610 1020 1640 1030
rect 1980 1020 2010 1030
rect 2840 1020 2900 1030
rect 4080 1020 4090 1030
rect 4200 1020 4210 1030
rect 4630 1020 5490 1030
rect 5550 1020 5570 1030
rect 5610 1020 5620 1030
rect 5640 1020 5670 1030
rect 5680 1020 5690 1030
rect 5710 1020 5790 1030
rect 5810 1020 5980 1030
rect 6000 1020 6290 1030
rect 6370 1020 6410 1030
rect 6810 1020 6820 1030
rect 7910 1020 7930 1030
rect 8150 1020 8180 1030
rect 9060 1020 9070 1030
rect 9530 1020 9550 1030
rect 9730 1020 9740 1030
rect 9950 1020 9960 1030
rect 330 1010 670 1020
rect 840 1010 960 1020
rect 1600 1010 1650 1020
rect 1980 1010 2000 1020
rect 2840 1010 2900 1020
rect 4100 1010 4110 1020
rect 4210 1010 4220 1020
rect 4660 1010 5490 1020
rect 5530 1010 5570 1020
rect 5590 1010 5600 1020
rect 5640 1010 5680 1020
rect 5710 1010 5840 1020
rect 5850 1010 5980 1020
rect 5990 1010 6290 1020
rect 6360 1010 6400 1020
rect 6810 1010 6820 1020
rect 7900 1010 7930 1020
rect 8150 1010 8180 1020
rect 9000 1010 9020 1020
rect 9050 1010 9070 1020
rect 9120 1010 9130 1020
rect 9530 1010 9540 1020
rect 9790 1010 9810 1020
rect 9820 1010 9830 1020
rect 330 1000 670 1010
rect 680 1000 690 1010
rect 720 1000 730 1010
rect 830 1000 960 1010
rect 1580 1000 1650 1010
rect 1980 1000 2000 1010
rect 2840 1000 2890 1010
rect 4190 1000 4200 1010
rect 4690 1000 5380 1010
rect 5390 1000 5470 1010
rect 5530 1000 5620 1010
rect 5630 1000 5670 1010
rect 5710 1000 5850 1010
rect 5860 1000 6280 1010
rect 6290 1000 6300 1010
rect 6360 1000 6410 1010
rect 6810 1000 6820 1010
rect 7900 1000 7930 1010
rect 8150 1000 8190 1010
rect 8990 1000 9030 1010
rect 9050 1000 9070 1010
rect 9120 1000 9130 1010
rect 9420 1000 9430 1010
rect 9520 1000 9540 1010
rect 9780 1000 9810 1010
rect 9820 1000 9830 1010
rect 320 990 680 1000
rect 720 990 730 1000
rect 820 990 960 1000
rect 1560 990 1640 1000
rect 1980 990 2000 1000
rect 2820 990 2830 1000
rect 2840 990 2890 1000
rect 4170 990 4180 1000
rect 4200 990 4210 1000
rect 4710 990 5400 1000
rect 5420 990 5450 1000
rect 5520 990 5580 1000
rect 5610 990 5670 1000
rect 5680 990 5690 1000
rect 5710 990 5870 1000
rect 5890 990 5900 1000
rect 5910 990 5920 1000
rect 5930 990 6000 1000
rect 6010 990 6300 1000
rect 6350 990 6410 1000
rect 6820 990 6830 1000
rect 7910 990 7930 1000
rect 8150 990 8180 1000
rect 8970 990 9030 1000
rect 9040 990 9080 1000
rect 9120 990 9130 1000
rect 9140 990 9150 1000
rect 9520 990 9530 1000
rect 9770 990 9810 1000
rect 9820 990 9830 1000
rect 320 980 680 990
rect 690 980 700 990
rect 820 980 950 990
rect 1550 980 1630 990
rect 1980 980 2000 990
rect 2830 980 2890 990
rect 4160 980 4170 990
rect 4740 980 5400 990
rect 5430 980 5450 990
rect 5490 980 5580 990
rect 5640 980 5670 990
rect 5680 980 5690 990
rect 5720 980 5730 990
rect 5740 980 5870 990
rect 5890 980 5900 990
rect 5920 980 6290 990
rect 6350 980 6400 990
rect 6820 980 6830 990
rect 7920 980 7940 990
rect 8150 980 8180 990
rect 8960 980 9020 990
rect 9040 980 9080 990
rect 9120 980 9130 990
rect 9490 980 9500 990
rect 9510 980 9530 990
rect 9760 980 9770 990
rect 9780 980 9790 990
rect 310 970 700 980
rect 710 970 720 980
rect 820 970 950 980
rect 1400 970 1410 980
rect 1540 970 1610 980
rect 1980 970 2000 980
rect 2820 970 2880 980
rect 4760 970 5400 980
rect 5470 970 5520 980
rect 5530 970 5560 980
rect 5720 970 5730 980
rect 5760 970 5850 980
rect 5860 970 5870 980
rect 5920 970 6280 980
rect 6290 970 6300 980
rect 6350 970 6400 980
rect 6820 970 6840 980
rect 7920 970 7940 980
rect 8150 970 8190 980
rect 8950 970 9080 980
rect 9120 970 9130 980
rect 9500 970 9520 980
rect 9760 970 9770 980
rect 9820 970 9830 980
rect 310 960 710 970
rect 810 960 950 970
rect 1390 960 1400 970
rect 1520 960 1600 970
rect 1980 960 2000 970
rect 2820 960 2870 970
rect 4770 960 5030 970
rect 5040 960 5210 970
rect 5220 960 5300 970
rect 5320 960 5330 970
rect 5380 960 5390 970
rect 5540 960 5550 970
rect 5690 960 5700 970
rect 5880 960 5990 970
rect 6000 960 6270 970
rect 6350 960 6410 970
rect 6820 960 6840 970
rect 7920 960 7940 970
rect 8150 960 8190 970
rect 8950 960 9070 970
rect 9120 960 9130 970
rect 9140 960 9160 970
rect 9510 960 9520 970
rect 9760 960 9770 970
rect 300 950 710 960
rect 810 950 940 960
rect 1520 950 1590 960
rect 1980 950 2000 960
rect 2820 950 2850 960
rect 4790 950 4820 960
rect 4860 950 4900 960
rect 5090 950 5220 960
rect 5230 950 5300 960
rect 5320 950 5330 960
rect 5680 950 5700 960
rect 5840 950 5850 960
rect 5880 950 5890 960
rect 5970 950 6020 960
rect 6040 950 6270 960
rect 6360 950 6410 960
rect 6820 950 6840 960
rect 7920 950 7940 960
rect 8140 950 8190 960
rect 8940 950 9070 960
rect 9140 950 9160 960
rect 9250 950 9260 960
rect 9510 950 9520 960
rect 300 940 710 950
rect 810 940 930 950
rect 1360 940 1370 950
rect 1510 940 1590 950
rect 1980 940 2000 950
rect 2810 940 2850 950
rect 4840 940 4850 950
rect 5140 940 5240 950
rect 5290 940 5310 950
rect 5320 940 5330 950
rect 5350 940 5360 950
rect 5590 940 5600 950
rect 5690 940 5700 950
rect 5870 940 5890 950
rect 5960 940 6030 950
rect 6040 940 6230 950
rect 6240 940 6250 950
rect 6360 940 6410 950
rect 6820 940 6840 950
rect 7920 940 7940 950
rect 8140 940 8190 950
rect 8940 940 9070 950
rect 290 930 700 940
rect 810 930 940 940
rect 1350 930 1360 940
rect 1500 930 1570 940
rect 1980 930 2000 940
rect 2790 930 2840 940
rect 3790 930 3800 940
rect 5010 930 5020 940
rect 5190 930 5250 940
rect 5270 930 5330 940
rect 5350 930 5370 940
rect 5590 930 5600 940
rect 5860 930 5870 940
rect 6020 930 6220 940
rect 6370 930 6420 940
rect 7920 930 7950 940
rect 8140 930 8200 940
rect 8930 930 9070 940
rect 9160 930 9170 940
rect 9210 930 9220 940
rect 9250 930 9260 940
rect 9490 930 9500 940
rect 280 920 700 930
rect 810 920 940 930
rect 1480 920 1570 930
rect 1990 920 2000 930
rect 2790 920 2820 930
rect 4910 920 4920 930
rect 4950 920 5080 930
rect 5210 920 5330 930
rect 5350 920 5360 930
rect 5580 920 5600 930
rect 5690 920 5700 930
rect 5860 920 5870 930
rect 6020 920 6220 930
rect 6370 920 6420 930
rect 7920 920 7950 930
rect 8150 920 8200 930
rect 8930 920 9080 930
rect 280 910 690 920
rect 810 910 940 920
rect 1470 910 1560 920
rect 1990 910 2000 920
rect 2770 910 2800 920
rect 4870 910 5130 920
rect 5250 910 5330 920
rect 5490 910 5500 920
rect 5590 910 5600 920
rect 5670 910 5700 920
rect 5850 910 5860 920
rect 6020 910 6030 920
rect 6040 910 6220 920
rect 6290 910 6300 920
rect 6380 910 6420 920
rect 6830 910 6840 920
rect 7420 910 7430 920
rect 7930 910 7960 920
rect 8150 910 8200 920
rect 8910 910 9080 920
rect 9480 910 9490 920
rect 270 900 690 910
rect 810 900 930 910
rect 1310 900 1320 910
rect 1450 900 1550 910
rect 1990 900 2000 910
rect 2760 900 2780 910
rect 4870 900 4920 910
rect 5000 900 5170 910
rect 5250 900 5270 910
rect 5300 900 5330 910
rect 5400 900 5410 910
rect 5770 900 5780 910
rect 5790 900 5810 910
rect 5850 900 5860 910
rect 6040 900 6230 910
rect 6370 900 6420 910
rect 7930 900 7960 910
rect 8150 900 8200 910
rect 8900 900 9090 910
rect 9470 900 9480 910
rect 260 890 690 900
rect 810 890 840 900
rect 880 890 890 900
rect 910 890 940 900
rect 1300 890 1310 900
rect 1440 890 1540 900
rect 1990 890 2000 900
rect 2750 890 2770 900
rect 4850 890 4880 900
rect 5080 890 5180 900
rect 5280 890 5290 900
rect 5300 890 5330 900
rect 5400 890 5410 900
rect 5680 890 5690 900
rect 5750 890 5780 900
rect 5790 890 5810 900
rect 5910 890 5930 900
rect 6000 890 6010 900
rect 6040 890 6220 900
rect 6370 890 6410 900
rect 6830 890 6840 900
rect 7420 890 7430 900
rect 7930 890 7960 900
rect 8150 890 8210 900
rect 8890 890 9080 900
rect 9440 890 9450 900
rect 9470 890 9480 900
rect 260 880 680 890
rect 920 880 930 890
rect 1420 880 1530 890
rect 2000 880 2010 890
rect 2730 880 2750 890
rect 5110 880 5180 890
rect 5290 880 5330 890
rect 5570 880 5580 890
rect 5680 880 5690 890
rect 5730 880 5810 890
rect 5970 880 5980 890
rect 6050 880 6220 890
rect 6280 880 6290 890
rect 6380 880 6420 890
rect 7420 880 7430 890
rect 7930 880 7960 890
rect 8150 880 8210 890
rect 8870 880 9070 890
rect 9170 880 9180 890
rect 9470 880 9480 890
rect 250 870 680 880
rect 920 870 930 880
rect 1410 870 1520 880
rect 2000 870 2010 880
rect 2720 870 2730 880
rect 3840 870 3850 880
rect 5170 870 5190 880
rect 5300 870 5340 880
rect 5520 870 5540 880
rect 5570 870 5600 880
rect 5630 870 5660 880
rect 5680 870 5690 880
rect 5710 870 5790 880
rect 5800 870 5810 880
rect 6010 870 6020 880
rect 6050 870 6210 880
rect 6380 870 6420 880
rect 7930 870 7960 880
rect 8150 870 8200 880
rect 8870 870 9070 880
rect 240 860 670 870
rect 920 860 930 870
rect 1260 860 1270 870
rect 1410 860 1500 870
rect 2000 860 2010 870
rect 2700 860 2710 870
rect 3850 860 3860 870
rect 5190 860 5220 870
rect 5240 860 5260 870
rect 5320 860 5350 870
rect 5430 860 5670 870
rect 5680 860 5690 870
rect 5710 860 5820 870
rect 5960 860 5970 870
rect 6010 860 6020 870
rect 6030 860 6220 870
rect 6390 860 6420 870
rect 7420 860 7430 870
rect 7930 860 7960 870
rect 8150 860 8200 870
rect 8870 860 9070 870
rect 9110 860 9120 870
rect 9420 860 9430 870
rect 240 850 670 860
rect 910 850 930 860
rect 1410 850 1490 860
rect 2010 850 2020 860
rect 2680 850 2690 860
rect 3860 850 3870 860
rect 4570 850 4590 860
rect 4870 850 4880 860
rect 4960 850 4970 860
rect 4980 850 4990 860
rect 5070 850 5080 860
rect 5210 850 5270 860
rect 5340 850 5370 860
rect 5440 850 5670 860
rect 5710 850 5820 860
rect 5960 850 5980 860
rect 6030 850 6220 860
rect 6280 850 6290 860
rect 6390 850 6440 860
rect 7420 850 7430 860
rect 7930 850 7950 860
rect 8150 850 8210 860
rect 8860 850 9080 860
rect 9110 850 9120 860
rect 9450 850 9460 860
rect 230 840 670 850
rect 910 840 930 850
rect 1400 840 1490 850
rect 2010 840 2020 850
rect 2660 840 2670 850
rect 3870 840 3880 850
rect 4570 840 4590 850
rect 5010 840 5030 850
rect 5060 840 5080 850
rect 5220 840 5280 850
rect 5350 840 5370 850
rect 5410 840 5470 850
rect 5490 840 5610 850
rect 5710 840 5770 850
rect 5780 840 5790 850
rect 5820 840 5830 850
rect 5840 840 5860 850
rect 5880 840 5890 850
rect 5920 840 5950 850
rect 6010 840 6210 850
rect 6280 840 6290 850
rect 6400 840 6440 850
rect 7420 840 7430 850
rect 7940 840 7960 850
rect 8150 840 8220 850
rect 8860 840 9080 850
rect 9110 840 9120 850
rect 9410 840 9420 850
rect 220 830 670 840
rect 910 830 920 840
rect 1220 830 1230 840
rect 1400 830 1470 840
rect 2020 830 2030 840
rect 2640 830 2650 840
rect 3880 830 3890 840
rect 5010 830 5040 840
rect 5230 830 5250 840
rect 5270 830 5290 840
rect 5360 830 5380 840
rect 5430 830 5460 840
rect 5520 830 5530 840
rect 5570 830 5610 840
rect 5630 830 5670 840
rect 5680 830 5690 840
rect 5710 830 5760 840
rect 5880 830 5890 840
rect 6000 830 6150 840
rect 6160 830 6200 840
rect 6280 830 6290 840
rect 6410 830 6450 840
rect 7420 830 7430 840
rect 7940 830 7960 840
rect 8140 830 8220 840
rect 8850 830 9080 840
rect 9110 830 9120 840
rect 9430 830 9440 840
rect 210 820 660 830
rect 880 820 920 830
rect 1390 820 1470 830
rect 2020 820 2030 830
rect 2620 820 2630 830
rect 4920 820 4930 830
rect 5130 820 5150 830
rect 5170 820 5180 830
rect 5240 820 5270 830
rect 5280 820 5310 830
rect 5370 820 5380 830
rect 5400 820 5420 830
rect 5430 820 5470 830
rect 5480 820 5490 830
rect 5510 820 5560 830
rect 5590 820 5600 830
rect 5680 820 5690 830
rect 5710 820 5770 830
rect 5880 820 5890 830
rect 6020 820 6190 830
rect 6410 820 6450 830
rect 7410 820 7430 830
rect 7940 820 7960 830
rect 8140 820 8220 830
rect 8850 820 9080 830
rect 9110 820 9120 830
rect 9190 820 9200 830
rect 9430 820 9440 830
rect 200 810 660 820
rect 860 810 920 820
rect 1380 810 1470 820
rect 2020 810 2040 820
rect 2600 810 2610 820
rect 5140 810 5150 820
rect 5160 810 5170 820
rect 5190 810 5200 820
rect 5250 810 5260 820
rect 5270 810 5280 820
rect 5300 810 5320 820
rect 5360 810 5370 820
rect 5380 810 5390 820
rect 5420 810 5670 820
rect 5680 810 5690 820
rect 5700 810 5770 820
rect 5880 810 5900 820
rect 6050 810 6190 820
rect 6290 810 6300 820
rect 6410 810 6460 820
rect 7420 810 7430 820
rect 7940 810 7970 820
rect 8140 810 8230 820
rect 8840 810 9080 820
rect 9110 810 9120 820
rect 9420 810 9430 820
rect 190 800 660 810
rect 850 800 920 810
rect 1180 800 1190 810
rect 1360 800 1480 810
rect 2030 800 2040 810
rect 2580 800 2590 810
rect 4300 800 4310 810
rect 5090 800 5120 810
rect 5170 800 5240 810
rect 5250 800 5300 810
rect 5310 800 5320 810
rect 5390 800 5400 810
rect 5420 800 5440 810
rect 5460 800 5470 810
rect 5490 800 5530 810
rect 5550 800 5670 810
rect 5680 800 5690 810
rect 5700 800 5780 810
rect 5790 800 5850 810
rect 6040 800 6190 810
rect 6290 800 6300 810
rect 6410 800 6460 810
rect 7420 800 7430 810
rect 7940 800 7970 810
rect 8140 800 8230 810
rect 8830 800 9090 810
rect 9100 800 9110 810
rect 9420 800 9430 810
rect 180 790 650 800
rect 830 790 920 800
rect 1340 790 1480 800
rect 2030 790 2040 800
rect 2560 790 2570 800
rect 3930 790 3940 800
rect 5210 790 5220 800
rect 5240 790 5250 800
rect 5270 790 5310 800
rect 5320 790 5350 800
rect 5400 790 5410 800
rect 5430 790 5450 800
rect 5550 790 5690 800
rect 5710 790 5780 800
rect 5790 790 5800 800
rect 5810 790 5820 800
rect 6040 790 6060 800
rect 6070 790 6150 800
rect 6160 790 6190 800
rect 6290 790 6300 800
rect 6420 790 6460 800
rect 6850 790 6860 800
rect 7410 790 7430 800
rect 7950 790 7970 800
rect 8140 790 8230 800
rect 8830 790 9090 800
rect 9100 790 9110 800
rect 9420 790 9430 800
rect 170 780 650 790
rect 820 780 910 790
rect 1150 780 1160 790
rect 1320 780 1470 790
rect 3660 780 3680 790
rect 4320 780 4330 790
rect 5310 780 5320 790
rect 5330 780 5350 790
rect 5400 780 5490 790
rect 5520 780 5690 790
rect 5700 780 5790 790
rect 5970 780 5980 790
rect 6060 780 6080 790
rect 6090 780 6160 790
rect 6290 780 6310 790
rect 6420 780 6460 790
rect 6850 780 6860 790
rect 7410 780 7430 790
rect 7950 780 7970 790
rect 8140 780 8150 790
rect 8160 780 8230 790
rect 8830 780 9090 790
rect 9100 780 9110 790
rect 9410 780 9420 790
rect 160 770 650 780
rect 800 770 910 780
rect 1310 770 1460 780
rect 3660 770 3670 780
rect 3730 770 3740 780
rect 3970 770 3980 780
rect 4330 770 4340 780
rect 5320 770 5360 780
rect 5410 770 5420 780
rect 5440 770 5490 780
rect 5520 770 5690 780
rect 5700 770 5770 780
rect 5870 770 5880 780
rect 5960 770 5970 780
rect 6090 770 6110 780
rect 6120 770 6180 780
rect 6290 770 6310 780
rect 6410 770 6470 780
rect 6850 770 6860 780
rect 7420 770 7430 780
rect 7950 770 7980 780
rect 8140 770 8150 780
rect 8160 770 8240 780
rect 8810 770 9090 780
rect 9100 770 9110 780
rect 9200 770 9210 780
rect 150 760 640 770
rect 780 760 900 770
rect 1280 760 1450 770
rect 3570 760 3590 770
rect 3650 760 3670 770
rect 4330 760 4350 770
rect 4910 760 4920 770
rect 5270 760 5280 770
rect 5330 760 5350 770
rect 5420 760 5430 770
rect 5440 760 5490 770
rect 5520 760 5690 770
rect 5710 760 5770 770
rect 6040 760 6050 770
rect 6160 760 6170 770
rect 6300 760 6310 770
rect 6420 760 6480 770
rect 6850 760 6860 770
rect 7400 760 7430 770
rect 7950 760 7980 770
rect 8140 760 8150 770
rect 8160 760 8250 770
rect 8800 760 9080 770
rect 9100 760 9110 770
rect 9400 760 9410 770
rect 140 750 640 760
rect 770 750 900 760
rect 1110 750 1120 760
rect 1290 750 1440 760
rect 2050 750 2060 760
rect 2490 750 2500 760
rect 3530 750 3540 760
rect 5170 750 5190 760
rect 5280 750 5300 760
rect 5340 750 5360 760
rect 5430 750 5450 760
rect 5460 750 5510 760
rect 5530 750 5690 760
rect 5700 750 5770 760
rect 6290 750 6320 760
rect 6430 750 6490 760
rect 6850 750 6860 760
rect 7400 750 7430 760
rect 7960 750 7980 760
rect 8140 750 8150 760
rect 8160 750 8250 760
rect 8790 750 9090 760
rect 130 740 640 750
rect 760 740 900 750
rect 1290 740 1420 750
rect 2060 740 2070 750
rect 3450 740 3520 750
rect 5290 740 5320 750
rect 5350 740 5360 750
rect 5440 740 5550 750
rect 5560 740 5570 750
rect 5580 740 5690 750
rect 5700 740 5770 750
rect 6300 740 6320 750
rect 6430 740 6490 750
rect 6850 740 6860 750
rect 7400 740 7430 750
rect 7960 740 7980 750
rect 8140 740 8150 750
rect 8160 740 8250 750
rect 8780 740 9080 750
rect 9100 740 9110 750
rect 120 730 630 740
rect 750 730 890 740
rect 1290 730 1410 740
rect 2060 730 2070 740
rect 2460 730 2470 740
rect 3420 730 3430 740
rect 4000 730 4010 740
rect 5360 730 5380 740
rect 5450 730 5510 740
rect 5520 730 5690 740
rect 5700 730 5740 740
rect 5750 730 5760 740
rect 5850 730 5860 740
rect 6020 730 6040 740
rect 6110 730 6120 740
rect 6300 730 6320 740
rect 6430 730 6490 740
rect 6850 730 6860 740
rect 7400 730 7430 740
rect 7970 730 7980 740
rect 8140 730 8240 740
rect 8770 730 9080 740
rect 9100 730 9110 740
rect 9210 730 9220 740
rect 110 720 630 730
rect 750 720 900 730
rect 1290 720 1410 730
rect 4010 720 4020 730
rect 5150 720 5170 730
rect 5180 720 5200 730
rect 5460 720 5500 730
rect 5520 720 5640 730
rect 5650 720 5690 730
rect 5700 720 5740 730
rect 5760 720 5770 730
rect 5810 720 5820 730
rect 5830 720 5840 730
rect 5980 720 6010 730
rect 6050 720 6060 730
rect 6290 720 6330 730
rect 6440 720 6490 730
rect 6850 720 6870 730
rect 7410 720 7430 730
rect 7970 720 7990 730
rect 8140 720 8230 730
rect 8780 720 9080 730
rect 9100 720 9110 730
rect 9120 720 9140 730
rect 90 710 630 720
rect 740 710 890 720
rect 1300 710 1400 720
rect 2070 710 2080 720
rect 3380 710 3390 720
rect 5050 710 5060 720
rect 5130 710 5190 720
rect 5370 710 5380 720
rect 5470 710 5490 720
rect 5500 710 5690 720
rect 5700 710 5780 720
rect 5970 710 6000 720
rect 6290 710 6330 720
rect 6460 710 6490 720
rect 6860 710 6870 720
rect 7400 710 7430 720
rect 7970 710 7990 720
rect 8140 710 8250 720
rect 8770 710 9080 720
rect 9110 710 9120 720
rect 80 700 620 710
rect 730 700 910 710
rect 1040 700 1050 710
rect 1300 700 1390 710
rect 2410 700 2420 710
rect 3360 700 3370 710
rect 4010 700 4020 710
rect 4920 700 4930 710
rect 5050 700 5060 710
rect 5140 700 5200 710
rect 5250 700 5260 710
rect 5350 700 5360 710
rect 5380 700 5400 710
rect 5480 700 5490 710
rect 5500 700 5510 710
rect 5520 700 5670 710
rect 5680 700 5690 710
rect 5700 700 5780 710
rect 5880 700 5890 710
rect 5940 700 5950 710
rect 6290 700 6330 710
rect 6460 700 6510 710
rect 6860 700 6870 710
rect 7400 700 7430 710
rect 7980 700 7990 710
rect 8140 700 8260 710
rect 8770 700 9080 710
rect 60 690 620 700
rect 730 690 910 700
rect 1300 690 1380 700
rect 2390 690 2400 700
rect 4770 690 4780 700
rect 4920 690 4930 700
rect 5140 690 5200 700
rect 5390 690 5410 700
rect 5490 690 5500 700
rect 5530 690 5580 700
rect 5590 690 5620 700
rect 5630 690 5650 700
rect 5660 690 5690 700
rect 5700 690 5770 700
rect 5780 690 5810 700
rect 5820 690 5840 700
rect 5990 690 6000 700
rect 6160 690 6170 700
rect 6290 690 6330 700
rect 6460 690 6520 700
rect 6860 690 6880 700
rect 7400 690 7420 700
rect 7980 690 8000 700
rect 8140 690 8260 700
rect 8750 690 9100 700
rect 9110 690 9120 700
rect 50 680 610 690
rect 720 680 920 690
rect 1010 680 1020 690
rect 1300 680 1360 690
rect 3330 680 3340 690
rect 4720 680 4770 690
rect 4920 680 4930 690
rect 5140 680 5210 690
rect 5400 680 5410 690
rect 5490 680 5500 690
rect 5540 680 5550 690
rect 5560 680 5580 690
rect 5610 680 5620 690
rect 5650 680 5690 690
rect 5700 680 5780 690
rect 5800 680 5810 690
rect 6290 680 6340 690
rect 6460 680 6520 690
rect 6860 680 6880 690
rect 7390 680 7420 690
rect 7980 680 8010 690
rect 8140 680 8280 690
rect 8750 680 9090 690
rect 9100 680 9110 690
rect 9350 680 9360 690
rect 30 670 610 680
rect 730 670 920 680
rect 1000 670 1010 680
rect 1300 670 1360 680
rect 2090 670 2100 680
rect 2360 670 2370 680
rect 4720 670 4770 680
rect 4920 670 4930 680
rect 5110 670 5120 680
rect 5150 670 5210 680
rect 5400 670 5420 680
rect 5540 670 5550 680
rect 5590 670 5600 680
rect 5660 670 5670 680
rect 5680 670 5690 680
rect 5700 670 5770 680
rect 5800 670 5810 680
rect 5860 670 5870 680
rect 6290 670 6340 680
rect 6470 670 6520 680
rect 6860 670 6880 680
rect 7390 670 7420 680
rect 7990 670 8010 680
rect 8140 670 8290 680
rect 8740 670 9090 680
rect 9330 670 9350 680
rect 10 660 600 670
rect 760 660 910 670
rect 930 660 950 670
rect 970 660 980 670
rect 1300 660 1350 670
rect 2090 660 2100 670
rect 2340 660 2350 670
rect 4140 660 4160 670
rect 4740 660 4780 670
rect 5140 660 5150 670
rect 5160 660 5180 670
rect 5190 660 5210 670
rect 5330 660 5340 670
rect 5400 660 5410 670
rect 5420 660 5430 670
rect 5560 660 5570 670
rect 5580 660 5610 670
rect 5680 660 5690 670
rect 5700 660 5760 670
rect 5860 660 5880 670
rect 5920 660 5930 670
rect 6290 660 6340 670
rect 6470 660 6540 670
rect 6870 660 6880 670
rect 7390 660 7420 670
rect 7990 660 8010 670
rect 8140 660 8310 670
rect 8740 660 9090 670
rect 9210 660 9220 670
rect 9310 660 9320 670
rect 9330 660 9340 670
rect 9600 660 9610 670
rect 0 650 590 660
rect 820 650 860 660
rect 1290 650 1340 660
rect 3270 650 3280 660
rect 4750 650 4780 660
rect 5140 650 5190 660
rect 5200 650 5210 660
rect 5290 650 5330 660
rect 5580 650 5600 660
rect 5660 650 5670 660
rect 5680 650 5690 660
rect 5700 650 5740 660
rect 5780 650 5810 660
rect 6290 650 6340 660
rect 6480 650 6540 660
rect 6870 650 6880 660
rect 7390 650 7420 660
rect 7990 650 8020 660
rect 8140 650 8320 660
rect 8730 650 9070 660
rect 9080 650 9090 660
rect 9110 650 9150 660
rect 9320 650 9340 660
rect 9590 650 9620 660
rect 0 640 580 650
rect 1290 640 1330 650
rect 2100 640 2110 650
rect 3250 640 3260 650
rect 4760 640 4830 650
rect 5160 640 5180 650
rect 5210 640 5220 650
rect 5290 640 5320 650
rect 5360 640 5370 650
rect 5430 640 5440 650
rect 5500 640 5510 650
rect 5530 640 5540 650
rect 5600 640 5610 650
rect 5700 640 5750 650
rect 5820 640 5850 650
rect 6280 640 6340 650
rect 6480 640 6530 650
rect 6870 640 6880 650
rect 7380 640 7420 650
rect 8000 640 8020 650
rect 8140 640 8330 650
rect 8710 640 9090 650
rect 9110 640 9130 650
rect 9300 640 9310 650
rect 9320 640 9330 650
rect 9590 640 9620 650
rect 0 630 520 640
rect 1280 630 1330 640
rect 2110 630 2120 640
rect 2290 630 2300 640
rect 3230 630 3240 640
rect 4760 630 4810 640
rect 5280 630 5290 640
rect 5300 630 5320 640
rect 5360 630 5370 640
rect 5400 630 5440 640
rect 5510 630 5520 640
rect 5530 630 5540 640
rect 5590 630 5600 640
rect 5700 630 5780 640
rect 5820 630 5850 640
rect 6280 630 6340 640
rect 6490 630 6530 640
rect 6870 630 6880 640
rect 7380 630 7420 640
rect 8000 630 8020 640
rect 8140 630 8340 640
rect 8690 630 8700 640
rect 8710 630 9080 640
rect 9110 630 9130 640
rect 9590 630 9630 640
rect 0 620 480 630
rect 1280 620 1330 630
rect 1360 620 1390 630
rect 2110 620 2120 630
rect 3160 620 3220 630
rect 4780 620 4790 630
rect 4930 620 4940 630
rect 5280 620 5290 630
rect 5310 620 5320 630
rect 5360 620 5370 630
rect 5400 620 5440 630
rect 5510 620 5520 630
rect 5540 620 5550 630
rect 5680 620 5690 630
rect 5700 620 5850 630
rect 6290 620 6340 630
rect 6500 620 6540 630
rect 6870 620 6890 630
rect 7380 620 7420 630
rect 8010 620 8030 630
rect 8140 620 8360 630
rect 8690 620 8700 630
rect 8720 620 9080 630
rect 9100 620 9140 630
rect 9290 620 9320 630
rect 0 610 450 620
rect 1260 610 1410 620
rect 2110 610 2120 620
rect 2260 610 2270 620
rect 3140 610 3150 620
rect 4770 610 4780 620
rect 5280 610 5290 620
rect 5360 610 5370 620
rect 5420 610 5430 620
rect 5440 610 5450 620
rect 5550 610 5560 620
rect 5590 610 5620 620
rect 5630 610 5640 620
rect 5680 610 5690 620
rect 5700 610 5820 620
rect 6300 610 6340 620
rect 6510 610 6540 620
rect 6870 610 6890 620
rect 7380 610 7420 620
rect 8010 610 8040 620
rect 8140 610 8360 620
rect 8700 610 9070 620
rect 9100 610 9140 620
rect 9210 610 9220 620
rect 0 600 420 610
rect 1250 600 1320 610
rect 1390 600 1400 610
rect 1410 600 1420 610
rect 2110 600 2120 610
rect 4760 600 4770 610
rect 5560 600 5570 610
rect 5680 600 5690 610
rect 5700 600 5850 610
rect 6300 600 6340 610
rect 6510 600 6550 610
rect 6880 600 6890 610
rect 7380 600 7420 610
rect 8010 600 8050 610
rect 8140 600 8370 610
rect 8670 600 9070 610
rect 9100 600 9120 610
rect 9210 600 9230 610
rect 0 590 390 600
rect 1250 590 1300 600
rect 1420 590 1430 600
rect 3120 590 3130 600
rect 4060 590 4080 600
rect 4550 590 4560 600
rect 4740 590 4760 600
rect 5450 590 5460 600
rect 5570 590 5590 600
rect 5680 590 5690 600
rect 5700 590 5850 600
rect 6310 590 6340 600
rect 6510 590 6560 600
rect 6880 590 6890 600
rect 7380 590 7420 600
rect 8020 590 8060 600
rect 8140 590 8390 600
rect 8650 590 9050 600
rect 9070 590 9100 600
rect 9290 590 9300 600
rect 0 580 370 590
rect 1230 580 1290 590
rect 2120 580 2130 590
rect 2210 580 2220 590
rect 3050 580 3090 590
rect 3110 580 3120 590
rect 4070 580 4080 590
rect 4550 580 4560 590
rect 4710 580 4720 590
rect 4730 580 4760 590
rect 4940 580 4950 590
rect 5240 580 5250 590
rect 5450 580 5460 590
rect 5540 580 5550 590
rect 5580 580 5590 590
rect 5680 580 5690 590
rect 5700 580 5880 590
rect 6320 580 6340 590
rect 6520 580 6570 590
rect 6880 580 6900 590
rect 7380 580 7420 590
rect 8030 580 8060 590
rect 8140 580 8400 590
rect 8650 580 9050 590
rect 9140 580 9170 590
rect 9290 580 9300 590
rect 0 570 350 580
rect 1210 570 1280 580
rect 3040 570 3050 580
rect 4540 570 4560 580
rect 4740 570 4750 580
rect 5230 570 5240 580
rect 5250 570 5260 580
rect 5280 570 5290 580
rect 5540 570 5550 580
rect 5580 570 5590 580
rect 5600 570 5610 580
rect 5680 570 5690 580
rect 5700 570 5880 580
rect 6320 570 6340 580
rect 6520 570 6570 580
rect 6890 570 6900 580
rect 7370 570 7420 580
rect 8040 570 8070 580
rect 8140 570 8430 580
rect 8570 570 8590 580
rect 8650 570 9050 580
rect 9150 570 9170 580
rect 9220 570 9230 580
rect 9280 570 9290 580
rect 0 560 330 570
rect 1190 560 1260 570
rect 3020 560 3030 570
rect 4530 560 4540 570
rect 4700 560 4710 570
rect 4730 560 4750 570
rect 5250 560 5270 570
rect 5460 560 5470 570
rect 5590 560 5610 570
rect 5680 560 5690 570
rect 5700 560 5850 570
rect 5910 560 5930 570
rect 6320 560 6340 570
rect 6520 560 6580 570
rect 6890 560 6900 570
rect 7370 560 7420 570
rect 8050 560 8080 570
rect 8130 560 8440 570
rect 8570 560 8600 570
rect 8610 560 9040 570
rect 9100 560 9120 570
rect 9160 560 9170 570
rect 9280 560 9290 570
rect 0 550 310 560
rect 1160 550 1250 560
rect 2140 550 2170 560
rect 4510 550 4530 560
rect 4540 550 4550 560
rect 4700 550 4710 560
rect 4730 550 4750 560
rect 5470 550 5480 560
rect 5570 550 5580 560
rect 5600 550 5630 560
rect 5680 550 5690 560
rect 5700 550 5850 560
rect 5880 550 5910 560
rect 5920 550 5930 560
rect 6320 550 6340 560
rect 6530 550 6580 560
rect 6890 550 6900 560
rect 7370 550 7420 560
rect 8060 550 8090 560
rect 8110 550 8440 560
rect 8450 550 8460 560
rect 8470 550 8480 560
rect 8560 550 9040 560
rect 9100 550 9140 560
rect 9170 550 9180 560
rect 9280 550 9290 560
rect 0 540 290 550
rect 1140 540 1240 550
rect 1470 540 1480 550
rect 4500 540 4510 550
rect 4680 540 4690 550
rect 4730 540 4750 550
rect 5470 540 5480 550
rect 5620 540 5630 550
rect 5680 540 5690 550
rect 5700 540 5840 550
rect 5850 540 5930 550
rect 6320 540 6340 550
rect 6540 540 6580 550
rect 6890 540 6900 550
rect 7360 540 7420 550
rect 8070 540 8470 550
rect 8500 540 8520 550
rect 8530 540 9070 550
rect 9080 540 9120 550
rect 9240 540 9250 550
rect 9270 540 9280 550
rect 0 530 260 540
rect 670 530 700 540
rect 1100 530 1230 540
rect 1480 530 1490 540
rect 2970 530 2980 540
rect 4480 530 4500 540
rect 4530 530 4540 540
rect 4680 530 4690 540
rect 4720 530 4740 540
rect 5430 530 5470 540
rect 5480 530 5490 540
rect 5570 530 5580 540
rect 5620 530 5630 540
rect 5670 530 5690 540
rect 5700 530 5890 540
rect 5900 530 5930 540
rect 5940 530 5950 540
rect 6000 530 6010 540
rect 6320 530 6340 540
rect 6540 530 6590 540
rect 6900 530 6910 540
rect 7360 530 7420 540
rect 8080 530 9040 540
rect 9060 530 9070 540
rect 9080 530 9100 540
rect 9160 530 9170 540
rect 9260 530 9270 540
rect 9960 530 9990 540
rect 0 520 230 530
rect 670 520 710 530
rect 750 520 780 530
rect 830 520 870 530
rect 1090 520 1220 530
rect 2950 520 2960 530
rect 4470 520 4480 530
rect 4530 520 4540 530
rect 4720 520 4740 530
rect 5390 520 5400 530
rect 5430 520 5500 530
rect 5590 520 5610 530
rect 5630 520 5640 530
rect 5670 520 5680 530
rect 5700 520 5970 530
rect 6330 520 6340 530
rect 6550 520 6600 530
rect 7370 520 7420 530
rect 8080 520 9040 530
rect 9070 520 9090 530
rect 9160 520 9170 530
rect 9250 520 9270 530
rect 9970 520 9990 530
rect 0 510 210 520
rect 320 510 340 520
rect 660 510 880 520
rect 1090 510 1210 520
rect 2900 510 2930 520
rect 4440 510 4470 520
rect 4530 510 4540 520
rect 4720 510 4740 520
rect 5370 510 5400 520
rect 5420 510 5480 520
rect 5640 510 5650 520
rect 5670 510 5680 520
rect 5700 510 5870 520
rect 5890 510 5930 520
rect 6320 510 6330 520
rect 6560 510 6600 520
rect 7360 510 7420 520
rect 8100 510 9050 520
rect 9070 510 9090 520
rect 9250 510 9260 520
rect 9930 510 9940 520
rect 9980 510 9990 520
rect 0 500 190 510
rect 320 500 350 510
rect 660 500 890 510
rect 1090 500 1190 510
rect 1510 500 1520 510
rect 2870 500 2880 510
rect 4410 500 4460 510
rect 4530 500 4540 510
rect 4720 500 4740 510
rect 5360 500 5400 510
rect 5420 500 5470 510
rect 5490 500 5500 510
rect 5650 500 5660 510
rect 5670 500 5680 510
rect 5700 500 5870 510
rect 5880 500 5930 510
rect 5950 500 5960 510
rect 6310 500 6330 510
rect 6560 500 6610 510
rect 7370 500 7420 510
rect 8100 500 9050 510
rect 9070 500 9100 510
rect 9130 500 9140 510
rect 9150 500 9160 510
rect 9170 500 9180 510
rect 9250 500 9260 510
rect 9920 500 9930 510
rect 0 490 170 500
rect 340 490 360 500
rect 650 490 900 500
rect 1090 490 1180 500
rect 1520 490 1530 500
rect 2850 490 2860 500
rect 4400 490 4430 500
rect 4530 490 4540 500
rect 4720 490 4740 500
rect 5360 490 5400 500
rect 5420 490 5470 500
rect 5490 490 5510 500
rect 5630 490 5640 500
rect 5660 490 5670 500
rect 5700 490 5800 500
rect 5820 490 5850 500
rect 5860 490 5870 500
rect 5900 490 5920 500
rect 6310 490 6330 500
rect 6570 490 6620 500
rect 7350 490 7420 500
rect 8110 490 9030 500
rect 9050 490 9080 500
rect 9210 490 9220 500
rect 9920 490 9930 500
rect 9940 490 9950 500
rect 9990 490 9990 500
rect 0 480 160 490
rect 350 480 370 490
rect 650 480 810 490
rect 830 480 900 490
rect 1090 480 1170 490
rect 2820 480 2830 490
rect 4310 480 4400 490
rect 4530 480 4550 490
rect 4720 480 4740 490
rect 4960 480 4970 490
rect 5360 480 5390 490
rect 5420 480 5460 490
rect 5630 480 5640 490
rect 5700 480 5810 490
rect 5830 480 5880 490
rect 5890 480 5910 490
rect 5920 480 5940 490
rect 6320 480 6330 490
rect 6570 480 6620 490
rect 7350 480 7410 490
rect 8120 480 9030 490
rect 9070 480 9080 490
rect 9120 480 9130 490
rect 9240 480 9250 490
rect 9860 480 9880 490
rect 9910 480 9940 490
rect 0 470 150 480
rect 350 470 380 480
rect 560 470 650 480
rect 660 470 690 480
rect 770 470 790 480
rect 820 470 920 480
rect 1090 470 1160 480
rect 2780 470 2790 480
rect 4260 470 4280 480
rect 4290 470 4380 480
rect 4450 470 4490 480
rect 4530 470 4550 480
rect 4720 470 4740 480
rect 5360 470 5380 480
rect 5430 470 5450 480
rect 5700 470 5800 480
rect 5840 470 5940 480
rect 6300 470 6320 480
rect 6570 470 6620 480
rect 7350 470 7420 480
rect 8160 470 9060 480
rect 9080 470 9110 480
rect 9230 470 9240 480
rect 9870 470 9880 480
rect 9910 470 9920 480
rect 0 460 140 470
rect 360 460 390 470
rect 550 460 640 470
rect 670 460 680 470
rect 820 460 940 470
rect 1080 460 1150 470
rect 2110 460 2120 470
rect 2150 460 2160 470
rect 2750 460 2760 470
rect 4260 460 4280 470
rect 4290 460 4330 470
rect 4440 460 4490 470
rect 4530 460 4550 470
rect 4710 460 4740 470
rect 5610 460 5620 470
rect 5700 460 5810 470
rect 5830 460 5840 470
rect 5860 460 5940 470
rect 5950 460 5970 470
rect 6290 460 6320 470
rect 6580 460 6620 470
rect 7350 460 7420 470
rect 8170 460 9040 470
rect 9080 460 9090 470
rect 9230 460 9240 470
rect 9860 460 9880 470
rect 0 450 130 460
rect 370 450 400 460
rect 550 450 630 460
rect 660 450 680 460
rect 810 450 950 460
rect 1060 450 1140 460
rect 1540 450 1550 460
rect 2700 450 2710 460
rect 4270 450 4290 460
rect 4440 450 4500 460
rect 4530 450 4560 460
rect 4700 450 4740 460
rect 5260 450 5270 460
rect 5700 450 5810 460
rect 5870 450 5950 460
rect 6270 450 6330 460
rect 6590 450 6630 460
rect 7350 450 7410 460
rect 8180 450 9010 460
rect 9040 450 9050 460
rect 9870 450 9880 460
rect 0 440 120 450
rect 380 440 410 450
rect 560 440 630 450
rect 670 440 680 450
rect 800 440 1010 450
rect 1020 440 1130 450
rect 2010 440 2020 450
rect 2660 440 2670 450
rect 4290 440 4310 450
rect 4430 440 4480 450
rect 4490 440 4510 450
rect 4540 440 4570 450
rect 4700 440 4720 450
rect 5230 440 5240 450
rect 5250 440 5270 450
rect 5710 440 5810 450
rect 5820 440 5830 450
rect 5870 440 5950 450
rect 6280 440 6330 450
rect 6600 440 6640 450
rect 7350 440 7410 450
rect 8210 440 9000 450
rect 9020 440 9030 450
rect 9040 440 9050 450
rect 0 430 110 440
rect 380 430 390 440
rect 400 430 410 440
rect 560 430 610 440
rect 670 430 680 440
rect 790 430 1120 440
rect 1850 430 1860 440
rect 1970 430 1980 440
rect 2630 430 2640 440
rect 4290 430 4320 440
rect 4430 430 4480 440
rect 4490 430 4510 440
rect 4540 430 4590 440
rect 4630 430 4690 440
rect 4700 430 4720 440
rect 5230 430 5240 440
rect 5260 430 5270 440
rect 5710 430 5840 440
rect 5860 430 5970 440
rect 6280 430 6340 440
rect 6600 430 6650 440
rect 7350 430 7410 440
rect 8230 430 8990 440
rect 9030 430 9050 440
rect 9090 430 9100 440
rect 9180 430 9190 440
rect 0 420 100 430
rect 390 420 400 430
rect 410 420 420 430
rect 550 420 560 430
rect 570 420 600 430
rect 670 420 680 430
rect 780 420 1120 430
rect 1810 420 1830 430
rect 2310 420 2320 430
rect 4270 420 4320 430
rect 4430 420 4510 430
rect 4550 420 4670 430
rect 4680 420 4690 430
rect 4700 420 4720 430
rect 5230 420 5240 430
rect 5260 420 5270 430
rect 5300 420 5310 430
rect 5710 420 5810 430
rect 5860 420 5980 430
rect 6270 420 6340 430
rect 6610 420 6650 430
rect 7350 420 7420 430
rect 8250 420 8990 430
rect 9090 420 9130 430
rect 0 410 90 420
rect 560 410 590 420
rect 670 410 680 420
rect 770 410 1110 420
rect 2360 410 2370 420
rect 4260 410 4310 420
rect 4340 410 4370 420
rect 4430 410 4480 420
rect 4490 410 4510 420
rect 4550 410 4690 420
rect 4710 410 4720 420
rect 5150 410 5160 420
rect 5230 410 5240 420
rect 5250 410 5270 420
rect 5340 410 5360 420
rect 5710 410 5820 420
rect 5850 410 5980 420
rect 6270 410 6340 420
rect 6620 410 6670 420
rect 7350 410 7420 420
rect 8260 410 8990 420
rect 9090 410 9100 420
rect 9120 410 9130 420
rect 9200 410 9210 420
rect 0 400 80 410
rect 400 400 410 410
rect 420 400 430 410
rect 560 400 570 410
rect 670 400 680 410
rect 770 400 1110 410
rect 4250 400 4310 410
rect 4320 400 4340 410
rect 4350 400 4380 410
rect 4420 400 4440 410
rect 4450 400 4460 410
rect 4490 400 4510 410
rect 4550 400 4680 410
rect 4700 400 4720 410
rect 5150 400 5160 410
rect 5220 400 5240 410
rect 5250 400 5270 410
rect 5340 400 5360 410
rect 5720 400 5990 410
rect 6000 400 6010 410
rect 6280 400 6340 410
rect 6620 400 6680 410
rect 7340 400 7420 410
rect 8270 400 9010 410
rect 9060 400 9080 410
rect 9090 400 9120 410
rect 0 390 80 400
rect 400 390 410 400
rect 420 390 430 400
rect 670 390 680 400
rect 770 390 1100 400
rect 4260 390 4300 400
rect 4310 390 4320 400
rect 4360 390 4380 400
rect 4430 390 4460 400
rect 4470 390 4500 400
rect 4550 390 4560 400
rect 4570 390 4680 400
rect 4710 390 4720 400
rect 5150 390 5160 400
rect 5220 390 5270 400
rect 5340 390 5360 400
rect 5730 390 6000 400
rect 6270 390 6340 400
rect 6620 390 6690 400
rect 7330 390 7420 400
rect 8290 390 8980 400
rect 9060 390 9070 400
rect 9080 390 9110 400
rect 9190 390 9200 400
rect 9330 390 9350 400
rect 0 380 70 390
rect 400 380 420 390
rect 430 380 440 390
rect 670 380 680 390
rect 770 380 1090 390
rect 4250 380 4290 390
rect 4300 380 4310 390
rect 4370 380 4390 390
rect 4430 380 4490 390
rect 4550 380 4560 390
rect 4580 380 4680 390
rect 4710 380 4720 390
rect 4970 380 4980 390
rect 5210 380 5270 390
rect 5330 380 5360 390
rect 5750 380 6010 390
rect 6290 380 6340 390
rect 6640 380 6700 390
rect 7330 380 7420 390
rect 8280 380 8970 390
rect 9060 380 9070 390
rect 9150 380 9160 390
rect 9180 380 9190 390
rect 9330 380 9390 390
rect 0 370 60 380
rect 410 370 420 380
rect 430 370 440 380
rect 670 370 680 380
rect 780 370 1080 380
rect 4250 370 4280 380
rect 4290 370 4300 380
rect 4380 370 4400 380
rect 4590 370 4670 380
rect 4710 370 4720 380
rect 4970 370 4980 380
rect 5210 370 5240 380
rect 5250 370 5260 380
rect 5330 370 5380 380
rect 5760 370 6000 380
rect 6290 370 6350 380
rect 6650 370 6700 380
rect 7330 370 7420 380
rect 8290 370 8840 380
rect 8860 370 8980 380
rect 9060 370 9070 380
rect 9090 370 9100 380
rect 9320 370 9400 380
rect 0 360 60 370
rect 410 360 420 370
rect 560 360 570 370
rect 580 360 600 370
rect 610 360 650 370
rect 670 360 680 370
rect 800 360 810 370
rect 920 360 1080 370
rect 4240 360 4270 370
rect 4280 360 4290 370
rect 4390 360 4420 370
rect 4600 360 4690 370
rect 4700 360 4720 370
rect 4970 360 4980 370
rect 5210 360 5250 370
rect 5320 360 5380 370
rect 5660 360 5670 370
rect 5770 360 5810 370
rect 5840 360 6000 370
rect 6280 360 6340 370
rect 6650 360 6710 370
rect 7330 360 7420 370
rect 8300 360 8830 370
rect 8860 360 8980 370
rect 9000 360 9030 370
rect 9060 360 9090 370
rect 9170 360 9180 370
rect 9250 360 9290 370
rect 9330 360 9400 370
rect 0 350 50 360
rect 410 350 420 360
rect 440 350 450 360
rect 530 350 650 360
rect 660 350 680 360
rect 950 350 1070 360
rect 4230 350 4240 360
rect 4250 350 4280 360
rect 4400 350 4470 360
rect 4500 350 4540 360
rect 4550 350 4560 360
rect 4610 350 4720 360
rect 5210 350 5250 360
rect 5330 350 5370 360
rect 5780 350 5790 360
rect 5840 350 6010 360
rect 6280 350 6340 360
rect 6670 350 6720 360
rect 7330 350 7420 360
rect 8310 350 8810 360
rect 8850 350 8980 360
rect 9000 350 9080 360
rect 9160 350 9170 360
rect 9250 350 9260 360
rect 9290 350 9310 360
rect 9320 350 9430 360
rect 9980 350 9990 360
rect 0 340 50 350
rect 440 340 450 350
rect 510 340 550 350
rect 1010 340 1060 350
rect 4260 340 4270 350
rect 4470 340 4480 350
rect 4490 340 4510 350
rect 4530 340 4560 350
rect 4620 340 4690 350
rect 4710 340 4720 350
rect 5120 340 5130 350
rect 5210 340 5250 350
rect 5330 340 5370 350
rect 5670 340 5680 350
rect 5740 340 5760 350
rect 5790 340 5800 350
rect 5850 340 6000 350
rect 6280 340 6340 350
rect 6680 340 6720 350
rect 7330 340 7420 350
rect 8320 340 8800 350
rect 8850 340 8980 350
rect 9020 340 9030 350
rect 9040 340 9100 350
rect 9130 340 9140 350
rect 9230 340 9240 350
rect 9260 340 9270 350
rect 9300 340 9380 350
rect 0 330 40 340
rect 420 330 430 340
rect 440 330 450 340
rect 700 330 720 340
rect 1030 330 1050 340
rect 4250 330 4260 340
rect 4470 330 4500 340
rect 4540 330 4570 340
rect 4600 330 4680 340
rect 5110 330 5140 340
rect 5210 330 5220 340
rect 5230 330 5240 340
rect 5340 330 5360 340
rect 5670 330 5680 340
rect 5730 330 5770 340
rect 5810 330 5820 340
rect 5860 330 6010 340
rect 6270 330 6340 340
rect 6680 330 6740 340
rect 7320 330 7420 340
rect 8320 330 8800 340
rect 8850 330 8880 340
rect 8900 330 8990 340
rect 9030 330 9040 340
rect 9230 330 9240 340
rect 9250 330 9280 340
rect 9300 330 9320 340
rect 9350 330 9380 340
rect 9410 330 9420 340
rect 0 320 30 330
rect 420 320 430 330
rect 440 320 480 330
rect 730 320 780 330
rect 1040 320 1050 330
rect 4480 320 4490 330
rect 4550 320 4660 330
rect 5110 320 5130 330
rect 5200 320 5220 330
rect 5670 320 5680 330
rect 5720 320 5790 330
rect 5820 320 5830 330
rect 5860 320 6010 330
rect 6280 320 6340 330
rect 6690 320 6740 330
rect 7320 320 7420 330
rect 8330 320 8800 330
rect 8810 320 8880 330
rect 8890 320 9000 330
rect 9140 320 9150 330
rect 9220 320 9320 330
rect 9360 320 9390 330
rect 0 310 30 320
rect 420 310 430 320
rect 450 310 470 320
rect 790 310 810 320
rect 1030 310 1040 320
rect 4480 310 4490 320
rect 4560 310 4620 320
rect 4650 310 4660 320
rect 5200 310 5210 320
rect 5680 310 5690 320
rect 5720 310 5810 320
rect 5840 310 5850 320
rect 5860 310 6010 320
rect 6260 310 6340 320
rect 6690 310 6750 320
rect 7320 310 7410 320
rect 8350 310 8940 320
rect 8950 310 9000 320
rect 9030 310 9040 320
rect 9110 310 9120 320
rect 9220 310 9300 320
rect 9400 310 9410 320
rect 0 300 30 310
rect 430 300 440 310
rect 450 300 470 310
rect 820 300 870 310
rect 880 300 930 310
rect 940 300 1000 310
rect 1030 300 1040 310
rect 1270 300 1290 310
rect 4560 300 4570 310
rect 4590 300 4620 310
rect 4650 300 4660 310
rect 5720 300 5800 310
rect 5810 300 5830 310
rect 5850 300 6000 310
rect 6270 300 6350 310
rect 6700 300 6770 310
rect 7320 300 7410 310
rect 8350 300 8900 310
rect 8940 300 9010 310
rect 9050 300 9070 310
rect 9130 300 9140 310
rect 9250 300 9300 310
rect 9390 300 9410 310
rect 0 290 20 300
rect 430 290 440 300
rect 450 290 460 300
rect 990 290 1030 300
rect 1260 290 1270 300
rect 1280 290 1310 300
rect 4560 290 4580 300
rect 4590 290 4630 300
rect 5720 290 5840 300
rect 5860 290 5990 300
rect 6280 290 6350 300
rect 6700 290 6780 300
rect 7320 290 7420 300
rect 8370 290 8900 300
rect 8930 290 9020 300
rect 9050 290 9060 300
rect 9210 290 9220 300
rect 9270 290 9310 300
rect 9400 290 9420 300
rect 0 280 20 290
rect 430 280 440 290
rect 1010 280 1030 290
rect 1250 280 1310 290
rect 4570 280 4590 290
rect 4620 280 4650 290
rect 4980 280 4990 290
rect 5070 280 5080 290
rect 5720 280 5830 290
rect 5880 280 5990 290
rect 6070 280 6130 290
rect 6270 280 6350 290
rect 6710 280 6790 290
rect 7320 280 7420 290
rect 8360 280 8910 290
rect 8930 280 8950 290
rect 8970 280 8990 290
rect 9020 280 9030 290
rect 9120 280 9130 290
rect 9280 280 9310 290
rect 9410 280 9420 290
rect 0 270 20 280
rect 430 270 440 280
rect 1000 270 1030 280
rect 1240 270 1290 280
rect 4570 270 4590 280
rect 4630 270 4650 280
rect 5730 270 5780 280
rect 5790 270 5830 280
rect 5900 270 6000 280
rect 6040 270 6060 280
rect 6110 270 6130 280
rect 6280 270 6360 280
rect 6710 270 6790 280
rect 7330 270 7410 280
rect 8370 270 8900 280
rect 8930 270 8940 280
rect 9020 270 9050 280
rect 9110 270 9120 280
rect 9210 270 9240 280
rect 9320 270 9330 280
rect 9420 270 9430 280
rect 0 260 10 270
rect 420 260 440 270
rect 1000 260 1020 270
rect 1240 260 1280 270
rect 4580 260 4590 270
rect 4630 260 4650 270
rect 5740 260 5830 270
rect 5920 260 6030 270
rect 6110 260 6130 270
rect 6280 260 6360 270
rect 6720 260 6810 270
rect 7320 260 7410 270
rect 8380 260 8890 270
rect 8930 260 8950 270
rect 9030 260 9050 270
rect 9110 260 9120 270
rect 9230 260 9240 270
rect 9260 260 9270 270
rect 9330 260 9340 270
rect 9420 260 9430 270
rect 0 250 10 260
rect 420 250 430 260
rect 1010 250 1020 260
rect 1240 250 1270 260
rect 4580 250 4590 260
rect 5740 250 5810 260
rect 5940 250 6010 260
rect 6100 250 6130 260
rect 6270 250 6360 260
rect 6730 250 6810 260
rect 7330 250 7410 260
rect 8390 250 8880 260
rect 8940 250 8960 260
rect 9230 250 9260 260
rect 9350 250 9370 260
rect 9410 250 9430 260
rect 0 240 10 250
rect 410 240 430 250
rect 4580 240 4590 250
rect 5710 240 5780 250
rect 6040 240 6070 250
rect 6090 240 6120 250
rect 6280 240 6360 250
rect 6740 240 6830 250
rect 7320 240 7410 250
rect 8400 240 8880 250
rect 8960 240 8970 250
rect 9030 240 9040 250
rect 9100 240 9110 250
rect 9200 240 9210 250
rect 9340 240 9360 250
rect 9790 240 9810 250
rect 0 230 10 240
rect 410 230 420 240
rect 5670 230 5680 240
rect 6010 230 6080 240
rect 6090 230 6110 240
rect 6290 230 6360 240
rect 6750 230 6830 240
rect 6840 230 6850 240
rect 7320 230 7410 240
rect 8400 230 8870 240
rect 9170 230 9190 240
rect 9330 230 9360 240
rect 9790 230 9810 240
rect 9830 230 9840 240
rect 0 220 10 230
rect 400 220 420 230
rect 5940 220 5950 230
rect 5970 220 6040 230
rect 6060 220 6110 230
rect 6290 220 6360 230
rect 6750 220 6850 230
rect 7320 220 7410 230
rect 8420 220 8870 230
rect 9020 220 9030 230
rect 9060 220 9070 230
rect 9090 220 9100 230
rect 9190 220 9200 230
rect 9330 220 9370 230
rect 9800 220 9810 230
rect 9820 220 9830 230
rect 0 210 10 220
rect 160 210 200 220
rect 400 210 420 220
rect 5610 210 5620 220
rect 5720 210 5730 220
rect 5990 210 6030 220
rect 6060 210 6110 220
rect 6290 210 6360 220
rect 6760 210 6850 220
rect 6860 210 6870 220
rect 7310 210 7410 220
rect 8430 210 8860 220
rect 9080 210 9090 220
rect 9170 210 9190 220
rect 9810 210 9840 220
rect 0 200 10 210
rect 140 200 210 210
rect 390 200 420 210
rect 1000 200 1010 210
rect 5720 200 5740 210
rect 6000 200 6010 210
rect 6020 200 6030 210
rect 6060 200 6100 210
rect 6300 200 6370 210
rect 6780 200 6880 210
rect 7310 200 7410 210
rect 8440 200 8700 210
rect 8710 200 8860 210
rect 8960 200 8970 210
rect 9010 200 9020 210
rect 9240 200 9280 210
rect 9810 200 9830 210
rect 110 190 180 200
rect 200 190 210 200
rect 380 190 420 200
rect 5720 190 5750 200
rect 6020 190 6030 200
rect 6040 190 6090 200
rect 6310 190 6370 200
rect 6790 190 6900 200
rect 6910 190 6920 200
rect 7320 190 7400 200
rect 8450 190 8600 200
rect 8630 190 8650 200
rect 8670 190 8690 200
rect 8740 190 8860 200
rect 8920 190 8950 200
rect 9070 190 9080 200
rect 9160 190 9170 200
rect 9230 190 9290 200
rect 9800 190 9810 200
rect 9820 190 9850 200
rect 120 180 160 190
rect 380 180 400 190
rect 420 180 430 190
rect 5000 180 5010 190
rect 5450 180 5490 190
rect 5610 180 5620 190
rect 5720 180 5740 190
rect 5970 180 5980 190
rect 6000 180 6010 190
rect 6020 180 6030 190
rect 6040 180 6090 190
rect 6310 180 6370 190
rect 6790 180 6930 190
rect 7330 180 7410 190
rect 8460 180 8570 190
rect 8680 180 8690 190
rect 8760 180 8840 190
rect 8910 180 8930 190
rect 9170 180 9180 190
rect 9210 180 9250 190
rect 9260 180 9270 190
rect 9290 180 9300 190
rect 9740 180 9790 190
rect 9820 180 9830 190
rect 9940 180 9950 190
rect 9970 180 9980 190
rect 140 170 180 180
rect 210 170 220 180
rect 370 170 400 180
rect 420 170 430 180
rect 5370 170 5420 180
rect 5450 170 5540 180
rect 5580 170 5590 180
rect 5690 170 5700 180
rect 5970 170 5980 180
rect 6000 170 6010 180
rect 6020 170 6080 180
rect 6310 170 6380 180
rect 6800 170 6940 180
rect 7320 170 7400 180
rect 8460 170 8580 180
rect 8750 170 8840 180
rect 9130 170 9140 180
rect 9200 170 9220 180
rect 9320 170 9330 180
rect 9730 170 9790 180
rect 9830 170 9840 180
rect 9890 170 9950 180
rect 9970 170 9980 180
rect 9990 170 9990 180
rect 140 160 220 170
rect 360 160 400 170
rect 430 160 440 170
rect 5350 160 5660 170
rect 5930 160 5980 170
rect 6000 160 6070 170
rect 6080 160 6090 170
rect 6320 160 6390 170
rect 6800 160 6960 170
rect 6970 160 6980 170
rect 7320 160 7400 170
rect 8480 160 8580 170
rect 8750 160 8830 170
rect 8900 160 8910 170
rect 9130 160 9140 170
rect 9150 160 9160 170
rect 9190 160 9200 170
rect 9320 160 9330 170
rect 9720 160 9750 170
rect 9760 160 9780 170
rect 9830 160 9840 170
rect 9890 160 9900 170
rect 9920 160 9940 170
rect 9980 160 9990 170
rect 150 150 230 160
rect 350 150 400 160
rect 430 150 450 160
rect 460 150 500 160
rect 4360 150 4380 160
rect 5360 150 5700 160
rect 5950 150 5980 160
rect 6000 150 6040 160
rect 6070 150 6100 160
rect 6330 150 6390 160
rect 6810 150 6990 160
rect 7330 150 7400 160
rect 8490 150 8570 160
rect 8730 150 8830 160
rect 8890 150 8900 160
rect 9070 150 9080 160
rect 9140 150 9150 160
rect 9180 150 9210 160
rect 9330 150 9340 160
rect 9710 150 9720 160
rect 9740 150 9750 160
rect 9760 150 9790 160
rect 9930 150 9940 160
rect 9970 150 9990 160
rect 150 140 230 150
rect 340 140 390 150
rect 450 140 570 150
rect 4340 140 4400 150
rect 5340 140 5720 150
rect 5970 140 5980 150
rect 5990 140 6030 150
rect 6050 140 6100 150
rect 6330 140 6400 150
rect 6810 140 6990 150
rect 7320 140 7400 150
rect 8500 140 8570 150
rect 8730 140 8830 150
rect 9140 140 9150 150
rect 9160 140 9170 150
rect 9180 140 9190 150
rect 9210 140 9220 150
rect 9310 140 9320 150
rect 9710 140 9720 150
rect 9740 140 9770 150
rect 9820 140 9830 150
rect 9880 140 9890 150
rect 9930 140 9940 150
rect 160 130 240 140
rect 330 130 390 140
rect 460 130 580 140
rect 4320 130 4430 140
rect 5340 130 5740 140
rect 5970 130 6010 140
rect 6040 130 6100 140
rect 6320 130 6400 140
rect 6820 130 7000 140
rect 7330 130 7390 140
rect 8500 130 8570 140
rect 8740 130 8830 140
rect 9080 130 9090 140
rect 9150 130 9170 140
rect 9180 130 9190 140
rect 9340 130 9350 140
rect 9750 130 9770 140
rect 9820 130 9830 140
rect 9920 130 9950 140
rect 160 120 250 130
rect 320 120 390 130
rect 480 120 560 130
rect 4290 120 4460 130
rect 4900 120 4940 130
rect 5340 120 5750 130
rect 5770 120 5790 130
rect 5870 120 5880 130
rect 5930 120 5990 130
rect 6010 120 6100 130
rect 6320 120 6410 130
rect 6820 120 7030 130
rect 7320 120 7390 130
rect 8510 120 8570 130
rect 8730 120 8830 130
rect 8930 120 8940 130
rect 9050 120 9060 130
rect 9160 120 9190 130
rect 9210 120 9220 130
rect 9340 120 9350 130
rect 9720 120 9730 130
rect 9740 120 9760 130
rect 9860 120 9870 130
rect 9910 120 9920 130
rect 9930 120 9940 130
rect 9960 120 9980 130
rect 150 110 220 120
rect 240 110 250 120
rect 320 110 390 120
rect 500 110 560 120
rect 4280 110 4470 120
rect 4880 110 4940 120
rect 5020 110 5030 120
rect 5350 110 5750 120
rect 5770 110 5840 120
rect 5890 110 5900 120
rect 6020 110 6100 120
rect 6330 110 6410 120
rect 6820 110 7030 120
rect 7320 110 7390 120
rect 8520 110 8570 120
rect 8730 110 8830 120
rect 8940 110 8960 120
rect 9090 110 9100 120
rect 9160 110 9180 120
rect 9210 110 9220 120
rect 9360 110 9370 120
rect 9740 110 9750 120
rect 9880 110 9890 120
rect 9940 110 9990 120
rect 160 100 220 110
rect 250 100 260 110
rect 320 100 380 110
rect 520 100 570 110
rect 760 100 780 110
rect 790 100 800 110
rect 4280 100 4490 110
rect 4850 100 4920 110
rect 5350 100 5750 110
rect 5770 100 5830 110
rect 6020 100 6100 110
rect 6330 100 6420 110
rect 6830 100 7030 110
rect 7320 100 7390 110
rect 8540 100 8570 110
rect 8720 100 8800 110
rect 8940 100 8970 110
rect 9030 100 9040 110
rect 9060 100 9070 110
rect 9160 100 9180 110
rect 9220 100 9230 110
rect 9370 100 9380 110
rect 9390 100 9410 110
rect 9580 100 9590 110
rect 9730 100 9750 110
rect 9840 100 9850 110
rect 160 90 220 100
rect 240 90 260 100
rect 330 90 380 100
rect 520 90 580 100
rect 730 90 800 100
rect 810 90 840 100
rect 4280 90 4490 100
rect 4840 90 4920 100
rect 5360 90 5750 100
rect 5770 90 5850 100
rect 6020 90 6100 100
rect 6360 90 6420 100
rect 6830 90 7040 100
rect 7320 90 7390 100
rect 8550 90 8590 100
rect 8720 90 8790 100
rect 8940 90 8970 100
rect 9050 90 9070 100
rect 9080 90 9090 100
rect 9150 90 9180 100
rect 9240 90 9250 100
rect 9570 90 9590 100
rect 9730 90 9750 100
rect 9850 90 9870 100
rect 160 80 230 90
rect 250 80 260 90
rect 320 80 370 90
rect 540 80 610 90
rect 630 80 640 90
rect 690 80 860 90
rect 4280 80 4490 90
rect 4520 80 4530 90
rect 4820 80 4910 90
rect 5290 80 5300 90
rect 5360 80 5750 90
rect 5770 80 5890 90
rect 6000 80 6100 90
rect 6360 80 6370 90
rect 6380 80 6420 90
rect 6840 80 7050 90
rect 7320 80 7380 90
rect 8550 80 8600 90
rect 8710 80 8770 90
rect 8940 80 8980 90
rect 9070 80 9080 90
rect 9170 80 9180 90
rect 9430 80 9440 90
rect 9560 80 9570 90
rect 9580 80 9590 90
rect 9730 80 9740 90
rect 9870 80 9880 90
rect 9970 80 9990 90
rect 160 70 220 80
rect 250 70 260 80
rect 320 70 360 80
rect 560 70 860 80
rect 4310 70 4530 80
rect 4820 70 4890 80
rect 5360 70 5720 80
rect 5790 70 5890 80
rect 5970 70 6100 80
rect 6400 70 6440 80
rect 6840 70 7060 80
rect 7320 70 7380 80
rect 8570 70 8600 80
rect 8710 70 8770 80
rect 8950 70 8960 80
rect 9150 70 9160 80
rect 9170 70 9180 80
rect 9230 70 9240 80
rect 9570 70 9580 80
rect 9600 70 9610 80
rect 9870 70 9890 80
rect 9900 70 9910 80
rect 9970 70 9990 80
rect 150 60 220 70
rect 260 60 270 70
rect 320 60 360 70
rect 590 60 860 70
rect 4320 60 4530 70
rect 4590 60 4610 70
rect 4810 60 4870 70
rect 5040 60 5050 70
rect 5250 60 5260 70
rect 5370 60 5700 70
rect 5800 60 6100 70
rect 6410 60 6430 70
rect 6840 60 7070 70
rect 7080 60 7090 70
rect 7320 60 7380 70
rect 8580 60 8610 70
rect 8700 60 8770 70
rect 8960 60 8970 70
rect 9180 60 9230 70
rect 9590 60 9610 70
rect 9670 60 9680 70
rect 9690 60 9700 70
rect 9830 60 9840 70
rect 9880 60 9910 70
rect 9960 60 9970 70
rect 160 50 220 60
rect 260 50 270 60
rect 310 50 360 60
rect 620 50 880 60
rect 4340 50 4520 60
rect 4570 50 4610 60
rect 4800 50 4850 60
rect 5250 50 5260 60
rect 5370 50 5680 60
rect 5810 50 6090 60
rect 6420 50 6430 60
rect 6850 50 7100 60
rect 7110 50 7120 60
rect 7320 50 7370 60
rect 8590 50 8620 60
rect 8690 50 8760 60
rect 9210 50 9230 60
rect 9270 50 9280 60
rect 9300 50 9310 60
rect 9480 50 9490 60
rect 9540 50 9550 60
rect 9670 50 9680 60
rect 9890 50 9900 60
rect 9910 50 9920 60
rect 9970 50 9980 60
rect 9990 50 9990 60
rect 170 40 220 50
rect 310 40 350 50
rect 640 40 880 50
rect 4340 40 4520 50
rect 4560 40 4600 50
rect 4790 40 4840 50
rect 5160 40 5170 50
rect 5320 40 5330 50
rect 5380 40 5670 50
rect 5820 40 6090 50
rect 6420 40 6460 50
rect 6850 40 7130 50
rect 7320 40 7360 50
rect 8600 40 8750 50
rect 8940 40 8960 50
rect 9260 40 9270 50
rect 9290 40 9300 50
rect 9530 40 9540 50
rect 9560 40 9570 50
rect 9630 40 9640 50
rect 9680 40 9690 50
rect 9700 40 9710 50
rect 9760 40 9770 50
rect 9900 40 9930 50
rect 170 30 220 40
rect 270 30 280 40
rect 310 30 350 40
rect 640 30 700 40
rect 710 30 890 40
rect 4360 30 4600 40
rect 4780 30 4830 40
rect 5380 30 5660 40
rect 5830 30 6080 40
rect 6430 30 6460 40
rect 6860 30 7120 40
rect 7310 30 7360 40
rect 8610 30 8740 40
rect 9530 30 9570 40
rect 9700 30 9710 40
rect 9780 30 9790 40
rect 9920 30 9930 40
rect 160 20 220 30
rect 270 20 280 30
rect 310 20 350 30
rect 620 20 690 30
rect 730 20 900 30
rect 4380 20 4600 30
rect 5050 20 5060 30
rect 5310 20 5320 30
rect 5390 20 5650 30
rect 5840 20 6090 30
rect 6430 20 6470 30
rect 6870 20 7120 30
rect 7310 20 7350 30
rect 8590 20 8600 30
rect 8640 20 8660 30
rect 8700 20 8720 30
rect 8990 20 9030 30
rect 9480 20 9500 30
rect 9670 20 9680 30
rect 170 10 220 20
rect 280 10 290 20
rect 310 10 350 20
rect 620 10 680 20
rect 730 10 900 20
rect 4380 10 4590 20
rect 5340 10 5350 20
rect 5390 10 5640 20
rect 5850 10 6090 20
rect 6440 10 6470 20
rect 6880 10 7140 20
rect 7300 10 7350 20
rect 8630 10 8660 20
rect 8700 10 8710 20
rect 9100 10 9110 20
rect 9180 10 9190 20
rect 9670 10 9710 20
rect 170 0 220 10
rect 270 0 290 10
rect 310 0 350 10
rect 600 0 680 10
rect 730 0 910 10
rect 4400 0 4580 10
rect 5340 0 5360 10
rect 5400 0 5640 10
rect 5860 0 5930 10
rect 5940 0 6090 10
rect 6440 0 6490 10
rect 6900 0 7160 10
rect 7290 0 7350 10
rect 8590 0 8600 10
rect 8680 0 8690 10
rect 9010 0 9020 10
rect 9180 0 9190 10
rect 9680 0 9710 10
<< metal2 >>
rect 2180 7490 2190 7500
rect 3740 7490 3750 7500
rect 3770 7490 3790 7500
rect 9760 7490 9810 7500
rect 2170 7480 2180 7490
rect 3780 7480 3800 7490
rect 9760 7480 9810 7490
rect 2160 7470 2170 7480
rect 3670 7470 3680 7480
rect 3740 7470 3760 7480
rect 3780 7470 3810 7480
rect 9680 7470 9690 7480
rect 9760 7470 9800 7480
rect 2150 7460 2170 7470
rect 3790 7460 3810 7470
rect 9640 7460 9670 7470
rect 9680 7460 9690 7470
rect 9760 7460 9800 7470
rect 2140 7450 2160 7460
rect 3790 7450 3820 7460
rect 9640 7450 9680 7460
rect 9750 7450 9800 7460
rect 9850 7450 9860 7460
rect 2130 7440 2160 7450
rect 3560 7440 3570 7450
rect 3790 7440 3820 7450
rect 9640 7440 9720 7450
rect 9730 7440 9780 7450
rect 9970 7440 9990 7450
rect 2110 7430 2150 7440
rect 3800 7430 3830 7440
rect 9640 7430 9770 7440
rect 9970 7430 9990 7440
rect 2110 7420 2140 7430
rect 3570 7420 3580 7430
rect 3810 7420 3830 7430
rect 9640 7420 9750 7430
rect 9950 7420 9990 7430
rect 2100 7410 2120 7420
rect 3640 7410 3650 7420
rect 3820 7410 3840 7420
rect 9640 7410 9690 7420
rect 9940 7410 9990 7420
rect 2090 7400 2110 7410
rect 3590 7400 3600 7410
rect 3640 7400 3650 7410
rect 3830 7400 3850 7410
rect 9640 7400 9670 7410
rect 9930 7400 9990 7410
rect 2090 7390 2110 7400
rect 3330 7390 3340 7400
rect 3840 7390 3850 7400
rect 9640 7390 9650 7400
rect 9930 7390 9990 7400
rect 2070 7380 2100 7390
rect 3620 7380 3630 7390
rect 3840 7380 3850 7390
rect 9940 7380 9970 7390
rect 3850 7370 3860 7380
rect 2050 7360 2080 7370
rect 3850 7360 3860 7370
rect 3350 7350 3360 7360
rect 3860 7350 3870 7360
rect 9630 7350 9640 7360
rect 2040 7340 2070 7350
rect 9630 7340 9640 7350
rect 2040 7330 2060 7340
rect 9620 7330 9640 7340
rect 9850 7330 9860 7340
rect 9980 7330 9990 7340
rect 2020 7320 2060 7330
rect 9630 7320 9640 7330
rect 9980 7320 9990 7330
rect 2020 7310 2050 7320
rect 9640 7310 9650 7320
rect 9960 7310 9990 7320
rect 2030 7300 2040 7310
rect 9640 7300 9660 7310
rect 9700 7300 9730 7310
rect 9940 7300 9990 7310
rect 2030 7290 2040 7300
rect 3360 7290 3370 7300
rect 3830 7290 3840 7300
rect 9640 7290 9670 7300
rect 9690 7290 9740 7300
rect 9780 7290 9840 7300
rect 9980 7290 9990 7300
rect 2010 7280 2020 7290
rect 3360 7280 3370 7290
rect 9560 7280 9570 7290
rect 9640 7280 9670 7290
rect 9690 7280 9850 7290
rect 9980 7280 9990 7290
rect 2010 7270 2020 7280
rect 9650 7270 9850 7280
rect 9970 7270 9990 7280
rect 1990 7260 2020 7270
rect 3380 7260 3390 7270
rect 3400 7260 3410 7270
rect 3840 7260 3850 7270
rect 3860 7260 3870 7270
rect 9640 7260 9850 7270
rect 9970 7260 9990 7270
rect 1990 7250 2010 7260
rect 3370 7250 3380 7260
rect 3400 7250 3410 7260
rect 3860 7250 3870 7260
rect 9650 7250 9760 7260
rect 9780 7250 9850 7260
rect 9960 7250 9990 7260
rect 1980 7240 2000 7250
rect 3370 7240 3380 7250
rect 9570 7240 9580 7250
rect 9640 7240 9750 7250
rect 9780 7240 9860 7250
rect 9950 7240 9990 7250
rect 1980 7230 2000 7240
rect 3410 7230 3420 7240
rect 3860 7230 3870 7240
rect 9650 7230 9750 7240
rect 9770 7230 9850 7240
rect 9950 7230 9990 7240
rect 1980 7220 1990 7230
rect 3380 7220 3390 7230
rect 3850 7220 3870 7230
rect 9610 7220 9620 7230
rect 9640 7220 9850 7230
rect 9950 7220 9990 7230
rect 1970 7210 1980 7220
rect 3440 7210 3450 7220
rect 3880 7210 3890 7220
rect 3900 7210 3910 7220
rect 9610 7210 9840 7220
rect 9950 7210 9990 7220
rect 1970 7200 1980 7210
rect 3870 7200 3910 7210
rect 9620 7200 9830 7210
rect 9960 7200 9990 7210
rect 1960 7190 1980 7200
rect 3870 7190 3920 7200
rect 9610 7190 9830 7200
rect 9970 7190 9990 7200
rect 1950 7180 1960 7190
rect 1970 7180 1980 7190
rect 3400 7180 3410 7190
rect 3860 7180 3920 7190
rect 9600 7180 9830 7190
rect 9970 7180 9990 7190
rect 1940 7170 1970 7180
rect 3440 7170 3450 7180
rect 3740 7170 3750 7180
rect 3880 7170 3920 7180
rect 9600 7170 9830 7180
rect 9970 7170 9990 7180
rect 1930 7160 1960 7170
rect 3730 7160 3750 7170
rect 3820 7160 3830 7170
rect 3880 7160 3930 7170
rect 9600 7160 9700 7170
rect 9710 7160 9830 7170
rect 9970 7160 9980 7170
rect 1930 7150 1950 7160
rect 3500 7150 3530 7160
rect 3690 7150 3700 7160
rect 3730 7150 3750 7160
rect 3820 7150 3850 7160
rect 3880 7150 3930 7160
rect 9600 7150 9690 7160
rect 9710 7150 9820 7160
rect 9860 7150 9870 7160
rect 9970 7150 9980 7160
rect 1920 7140 1950 7150
rect 3490 7140 3500 7150
rect 3530 7140 3540 7150
rect 3680 7140 3690 7150
rect 3740 7140 3750 7150
rect 3820 7140 3830 7150
rect 3880 7140 3930 7150
rect 9590 7140 9700 7150
rect 9720 7140 9820 7150
rect 9970 7140 9990 7150
rect 1920 7130 1950 7140
rect 2150 7130 2160 7140
rect 3500 7130 3510 7140
rect 3660 7130 3670 7140
rect 3820 7130 3840 7140
rect 3880 7130 3930 7140
rect 6610 7130 6620 7140
rect 9590 7130 9700 7140
rect 9720 7130 9820 7140
rect 9970 7130 9990 7140
rect 1930 7120 1940 7130
rect 2140 7120 2150 7130
rect 3410 7120 3420 7130
rect 3430 7120 3450 7130
rect 3650 7120 3660 7130
rect 3700 7120 3710 7130
rect 3770 7120 3780 7130
rect 3820 7120 3840 7130
rect 3870 7120 3930 7130
rect 6590 7120 6620 7130
rect 9590 7120 9680 7130
rect 9730 7120 9820 7130
rect 9970 7120 9990 7130
rect 1920 7110 1930 7120
rect 2140 7110 2160 7120
rect 3460 7110 3470 7120
rect 3640 7110 3660 7120
rect 3710 7110 3720 7120
rect 3770 7110 3790 7120
rect 3820 7110 3830 7120
rect 3870 7110 3930 7120
rect 6580 7110 6620 7120
rect 9580 7110 9660 7120
rect 9730 7110 9820 7120
rect 9970 7110 9990 7120
rect 1920 7100 1930 7110
rect 2120 7100 2150 7110
rect 3470 7100 3480 7110
rect 3520 7100 3530 7110
rect 3730 7100 3790 7110
rect 3820 7100 3830 7110
rect 3870 7100 3930 7110
rect 6570 7100 6620 7110
rect 9570 7100 9670 7110
rect 9730 7100 9810 7110
rect 1910 7090 1930 7100
rect 2080 7090 2090 7100
rect 2110 7090 2130 7100
rect 3480 7090 3490 7100
rect 3520 7090 3530 7100
rect 3560 7090 3570 7100
rect 3700 7090 3740 7100
rect 3760 7090 3800 7100
rect 3820 7090 3830 7100
rect 3870 7090 3930 7100
rect 6570 7090 6620 7100
rect 9570 7090 9670 7100
rect 9740 7090 9800 7100
rect 1910 7080 1930 7090
rect 1990 7080 2020 7090
rect 2060 7080 2120 7090
rect 3490 7080 3500 7090
rect 3530 7080 3540 7090
rect 3550 7080 3580 7090
rect 3700 7080 3730 7090
rect 3750 7080 3790 7090
rect 3820 7080 3840 7090
rect 3860 7080 3940 7090
rect 6560 7080 6610 7090
rect 9570 7080 9590 7090
rect 9620 7080 9670 7090
rect 9740 7080 9800 7090
rect 1900 7070 1930 7080
rect 2050 7070 2070 7080
rect 2090 7070 2110 7080
rect 3500 7070 3510 7080
rect 3540 7070 3550 7080
rect 3560 7070 3580 7080
rect 3620 7070 3630 7080
rect 3690 7070 3710 7080
rect 3730 7070 3740 7080
rect 3770 7070 3790 7080
rect 3820 7070 3830 7080
rect 3870 7070 3940 7080
rect 6550 7070 6610 7080
rect 9570 7070 9580 7080
rect 9620 7070 9680 7080
rect 9740 7070 9780 7080
rect 1910 7060 1930 7070
rect 2010 7060 2020 7070
rect 2030 7060 2060 7070
rect 2090 7060 2100 7070
rect 3510 7060 3520 7070
rect 3620 7060 3630 7070
rect 3690 7060 3710 7070
rect 3740 7060 3750 7070
rect 3780 7060 3790 7070
rect 3820 7060 3850 7070
rect 3860 7060 3940 7070
rect 6560 7060 6600 7070
rect 9610 7060 9680 7070
rect 9750 7060 9770 7070
rect 1910 7050 1930 7060
rect 2010 7050 2050 7060
rect 2070 7050 2090 7060
rect 3580 7050 3590 7060
rect 3690 7050 3710 7060
rect 3740 7050 3750 7060
rect 3770 7050 3790 7060
rect 3820 7050 3850 7060
rect 3860 7050 3940 7060
rect 9570 7050 9580 7060
rect 9600 7050 9680 7060
rect 1900 7040 1930 7050
rect 1950 7040 1980 7050
rect 2010 7040 2020 7050
rect 2260 7040 2290 7050
rect 3690 7040 3700 7050
rect 3710 7040 3720 7050
rect 3750 7040 3780 7050
rect 3820 7040 3940 7050
rect 9570 7040 9680 7050
rect 1900 7030 1930 7040
rect 1940 7030 1950 7040
rect 1970 7030 1980 7040
rect 2020 7030 2030 7040
rect 2050 7030 2070 7040
rect 2260 7030 2300 7040
rect 2340 7030 2350 7040
rect 2360 7030 2370 7040
rect 3630 7030 3650 7040
rect 3720 7030 3730 7040
rect 3770 7030 3780 7040
rect 3830 7030 3940 7040
rect 9580 7030 9670 7040
rect 1900 7020 1930 7030
rect 2000 7020 2030 7030
rect 2050 7020 2060 7030
rect 2240 7020 2410 7030
rect 3010 7020 3070 7030
rect 3630 7020 3640 7030
rect 3700 7020 3710 7030
rect 3770 7020 3780 7030
rect 3810 7020 3820 7030
rect 3830 7020 3940 7030
rect 9580 7020 9670 7030
rect 1910 7010 1920 7020
rect 2000 7010 2050 7020
rect 2260 7010 2420 7020
rect 2880 7010 2900 7020
rect 2980 7010 3120 7020
rect 3640 7010 3650 7020
rect 3700 7010 3730 7020
rect 3810 7010 3930 7020
rect 9580 7010 9670 7020
rect 1970 7000 2000 7010
rect 2260 7000 2440 7010
rect 2560 7000 2580 7010
rect 2720 7000 2730 7010
rect 2780 7000 2800 7010
rect 2820 7000 2930 7010
rect 2980 7000 3170 7010
rect 3710 7000 3730 7010
rect 3810 7000 3930 7010
rect 9600 7000 9670 7010
rect 1890 6990 1910 7000
rect 1950 6990 1980 7000
rect 2010 6990 2020 7000
rect 2260 6990 2450 7000
rect 2500 6990 2510 7000
rect 2560 6990 2590 7000
rect 2640 6990 2660 7000
rect 2720 6990 2750 7000
rect 2780 6990 3150 7000
rect 3160 6990 3170 7000
rect 3190 6990 3200 7000
rect 3610 6990 3620 7000
rect 3670 6990 3680 7000
rect 3720 6990 3730 7000
rect 3820 6990 3930 7000
rect 9610 6990 9670 7000
rect 1950 6980 1980 6990
rect 1990 6980 2000 6990
rect 2270 6980 2470 6990
rect 2510 6980 2520 6990
rect 2580 6980 2610 6990
rect 2640 6980 2690 6990
rect 2720 6980 2970 6990
rect 2980 6980 3160 6990
rect 3170 6980 3180 6990
rect 3230 6980 3240 6990
rect 3700 6980 3730 6990
rect 3830 6980 3910 6990
rect 9610 6980 9670 6990
rect 1970 6970 1990 6980
rect 2280 6970 2490 6980
rect 2520 6970 2540 6980
rect 2580 6970 2630 6980
rect 2660 6970 3170 6980
rect 3260 6970 3270 6980
rect 3640 6970 3650 6980
rect 3840 6970 3910 6980
rect 9610 6970 9670 6980
rect 9770 6970 9780 6980
rect 1940 6960 1950 6970
rect 1970 6960 1980 6970
rect 2270 6960 2490 6970
rect 2530 6960 2560 6970
rect 2600 6960 2640 6970
rect 2660 6960 3170 6970
rect 3290 6960 3300 6970
rect 3660 6960 3670 6970
rect 3850 6960 3910 6970
rect 9610 6960 9660 6970
rect 9750 6960 9780 6970
rect 9790 6960 9800 6970
rect 9810 6960 9820 6970
rect 1940 6950 1950 6960
rect 2300 6950 2450 6960
rect 2460 6950 2480 6960
rect 2490 6950 2500 6960
rect 2540 6950 2580 6960
rect 2610 6950 3180 6960
rect 3310 6950 3320 6960
rect 3680 6950 3700 6960
rect 3860 6950 3910 6960
rect 9620 6950 9650 6960
rect 9740 6950 9790 6960
rect 1940 6940 1950 6950
rect 2310 6940 2440 6950
rect 2460 6940 2470 6950
rect 2500 6940 2520 6950
rect 2560 6940 2600 6950
rect 2610 6940 3180 6950
rect 3340 6940 3350 6950
rect 3720 6940 3780 6950
rect 3870 6940 3910 6950
rect 9630 6940 9650 6950
rect 9720 6940 9770 6950
rect 2310 6930 2450 6940
rect 2520 6930 2540 6940
rect 2580 6930 2700 6940
rect 2710 6930 3190 6940
rect 3370 6930 3380 6940
rect 3730 6930 3790 6940
rect 3870 6930 3910 6940
rect 9630 6930 9650 6940
rect 9710 6930 9750 6940
rect 1920 6920 1930 6930
rect 2330 6920 2470 6930
rect 2480 6920 2490 6930
rect 2540 6920 2550 6930
rect 2580 6920 2720 6930
rect 2730 6920 3200 6930
rect 3740 6920 3780 6930
rect 3790 6920 3810 6930
rect 3870 6920 3890 6930
rect 9630 6920 9650 6930
rect 9690 6920 9700 6930
rect 1890 6910 1920 6920
rect 2360 6910 2480 6920
rect 2560 6910 2580 6920
rect 2590 6910 2890 6920
rect 2900 6910 3040 6920
rect 3060 6910 3090 6920
rect 3100 6910 3220 6920
rect 3420 6910 3430 6920
rect 3740 6910 3790 6920
rect 3800 6910 3810 6920
rect 3870 6910 3890 6920
rect 9610 6910 9650 6920
rect 9680 6910 9700 6920
rect 1890 6900 1900 6910
rect 2360 6900 2510 6910
rect 2580 6900 2680 6910
rect 2690 6900 2910 6910
rect 2920 6900 3030 6910
rect 3060 6900 3100 6910
rect 3120 6900 3230 6910
rect 3760 6900 3820 6910
rect 3870 6900 3900 6910
rect 9590 6900 9680 6910
rect 1880 6890 1890 6900
rect 2380 6890 2510 6900
rect 2600 6890 2700 6900
rect 2710 6890 2830 6900
rect 2850 6890 2920 6900
rect 2950 6890 3000 6900
rect 3020 6890 3070 6900
rect 3090 6890 3120 6900
rect 3140 6890 3230 6900
rect 3770 6890 3810 6900
rect 3820 6890 3840 6900
rect 3880 6890 3900 6900
rect 9590 6890 9680 6900
rect 1880 6880 1890 6890
rect 2410 6880 2520 6890
rect 2610 6880 2880 6890
rect 2890 6880 2940 6890
rect 2990 6880 3110 6890
rect 3120 6880 3160 6890
rect 3170 6880 3240 6890
rect 3250 6880 3260 6890
rect 3780 6880 3850 6890
rect 3870 6880 3880 6890
rect 3890 6880 3900 6890
rect 9590 6880 9680 6890
rect 1880 6870 1900 6880
rect 2420 6870 2520 6880
rect 2640 6870 2710 6880
rect 2740 6870 2890 6880
rect 2940 6870 2980 6880
rect 3020 6870 3030 6880
rect 3040 6870 3070 6880
rect 3080 6870 3090 6880
rect 3120 6870 3160 6880
rect 3250 6870 3260 6880
rect 3780 6870 3880 6880
rect 9590 6870 9680 6880
rect 1910 6860 1920 6870
rect 2440 6860 2540 6870
rect 2670 6860 2720 6870
rect 2750 6860 2840 6870
rect 2850 6860 2920 6870
rect 2970 6860 2990 6870
rect 3060 6860 3080 6870
rect 3130 6860 3150 6870
rect 3790 6860 3880 6870
rect 9590 6860 9680 6870
rect 1900 6850 1910 6860
rect 2470 6850 2560 6860
rect 2690 6850 2720 6860
rect 2730 6850 2750 6860
rect 2770 6850 2910 6860
rect 2920 6850 2960 6860
rect 2970 6850 3050 6860
rect 3810 6850 3830 6860
rect 3880 6850 3890 6860
rect 9590 6850 9680 6860
rect 2490 6840 2560 6850
rect 2730 6840 2900 6850
rect 2950 6840 3040 6850
rect 3060 6840 3070 6850
rect 3820 6840 3840 6850
rect 9590 6840 9680 6850
rect 1890 6830 1900 6840
rect 2500 6830 2590 6840
rect 2780 6830 2940 6840
rect 2950 6830 3070 6840
rect 3120 6830 3130 6840
rect 3820 6830 3890 6840
rect 9590 6830 9680 6840
rect 2510 6820 2620 6830
rect 2830 6820 2870 6830
rect 2920 6820 2990 6830
rect 3020 6820 3080 6830
rect 3140 6820 3160 6830
rect 3600 6820 3610 6830
rect 3830 6820 3890 6830
rect 9590 6820 9680 6830
rect 2550 6810 2690 6820
rect 2900 6810 2930 6820
rect 3000 6810 3010 6820
rect 3040 6810 3060 6820
rect 3830 6810 3890 6820
rect 9590 6810 9630 6820
rect 9640 6810 9680 6820
rect 1850 6800 1860 6810
rect 2560 6800 2570 6810
rect 2580 6800 2740 6810
rect 3830 6800 3900 6810
rect 9590 6800 9680 6810
rect 1870 6790 1880 6800
rect 2680 6790 2790 6800
rect 3840 6790 3900 6800
rect 9600 6790 9620 6800
rect 9640 6790 9680 6800
rect 1970 6780 2010 6790
rect 2710 6780 2830 6790
rect 3850 6780 3910 6790
rect 9600 6780 9610 6790
rect 9650 6780 9680 6790
rect 1870 6770 1890 6780
rect 1990 6770 2000 6780
rect 2300 6770 2380 6780
rect 2730 6770 2750 6780
rect 2800 6770 2880 6780
rect 3720 6770 3730 6780
rect 3850 6770 3900 6780
rect 3910 6770 3920 6780
rect 9650 6770 9680 6780
rect 1870 6760 1890 6770
rect 1960 6760 1970 6770
rect 1980 6760 1990 6770
rect 2290 6760 2400 6770
rect 2860 6760 2980 6770
rect 3850 6760 3920 6770
rect 9640 6760 9690 6770
rect 1950 6750 1960 6760
rect 1980 6750 1990 6760
rect 2280 6750 2400 6760
rect 2920 6750 3060 6760
rect 3850 6750 3920 6760
rect 9570 6750 9580 6760
rect 9640 6750 9690 6760
rect 1870 6740 1880 6750
rect 1950 6740 1970 6750
rect 2260 6740 2360 6750
rect 3030 6740 3140 6750
rect 3870 6740 3930 6750
rect 9550 6740 9580 6750
rect 9640 6740 9690 6750
rect 1930 6730 1980 6740
rect 2260 6730 2340 6740
rect 2460 6730 2470 6740
rect 3080 6730 3110 6740
rect 3120 6730 3230 6740
rect 3870 6730 3930 6740
rect 9560 6730 9570 6740
rect 9640 6730 9690 6740
rect 1870 6720 1890 6730
rect 2240 6720 2310 6730
rect 2480 6720 2490 6730
rect 3150 6720 3190 6730
rect 3200 6720 3260 6730
rect 3750 6720 3760 6730
rect 3780 6720 3790 6730
rect 3880 6720 3940 6730
rect 9640 6720 9690 6730
rect 1840 6710 1850 6720
rect 1860 6710 1870 6720
rect 1880 6710 1890 6720
rect 2240 6710 2300 6720
rect 2500 6710 2510 6720
rect 3240 6710 3310 6720
rect 3320 6710 3330 6720
rect 3890 6710 3940 6720
rect 9640 6710 9690 6720
rect 1870 6700 1880 6710
rect 2240 6700 2290 6710
rect 2500 6700 2540 6710
rect 3290 6700 3360 6710
rect 3900 6700 3940 6710
rect 9530 6700 9540 6710
rect 9640 6700 9690 6710
rect 1860 6690 1870 6700
rect 2250 6690 2270 6700
rect 2510 6690 2540 6700
rect 2560 6690 2570 6700
rect 3350 6690 3420 6700
rect 3910 6690 3940 6700
rect 9560 6690 9570 6700
rect 9640 6690 9690 6700
rect 9990 6690 9990 6700
rect 1800 6680 1830 6690
rect 1840 6680 1860 6690
rect 1890 6680 1910 6690
rect 2250 6680 2260 6690
rect 2520 6680 2580 6690
rect 3410 6680 3440 6690
rect 3820 6680 3830 6690
rect 3910 6680 3930 6690
rect 9550 6680 9570 6690
rect 9600 6680 9610 6690
rect 9640 6680 9690 6690
rect 9970 6680 9980 6690
rect 1840 6670 1850 6680
rect 1900 6670 1910 6680
rect 2240 6670 2250 6680
rect 2550 6670 2580 6680
rect 3430 6670 3470 6680
rect 3810 6670 3820 6680
rect 3830 6670 3840 6680
rect 3910 6670 3950 6680
rect 9510 6670 9520 6680
rect 9540 6670 9550 6680
rect 9600 6670 9610 6680
rect 9650 6670 9690 6680
rect 9940 6670 9950 6680
rect 1870 6660 1880 6670
rect 2240 6660 2250 6670
rect 2550 6660 2580 6670
rect 3480 6660 3490 6670
rect 3920 6660 3950 6670
rect 9500 6660 9510 6670
rect 9530 6660 9550 6670
rect 9650 6660 9690 6670
rect 1850 6650 1880 6660
rect 2230 6650 2240 6660
rect 2560 6650 2590 6660
rect 3500 6650 3550 6660
rect 3930 6650 3960 6660
rect 9510 6650 9540 6660
rect 9640 6650 9690 6660
rect 9870 6650 9890 6660
rect 1840 6640 1850 6650
rect 2220 6640 2230 6650
rect 2560 6640 2600 6650
rect 3530 6640 3570 6650
rect 3860 6640 3870 6650
rect 3940 6640 3960 6650
rect 9490 6640 9500 6650
rect 9520 6640 9540 6650
rect 9610 6640 9620 6650
rect 9650 6640 9690 6650
rect 9840 6640 9850 6650
rect 1760 6630 1820 6640
rect 1850 6630 1860 6640
rect 2210 6630 2220 6640
rect 2570 6630 2600 6640
rect 3550 6630 3610 6640
rect 3940 6630 3970 6640
rect 9520 6630 9540 6640
rect 9610 6630 9620 6640
rect 9650 6630 9700 6640
rect 9810 6630 9820 6640
rect 1740 6620 1750 6630
rect 2210 6620 2220 6630
rect 2570 6620 2610 6630
rect 3600 6620 3630 6630
rect 3950 6620 3970 6630
rect 9500 6620 9520 6630
rect 9610 6620 9620 6630
rect 9630 6620 9640 6630
rect 9650 6620 9690 6630
rect 9780 6620 9790 6630
rect 2190 6610 2220 6620
rect 2580 6610 2620 6620
rect 3620 6610 3650 6620
rect 3950 6610 3970 6620
rect 9480 6610 9490 6620
rect 9500 6610 9520 6620
rect 9610 6610 9630 6620
rect 9640 6610 9690 6620
rect 9750 6610 9760 6620
rect 1600 6600 1610 6610
rect 2180 6600 2210 6610
rect 2580 6600 2610 6610
rect 3640 6600 3680 6610
rect 3960 6600 3970 6610
rect 9480 6600 9490 6610
rect 9510 6600 9520 6610
rect 9610 6600 9630 6610
rect 9640 6600 9700 6610
rect 9720 6600 9730 6610
rect 1590 6590 1600 6600
rect 2180 6590 2200 6600
rect 2590 6590 2620 6600
rect 3680 6590 3690 6600
rect 3960 6590 3980 6600
rect 6080 6590 6090 6600
rect 9480 6590 9490 6600
rect 9510 6590 9520 6600
rect 9610 6590 9680 6600
rect 1570 6580 1580 6590
rect 1610 6580 1620 6590
rect 1630 6580 1640 6590
rect 1770 6580 1780 6590
rect 2070 6580 2090 6590
rect 2170 6580 2190 6590
rect 2590 6580 2620 6590
rect 3700 6580 3730 6590
rect 3960 6580 3990 6590
rect 6080 6580 6090 6590
rect 9500 6580 9530 6590
rect 9610 6580 9670 6590
rect 1550 6570 1560 6580
rect 1780 6570 1790 6580
rect 2120 6570 2130 6580
rect 2170 6570 2190 6580
rect 2600 6570 2620 6580
rect 3720 6570 3740 6580
rect 3970 6570 4000 6580
rect 6270 6570 6280 6580
rect 9490 6570 9520 6580
rect 9630 6570 9640 6580
rect 1360 6560 1370 6570
rect 1540 6560 1550 6570
rect 1590 6560 1610 6570
rect 1790 6560 1800 6570
rect 2000 6560 2020 6570
rect 2040 6560 2050 6570
rect 2600 6560 2620 6570
rect 3740 6560 3760 6570
rect 3920 6560 3930 6570
rect 3980 6560 4000 6570
rect 6010 6560 6020 6570
rect 6220 6560 6230 6570
rect 6260 6560 6270 6570
rect 9500 6560 9520 6570
rect 1360 6550 1380 6560
rect 1590 6550 1610 6560
rect 1620 6550 1630 6560
rect 1780 6550 1810 6560
rect 2030 6550 2040 6560
rect 2590 6550 2620 6560
rect 3760 6550 3780 6560
rect 3990 6550 4000 6560
rect 6010 6550 6030 6560
rect 6220 6550 6240 6560
rect 9500 6550 9510 6560
rect 1360 6540 1390 6550
rect 1460 6540 1490 6550
rect 1590 6540 1630 6550
rect 1730 6540 1750 6550
rect 1800 6540 1820 6550
rect 2010 6540 2050 6550
rect 2600 6540 2630 6550
rect 3770 6540 3790 6550
rect 5970 6540 5980 6550
rect 6030 6540 6040 6550
rect 6060 6540 6070 6550
rect 6220 6540 6240 6550
rect 6250 6540 6270 6550
rect 6360 6540 6380 6550
rect 6420 6540 6450 6550
rect 6540 6540 6560 6550
rect 1440 6530 1450 6540
rect 1480 6530 1500 6540
rect 1750 6530 1760 6540
rect 1800 6530 1830 6540
rect 2580 6530 2630 6540
rect 3800 6530 3820 6540
rect 4000 6530 4010 6540
rect 6030 6530 6050 6540
rect 6220 6530 6240 6540
rect 6250 6530 6270 6540
rect 6350 6530 6460 6540
rect 6480 6530 6490 6540
rect 6510 6530 6570 6540
rect 1420 6520 1440 6530
rect 1770 6520 1780 6530
rect 1800 6520 1840 6530
rect 2570 6520 2580 6530
rect 3820 6520 3840 6530
rect 4000 6520 4010 6530
rect 6000 6520 6020 6530
rect 6040 6520 6050 6530
rect 6060 6520 6080 6530
rect 6230 6520 6240 6530
rect 6260 6520 6280 6530
rect 6310 6520 6340 6530
rect 6360 6520 6450 6530
rect 6460 6520 6560 6530
rect 6620 6520 6630 6530
rect 9420 6520 9430 6530
rect 9980 6520 9990 6530
rect 1320 6510 1370 6520
rect 1430 6510 1480 6520
rect 1780 6510 1840 6520
rect 2540 6510 2550 6520
rect 3840 6510 3850 6520
rect 4000 6510 4010 6520
rect 6010 6510 6030 6520
rect 6050 6510 6080 6520
rect 6170 6510 6210 6520
rect 6270 6510 6280 6520
rect 6310 6510 6380 6520
rect 6390 6510 6520 6520
rect 6530 6510 6560 6520
rect 6580 6510 6630 6520
rect 9420 6510 9440 6520
rect 9950 6510 9970 6520
rect 1300 6500 1310 6510
rect 1790 6500 1850 6510
rect 2090 6500 2100 6510
rect 2250 6500 2270 6510
rect 2420 6500 2440 6510
rect 2500 6500 2520 6510
rect 3860 6500 3870 6510
rect 4000 6500 4010 6510
rect 6000 6500 6010 6510
rect 6020 6500 6030 6510
rect 6060 6500 6090 6510
rect 6110 6500 6240 6510
rect 6270 6500 6310 6510
rect 6330 6500 6380 6510
rect 6430 6500 6480 6510
rect 6540 6500 6600 6510
rect 6610 6500 6620 6510
rect 9910 6500 9940 6510
rect 1260 6490 1270 6500
rect 1800 6490 1850 6500
rect 2110 6490 2120 6500
rect 2260 6490 2270 6500
rect 2400 6490 2410 6500
rect 2440 6490 2480 6500
rect 4010 6490 4020 6500
rect 5810 6490 5820 6500
rect 6070 6490 6240 6500
rect 6250 6490 6320 6500
rect 6340 6490 6380 6500
rect 6430 6490 6450 6500
rect 6540 6490 6610 6500
rect 9880 6490 9890 6500
rect 1250 6480 1260 6490
rect 1270 6480 1280 6490
rect 1710 6480 1760 6490
rect 1800 6480 1810 6490
rect 1820 6480 1840 6490
rect 2120 6480 2130 6490
rect 2260 6480 2280 6490
rect 2400 6480 2410 6490
rect 2470 6480 2480 6490
rect 3980 6480 3990 6490
rect 4010 6480 4020 6490
rect 6080 6480 6340 6490
rect 6360 6480 6390 6490
rect 6540 6480 6620 6490
rect 9860 6480 9870 6490
rect 1240 6470 1270 6480
rect 1340 6470 1370 6480
rect 1690 6470 1770 6480
rect 1830 6470 1850 6480
rect 2130 6470 2150 6480
rect 2540 6470 2560 6480
rect 3910 6470 3920 6480
rect 6090 6470 6350 6480
rect 6360 6470 6400 6480
rect 6530 6470 6610 6480
rect 9810 6470 9850 6480
rect 1240 6460 1250 6470
rect 1330 6460 1360 6470
rect 1370 6460 1380 6470
rect 1680 6460 1690 6470
rect 1720 6460 1770 6470
rect 1810 6460 1820 6470
rect 1830 6460 1860 6470
rect 2390 6460 2400 6470
rect 4000 6460 4010 6470
rect 4020 6460 4030 6470
rect 6100 6460 6140 6470
rect 6150 6460 6160 6470
rect 6170 6460 6400 6470
rect 6520 6460 6590 6470
rect 9770 6460 9780 6470
rect 1300 6450 1360 6460
rect 1660 6450 1670 6460
rect 1730 6450 1770 6460
rect 1810 6450 1820 6460
rect 1830 6450 1890 6460
rect 1900 6450 1940 6460
rect 2100 6450 2120 6460
rect 2290 6450 2300 6460
rect 3940 6450 3950 6460
rect 4030 6450 4040 6460
rect 6100 6450 6120 6460
rect 6190 6450 6410 6460
rect 6530 6450 6540 6460
rect 6570 6450 6600 6460
rect 9740 6450 9750 6460
rect 1240 6440 1250 6450
rect 1290 6440 1300 6450
rect 1340 6440 1380 6450
rect 1650 6440 1660 6450
rect 1740 6440 1770 6450
rect 1830 6440 1940 6450
rect 2080 6440 2120 6450
rect 2140 6440 2150 6450
rect 2260 6440 2270 6450
rect 2280 6440 2290 6450
rect 3960 6440 3970 6450
rect 6090 6440 6120 6450
rect 6210 6440 6310 6450
rect 6330 6440 6420 6450
rect 6570 6440 6610 6450
rect 6660 6440 6670 6450
rect 9680 6440 9700 6450
rect 1240 6430 1250 6440
rect 1350 6430 1370 6440
rect 1740 6430 1770 6440
rect 1810 6430 1820 6440
rect 1830 6430 1870 6440
rect 1890 6430 1920 6440
rect 1930 6430 1960 6440
rect 2100 6430 2130 6440
rect 2310 6430 2330 6440
rect 3970 6430 3980 6440
rect 5810 6430 5970 6440
rect 6080 6430 6120 6440
rect 6210 6430 6220 6440
rect 6230 6430 6280 6440
rect 6290 6430 6320 6440
rect 6340 6430 6420 6440
rect 6590 6430 6630 6440
rect 6670 6430 6680 6440
rect 9670 6430 9680 6440
rect 9950 6430 9970 6440
rect 1280 6420 1290 6430
rect 1330 6420 1370 6430
rect 1640 6420 1650 6430
rect 1740 6420 1790 6430
rect 1830 6420 1870 6430
rect 1940 6420 1960 6430
rect 2070 6420 2080 6430
rect 2090 6420 2110 6430
rect 2320 6420 2330 6430
rect 2500 6420 2510 6430
rect 3990 6420 4000 6430
rect 5810 6420 5840 6430
rect 5870 6420 5960 6430
rect 6100 6420 6110 6430
rect 6220 6420 6230 6430
rect 6240 6420 6260 6430
rect 6290 6420 6340 6430
rect 6350 6420 6370 6430
rect 6570 6420 6640 6430
rect 6690 6420 6700 6430
rect 9650 6420 9660 6430
rect 9940 6420 9980 6430
rect 1270 6410 1280 6420
rect 1330 6410 1370 6420
rect 1440 6410 1450 6420
rect 1460 6410 1470 6420
rect 1840 6410 1850 6420
rect 1940 6410 1970 6420
rect 2040 6410 2060 6420
rect 2500 6410 2510 6420
rect 5820 6410 5880 6420
rect 6100 6410 6120 6420
rect 6180 6410 6360 6420
rect 6550 6410 6560 6420
rect 6580 6410 6660 6420
rect 6690 6410 6720 6420
rect 8650 6410 8660 6420
rect 9640 6410 9650 6420
rect 9940 6410 9990 6420
rect 1230 6400 1240 6410
rect 1250 6400 1260 6410
rect 1320 6400 1370 6410
rect 1420 6400 1430 6410
rect 1480 6400 1490 6410
rect 1630 6400 1640 6410
rect 1940 6400 2060 6410
rect 4020 6400 4030 6410
rect 5760 6400 5770 6410
rect 5780 6400 5800 6410
rect 6050 6400 6090 6410
rect 6110 6400 6360 6410
rect 6590 6400 6670 6410
rect 6690 6400 6720 6410
rect 6770 6400 6780 6410
rect 9640 6400 9650 6410
rect 9940 6400 9990 6410
rect 1380 6390 1400 6400
rect 1450 6390 1460 6400
rect 1970 6390 2050 6400
rect 6070 6390 6090 6400
rect 6110 6390 6380 6400
rect 6590 6390 6780 6400
rect 9940 6390 9990 6400
rect 1240 6380 1250 6390
rect 1410 6380 1430 6390
rect 1620 6380 1630 6390
rect 1760 6380 1820 6390
rect 1970 6380 2010 6390
rect 4050 6380 4060 6390
rect 5890 6380 5930 6390
rect 5960 6380 6010 6390
rect 6120 6380 6280 6390
rect 6310 6380 6390 6390
rect 6600 6380 6800 6390
rect 9630 6380 9640 6390
rect 9940 6380 9990 6390
rect 1240 6370 1250 6380
rect 1390 6370 1430 6380
rect 1440 6370 1460 6380
rect 1610 6370 1620 6380
rect 1730 6370 1750 6380
rect 1830 6370 1840 6380
rect 2470 6370 2480 6380
rect 4060 6370 4070 6380
rect 5800 6370 5930 6380
rect 5960 6370 5990 6380
rect 6140 6370 6260 6380
rect 6350 6370 6380 6380
rect 6390 6370 6400 6380
rect 6600 6370 6800 6380
rect 9950 6370 9970 6380
rect 1230 6360 1240 6370
rect 1400 6360 1460 6370
rect 1710 6360 1740 6370
rect 1830 6360 1840 6370
rect 2400 6360 2410 6370
rect 5790 6360 5910 6370
rect 6350 6360 6410 6370
rect 6600 6360 6810 6370
rect 9780 6360 9790 6370
rect 1230 6350 1250 6360
rect 1410 6350 1460 6360
rect 1600 6350 1610 6360
rect 1680 6350 1720 6360
rect 2400 6350 2410 6360
rect 5750 6350 5880 6360
rect 6360 6350 6430 6360
rect 6610 6350 6830 6360
rect 9460 6350 9470 6360
rect 9780 6350 9800 6360
rect 1250 6340 1270 6350
rect 1410 6340 1430 6350
rect 1670 6340 1710 6350
rect 2410 6340 2420 6350
rect 2470 6340 2480 6350
rect 4100 6340 4110 6350
rect 5730 6340 5740 6350
rect 5780 6340 5820 6350
rect 6380 6340 6450 6350
rect 6670 6340 6810 6350
rect 9460 6340 9500 6350
rect 9630 6340 9640 6350
rect 9780 6340 9810 6350
rect 1410 6330 1430 6340
rect 1590 6330 1600 6340
rect 1660 6330 1710 6340
rect 2450 6330 2460 6340
rect 2470 6330 2480 6340
rect 4110 6330 4120 6340
rect 5560 6330 5670 6340
rect 5710 6330 5750 6340
rect 5790 6330 5820 6340
rect 6400 6330 6480 6340
rect 6500 6330 6510 6340
rect 6680 6330 6710 6340
rect 6720 6330 6810 6340
rect 9400 6330 9410 6340
rect 9460 6330 9480 6340
rect 9770 6330 9820 6340
rect 1220 6320 1250 6330
rect 1280 6320 1290 6330
rect 1410 6320 1420 6330
rect 1650 6320 1700 6330
rect 2400 6320 2410 6330
rect 4120 6320 4130 6330
rect 5480 6320 5500 6330
rect 5510 6320 5650 6330
rect 5690 6320 5710 6330
rect 5720 6320 5740 6330
rect 5790 6320 5820 6330
rect 6430 6320 6520 6330
rect 6700 6320 6720 6330
rect 6730 6320 6800 6330
rect 9400 6320 9410 6330
rect 9790 6320 9800 6330
rect 1240 6310 1270 6320
rect 1290 6310 1300 6320
rect 1410 6310 1420 6320
rect 1630 6310 1680 6320
rect 1830 6310 1840 6320
rect 2400 6310 2420 6320
rect 4130 6310 4140 6320
rect 5440 6310 5480 6320
rect 5500 6310 5630 6320
rect 5660 6310 5700 6320
rect 5720 6310 5760 6320
rect 5770 6310 5820 6320
rect 6440 6310 6540 6320
rect 6750 6310 6800 6320
rect 9330 6310 9340 6320
rect 9400 6310 9410 6320
rect 9490 6310 9510 6320
rect 1270 6300 1280 6310
rect 1300 6300 1310 6310
rect 1410 6300 1420 6310
rect 1580 6300 1590 6310
rect 1620 6300 1660 6310
rect 1830 6300 1840 6310
rect 2400 6300 2410 6310
rect 4140 6300 4150 6310
rect 5390 6300 5410 6310
rect 5500 6300 5520 6310
rect 5570 6300 5620 6310
rect 5640 6300 5660 6310
rect 5670 6300 5810 6310
rect 6460 6300 6560 6310
rect 6610 6300 6620 6310
rect 6750 6300 6770 6310
rect 9300 6300 9330 6310
rect 9410 6300 9420 6310
rect 9470 6300 9500 6310
rect 9980 6300 9990 6310
rect 1230 6290 1250 6300
rect 1270 6290 1290 6300
rect 1300 6290 1320 6300
rect 1400 6290 1410 6300
rect 1580 6290 1590 6300
rect 1620 6290 1640 6300
rect 2460 6290 2470 6300
rect 5370 6290 5410 6300
rect 5510 6290 5640 6300
rect 5670 6290 5710 6300
rect 6490 6290 6570 6300
rect 6770 6290 6780 6300
rect 8590 6290 8600 6300
rect 9400 6290 9420 6300
rect 9480 6290 9500 6300
rect 9590 6290 9610 6300
rect 9960 6290 9970 6300
rect 1230 6280 1270 6290
rect 1310 6280 1320 6290
rect 1580 6280 1590 6290
rect 1610 6280 1630 6290
rect 1820 6280 1830 6290
rect 2440 6280 2450 6290
rect 5380 6280 5400 6290
rect 5550 6280 5600 6290
rect 5620 6280 5680 6290
rect 6520 6280 6570 6290
rect 6610 6280 6620 6290
rect 6770 6280 6780 6290
rect 6800 6280 6820 6290
rect 9280 6280 9300 6290
rect 9400 6280 9410 6290
rect 9420 6280 9430 6290
rect 9480 6280 9500 6290
rect 9910 6280 9930 6290
rect 9950 6280 9960 6290
rect 1240 6270 1260 6280
rect 1310 6270 1330 6280
rect 1390 6270 1400 6280
rect 1580 6270 1590 6280
rect 1600 6270 1620 6280
rect 1820 6270 1830 6280
rect 2440 6270 2450 6280
rect 5360 6270 5370 6280
rect 5540 6270 5630 6280
rect 6530 6270 6580 6280
rect 6660 6270 6680 6280
rect 6770 6270 6830 6280
rect 8570 6270 8580 6280
rect 9280 6270 9320 6280
rect 9400 6270 9410 6280
rect 9480 6270 9500 6280
rect 9870 6270 9880 6280
rect 9890 6270 9940 6280
rect 9960 6270 9970 6280
rect 9980 6270 9990 6280
rect 1240 6260 1290 6270
rect 1320 6260 1330 6270
rect 1390 6260 1400 6270
rect 1540 6260 1550 6270
rect 1570 6260 1610 6270
rect 1810 6260 1820 6270
rect 2400 6260 2410 6270
rect 2440 6260 2450 6270
rect 5340 6260 5360 6270
rect 5530 6260 5620 6270
rect 6540 6260 6590 6270
rect 6650 6260 6680 6270
rect 6770 6260 6790 6270
rect 6810 6260 6840 6270
rect 8570 6260 8580 6270
rect 9270 6260 9320 6270
rect 9420 6260 9430 6270
rect 9480 6260 9500 6270
rect 9570 6260 9590 6270
rect 9850 6260 9870 6270
rect 9910 6260 9950 6270
rect 9990 6260 9990 6270
rect 1250 6250 1260 6260
rect 1320 6250 1340 6260
rect 1580 6250 1610 6260
rect 2440 6250 2450 6260
rect 5390 6250 5410 6260
rect 5520 6250 5610 6260
rect 6540 6250 6590 6260
rect 6650 6250 6660 6260
rect 6770 6250 6800 6260
rect 6810 6250 6850 6260
rect 9260 6250 9310 6260
rect 9410 6250 9420 6260
rect 9540 6250 9560 6260
rect 9640 6250 9650 6260
rect 9820 6250 9830 6260
rect 9860 6250 9870 6260
rect 9920 6250 9930 6260
rect 1230 6240 1260 6250
rect 1380 6240 1390 6250
rect 1570 6240 1600 6250
rect 1800 6240 1810 6250
rect 5310 6240 5330 6250
rect 5380 6240 5400 6250
rect 5520 6240 5590 6250
rect 6560 6240 6610 6250
rect 6650 6240 6660 6250
rect 6770 6240 6840 6250
rect 9260 6240 9300 6250
rect 9410 6240 9440 6250
rect 9510 6240 9520 6250
rect 1330 6230 1350 6240
rect 1380 6230 1390 6240
rect 1570 6230 1600 6240
rect 1790 6230 1800 6240
rect 5310 6230 5320 6240
rect 5510 6230 5580 6240
rect 6570 6230 6620 6240
rect 6630 6230 6650 6240
rect 6750 6230 6850 6240
rect 9250 6230 9260 6240
rect 9410 6230 9420 6240
rect 9480 6230 9490 6240
rect 9630 6230 9640 6240
rect 9650 6230 9660 6240
rect 1300 6220 1320 6230
rect 1330 6220 1360 6230
rect 1370 6220 1390 6230
rect 1570 6220 1600 6230
rect 1790 6220 1800 6230
rect 2450 6220 2460 6230
rect 5330 6220 5340 6230
rect 5500 6220 5550 6230
rect 6570 6220 6650 6230
rect 6750 6220 6780 6230
rect 6800 6220 6850 6230
rect 9250 6220 9290 6230
rect 9410 6220 9420 6230
rect 1280 6210 1290 6220
rect 1300 6210 1320 6220
rect 1330 6210 1340 6220
rect 1350 6210 1400 6220
rect 1580 6210 1610 6220
rect 1780 6210 1790 6220
rect 2450 6210 2460 6220
rect 4230 6210 4240 6220
rect 5290 6210 5300 6220
rect 5340 6210 5350 6220
rect 5480 6210 5540 6220
rect 6590 6210 6670 6220
rect 6760 6210 6780 6220
rect 6820 6210 6860 6220
rect 9240 6210 9290 6220
rect 9380 6210 9420 6220
rect 9630 6210 9640 6220
rect 9660 6210 9670 6220
rect 9800 6210 9810 6220
rect 9910 6210 9920 6220
rect 9940 6210 9950 6220
rect 1280 6200 1300 6210
rect 1360 6200 1370 6210
rect 1380 6200 1400 6210
rect 1580 6200 1620 6210
rect 1730 6200 1740 6210
rect 1760 6200 1780 6210
rect 5290 6200 5310 6210
rect 5320 6200 5350 6210
rect 5470 6200 5520 6210
rect 6610 6200 6670 6210
rect 6760 6200 6780 6210
rect 6840 6200 6870 6210
rect 9240 6200 9280 6210
rect 9310 6200 9320 6210
rect 9330 6200 9350 6210
rect 9800 6200 9810 6210
rect 1290 6190 1310 6200
rect 1320 6190 1330 6200
rect 1360 6190 1370 6200
rect 1380 6190 1400 6200
rect 1580 6190 1630 6200
rect 1720 6190 1780 6200
rect 5280 6190 5290 6200
rect 5310 6190 5320 6200
rect 5460 6190 5510 6200
rect 6630 6190 6670 6200
rect 6750 6190 6800 6200
rect 6830 6190 6880 6200
rect 9230 6190 9280 6200
rect 9310 6190 9360 6200
rect 9610 6190 9620 6200
rect 9800 6190 9820 6200
rect 1260 6180 1280 6190
rect 1290 6180 1310 6190
rect 1320 6180 1330 6190
rect 1340 6180 1350 6190
rect 1380 6180 1400 6190
rect 1590 6180 1630 6190
rect 1720 6180 1780 6190
rect 2390 6180 2400 6190
rect 2420 6180 2430 6190
rect 5300 6180 5310 6190
rect 5450 6180 5490 6190
rect 6650 6180 6680 6190
rect 6740 6180 6810 6190
rect 6820 6180 6890 6190
rect 7650 6180 7660 6190
rect 9220 6180 9230 6190
rect 9300 6180 9320 6190
rect 9610 6180 9620 6190
rect 9810 6180 9820 6190
rect 1260 6170 1280 6180
rect 1310 6170 1340 6180
rect 1370 6170 1400 6180
rect 1420 6170 1430 6180
rect 1590 6170 1600 6180
rect 1620 6170 1640 6180
rect 1720 6170 1780 6180
rect 2420 6170 2430 6180
rect 4260 6170 4270 6180
rect 5290 6170 5320 6180
rect 5440 6170 5470 6180
rect 6650 6170 6680 6180
rect 6740 6170 6900 6180
rect 7650 6170 7660 6180
rect 9220 6170 9240 6180
rect 9290 6170 9300 6180
rect 9610 6170 9620 6180
rect 9820 6170 9830 6180
rect 1260 6160 1270 6170
rect 1300 6160 1330 6170
rect 1420 6160 1430 6170
rect 1600 6160 1610 6170
rect 1630 6160 1650 6170
rect 1720 6160 1750 6170
rect 1770 6160 1780 6170
rect 2420 6160 2430 6170
rect 5300 6160 5310 6170
rect 5430 6160 5460 6170
rect 6660 6160 6690 6170
rect 6740 6160 6900 6170
rect 7650 6160 7660 6170
rect 9260 6160 9270 6170
rect 9650 6160 9670 6170
rect 9820 6160 9830 6170
rect 1290 6150 1300 6160
rect 1310 6150 1340 6160
rect 1350 6150 1360 6160
rect 1380 6150 1390 6160
rect 1610 6150 1630 6160
rect 1640 6150 1680 6160
rect 1720 6150 1740 6160
rect 2420 6150 2430 6160
rect 5280 6150 5290 6160
rect 5420 6150 5440 6160
rect 6660 6150 6690 6160
rect 6750 6150 6780 6160
rect 6800 6150 6900 6160
rect 7650 6150 7670 6160
rect 9230 6150 9240 6160
rect 9630 6150 9640 6160
rect 9820 6150 9830 6160
rect 1270 6140 1280 6150
rect 1300 6140 1310 6150
rect 1320 6140 1330 6150
rect 1400 6140 1420 6150
rect 1630 6140 1650 6150
rect 1680 6140 1740 6150
rect 2420 6140 2430 6150
rect 5270 6140 5280 6150
rect 5290 6140 5300 6150
rect 5420 6140 5430 6150
rect 6670 6140 6710 6150
rect 6750 6140 6780 6150
rect 6810 6140 6900 6150
rect 7650 6140 7670 6150
rect 9210 6140 9220 6150
rect 9830 6140 9840 6150
rect 1120 6130 1140 6140
rect 1390 6130 1400 6140
rect 1410 6130 1420 6140
rect 1430 6130 1440 6140
rect 1640 6130 1650 6140
rect 1770 6130 1790 6140
rect 4290 6130 4300 6140
rect 5270 6130 5290 6140
rect 5410 6130 5430 6140
rect 6680 6130 6720 6140
rect 6760 6130 6780 6140
rect 6810 6130 6830 6140
rect 6840 6130 6900 6140
rect 8520 6130 8550 6140
rect 9190 6130 9200 6140
rect 9950 6130 9960 6140
rect 1120 6120 1130 6130
rect 1270 6120 1290 6130
rect 1320 6120 1350 6130
rect 1360 6120 1370 6130
rect 1390 6120 1420 6130
rect 1430 6120 1440 6130
rect 1640 6120 1650 6130
rect 1770 6120 1790 6130
rect 2430 6120 2440 6130
rect 5260 6120 5270 6130
rect 5400 6120 5420 6130
rect 6690 6120 6730 6130
rect 6760 6120 6780 6130
rect 6840 6120 6900 6130
rect 6910 6120 6920 6130
rect 8520 6120 8540 6130
rect 9160 6120 9180 6130
rect 9840 6120 9850 6130
rect 9910 6120 9920 6130
rect 1280 6110 1290 6120
rect 1330 6110 1370 6120
rect 1400 6110 1430 6120
rect 1650 6110 1660 6120
rect 1760 6110 1790 6120
rect 2430 6110 2440 6120
rect 4300 6110 4310 6120
rect 5270 6110 5280 6120
rect 5390 6110 5410 6120
rect 6690 6110 6730 6120
rect 6830 6110 6920 6120
rect 7690 6110 7700 6120
rect 9130 6110 9180 6120
rect 9900 6110 9920 6120
rect 1290 6100 1300 6110
rect 1340 6100 1370 6110
rect 1400 6100 1430 6110
rect 1650 6100 1670 6110
rect 1750 6100 1790 6110
rect 3910 6100 3920 6110
rect 5250 6100 5260 6110
rect 5390 6100 5400 6110
rect 6700 6100 6730 6110
rect 6830 6100 6930 6110
rect 9100 6100 9160 6110
rect 9410 6100 9420 6110
rect 9450 6100 9460 6110
rect 9900 6100 9920 6110
rect 1360 6090 1370 6100
rect 1410 6090 1430 6100
rect 1640 6090 1680 6100
rect 1750 6090 1770 6100
rect 1780 6090 1790 6100
rect 3890 6090 3900 6100
rect 4310 6090 4320 6100
rect 5250 6090 5270 6100
rect 5380 6090 5390 6100
rect 6710 6090 6750 6100
rect 6840 6090 6950 6100
rect 9080 6090 9120 6100
rect 9470 6090 9480 6100
rect 9850 6090 9860 6100
rect 9940 6090 9950 6100
rect 1300 6080 1310 6090
rect 1420 6080 1430 6090
rect 1630 6080 1680 6090
rect 1750 6080 1770 6090
rect 1790 6080 1800 6090
rect 2440 6080 2450 6090
rect 2470 6080 2480 6090
rect 3880 6080 3890 6090
rect 5240 6080 5250 6090
rect 5380 6080 5390 6090
rect 6710 6080 6760 6090
rect 6840 6080 6950 6090
rect 9060 6080 9120 6090
rect 9480 6080 9490 6090
rect 9890 6080 9910 6090
rect 9930 6080 9960 6090
rect 1120 6070 1140 6080
rect 1300 6070 1310 6080
rect 1420 6070 1430 6080
rect 1610 6070 1690 6080
rect 1760 6070 1780 6080
rect 1790 6070 1800 6080
rect 4320 6070 4330 6080
rect 5210 6070 5220 6080
rect 5250 6070 5260 6080
rect 5370 6070 5380 6080
rect 6720 6070 6760 6080
rect 6770 6070 6780 6080
rect 6850 6070 6970 6080
rect 9010 6070 9020 6080
rect 9030 6070 9090 6080
rect 9900 6070 9950 6080
rect 1100 6060 1110 6070
rect 1300 6060 1310 6070
rect 1420 6060 1430 6070
rect 1610 6060 1700 6070
rect 1780 6060 1800 6070
rect 3780 6060 3790 6070
rect 5200 6060 5210 6070
rect 5240 6060 5250 6070
rect 5370 6060 5380 6070
rect 6720 6060 6790 6070
rect 6850 6060 6960 6070
rect 8980 6060 9010 6070
rect 9020 6060 9080 6070
rect 9400 6060 9430 6070
rect 1290 6050 1320 6060
rect 1610 6050 1730 6060
rect 3790 6050 3840 6060
rect 3980 6050 3990 6060
rect 5190 6050 5200 6060
rect 5370 6050 5380 6060
rect 6730 6050 6770 6060
rect 6830 6050 6960 6060
rect 8940 6050 9080 6060
rect 9240 6050 9250 6060
rect 9440 6050 9450 6060
rect 9860 6050 9870 6060
rect 830 6040 840 6050
rect 1200 6040 1230 6050
rect 1250 6040 1260 6050
rect 1270 6040 1320 6050
rect 1610 6040 1730 6050
rect 2460 6040 2470 6050
rect 3780 6040 3790 6050
rect 3810 6040 3820 6050
rect 3990 6040 4000 6050
rect 5230 6040 5240 6050
rect 5370 6040 5380 6050
rect 6730 6040 6780 6050
rect 6810 6040 6960 6050
rect 8930 6040 9050 6050
rect 9060 6040 9070 6050
rect 9210 6040 9220 6050
rect 9340 6040 9350 6050
rect 9860 6040 9870 6050
rect 830 6030 840 6040
rect 860 6030 880 6040
rect 1160 6030 1210 6040
rect 1250 6030 1320 6040
rect 1620 6030 1730 6040
rect 5220 6030 5240 6040
rect 5370 6030 5380 6040
rect 6740 6030 6770 6040
rect 6810 6030 6840 6040
rect 6850 6030 6970 6040
rect 8860 6030 9020 6040
rect 9340 6030 9350 6040
rect 9390 6030 9400 6040
rect 9430 6030 9440 6040
rect 9480 6030 9490 6040
rect 9860 6030 9870 6040
rect 840 6020 890 6030
rect 900 6020 940 6030
rect 1130 6020 1170 6030
rect 1190 6020 1210 6030
rect 1230 6020 1240 6030
rect 1260 6020 1300 6030
rect 1310 6020 1320 6030
rect 1620 6020 1680 6030
rect 1700 6020 1720 6030
rect 3230 6020 3240 6030
rect 4340 6020 4350 6030
rect 5200 6020 5220 6030
rect 6740 6020 6770 6030
rect 6820 6020 6980 6030
rect 8830 6020 8850 6030
rect 8900 6020 8910 6030
rect 9270 6020 9280 6030
rect 9390 6020 9400 6030
rect 9410 6020 9420 6030
rect 9860 6020 9870 6030
rect 830 6010 850 6020
rect 890 6010 940 6020
rect 1130 6010 1150 6020
rect 1170 6010 1190 6020
rect 1250 6010 1280 6020
rect 1310 6010 1320 6020
rect 1640 6010 1660 6020
rect 1670 6010 1680 6020
rect 1710 6010 1720 6020
rect 2480 6010 2490 6020
rect 4030 6010 4040 6020
rect 5190 6010 5220 6020
rect 5360 6010 5370 6020
rect 6740 6010 6790 6020
rect 6810 6010 6980 6020
rect 8420 6010 8430 6020
rect 8800 6010 8830 6020
rect 9100 6010 9110 6020
rect 9130 6010 9140 6020
rect 9240 6010 9250 6020
rect 760 6000 770 6010
rect 830 6000 850 6010
rect 910 6000 950 6010
rect 1120 6000 1160 6010
rect 1170 6000 1190 6010
rect 1250 6000 1280 6010
rect 1640 6000 1660 6010
rect 1670 6000 1680 6010
rect 1700 6000 1720 6010
rect 3200 6000 3230 6010
rect 4040 6000 4050 6010
rect 5180 6000 5210 6010
rect 5350 6000 5370 6010
rect 6750 6000 6800 6010
rect 6810 6000 6820 6010
rect 6850 6000 6920 6010
rect 6930 6000 6980 6010
rect 8770 6000 8820 6010
rect 9090 6000 9100 6010
rect 9140 6000 9150 6010
rect 9170 6000 9180 6010
rect 9350 6000 9360 6010
rect 9930 6000 9950 6010
rect 760 5990 770 6000
rect 830 5990 850 6000
rect 920 5990 950 6000
rect 1120 5990 1170 6000
rect 1200 5990 1210 6000
rect 1250 5990 1270 6000
rect 1650 5990 1660 6000
rect 1700 5990 1720 6000
rect 3180 5990 3240 6000
rect 3810 5990 3830 6000
rect 5180 5990 5200 6000
rect 5360 5990 5370 6000
rect 6750 5990 6800 6000
rect 6860 5990 6910 6000
rect 6940 5990 6980 6000
rect 8410 5990 8420 6000
rect 8760 5990 8800 6000
rect 9040 5990 9050 6000
rect 9060 5990 9070 6000
rect 9080 5990 9100 6000
rect 9170 5990 9180 6000
rect 9350 5990 9360 6000
rect 9940 5990 9960 6000
rect 750 5980 770 5990
rect 840 5980 850 5990
rect 880 5980 910 5990
rect 920 5980 970 5990
rect 1130 5980 1140 5990
rect 1170 5980 1180 5990
rect 1190 5980 1200 5990
rect 1650 5980 1660 5990
rect 1690 5980 1710 5990
rect 3180 5980 3250 5990
rect 4070 5980 4080 5990
rect 5170 5980 5190 5990
rect 5360 5980 5370 5990
rect 6760 5980 6810 5990
rect 6950 5980 6990 5990
rect 8720 5980 8730 5990
rect 8740 5980 8770 5990
rect 9020 5980 9030 5990
rect 9070 5980 9100 5990
rect 9160 5980 9190 5990
rect 9230 5980 9240 5990
rect 9280 5980 9300 5990
rect 9350 5980 9360 5990
rect 9890 5980 9900 5990
rect 9910 5980 9920 5990
rect 9940 5980 9950 5990
rect 750 5970 770 5980
rect 840 5970 850 5980
rect 900 5970 910 5980
rect 930 5970 980 5980
rect 1120 5970 1130 5980
rect 1180 5970 1190 5980
rect 1690 5970 1720 5980
rect 2510 5970 2520 5980
rect 3170 5970 3250 5980
rect 5160 5970 5190 5980
rect 5350 5970 5360 5980
rect 6760 5970 6820 5980
rect 6950 5970 6990 5980
rect 8400 5970 8410 5980
rect 8670 5970 8760 5980
rect 8970 5970 9000 5980
rect 9010 5970 9030 5980
rect 9080 5970 9100 5980
rect 9150 5970 9190 5980
rect 9240 5970 9260 5980
rect 9410 5970 9420 5980
rect 740 5960 770 5970
rect 840 5960 850 5970
rect 860 5960 870 5970
rect 910 5960 920 5970
rect 950 5960 1050 5970
rect 1080 5960 1100 5970
rect 1110 5960 1120 5970
rect 1160 5960 1180 5970
rect 1680 5960 1720 5970
rect 1780 5960 1790 5970
rect 1800 5960 1810 5970
rect 2520 5960 2530 5970
rect 3170 5960 3250 5970
rect 3770 5960 3780 5970
rect 3860 5960 3870 5970
rect 6770 5960 6820 5970
rect 6960 5960 6990 5970
rect 8640 5960 8650 5970
rect 8670 5960 8680 5970
rect 8960 5960 8970 5970
rect 9000 5960 9030 5970
rect 9090 5960 9100 5970
rect 9160 5960 9190 5970
rect 9360 5960 9370 5970
rect 9410 5960 9420 5970
rect 9490 5960 9500 5970
rect 9890 5960 9900 5970
rect 9930 5960 9950 5970
rect 9960 5960 9980 5970
rect 740 5950 760 5960
rect 840 5950 850 5960
rect 920 5950 980 5960
rect 1000 5950 1070 5960
rect 1090 5950 1100 5960
rect 1160 5950 1170 5960
rect 1680 5950 1710 5960
rect 1720 5950 1730 5960
rect 2530 5950 2540 5960
rect 3160 5950 3190 5960
rect 3200 5950 3250 5960
rect 3870 5950 3880 5960
rect 4120 5950 4130 5960
rect 4340 5950 4350 5960
rect 5340 5950 5350 5960
rect 6780 5950 6820 5960
rect 6950 5950 6960 5960
rect 6970 5950 7000 5960
rect 8610 5950 8620 5960
rect 8630 5950 8640 5960
rect 9010 5950 9030 5960
rect 9150 5950 9200 5960
rect 9300 5950 9310 5960
rect 9360 5950 9370 5960
rect 9440 5950 9450 5960
rect 9900 5950 9920 5960
rect 9940 5950 9950 5960
rect 730 5940 760 5950
rect 800 5940 840 5950
rect 920 5940 960 5950
rect 1040 5940 1060 5950
rect 1680 5940 1700 5950
rect 2540 5940 2550 5950
rect 3150 5940 3180 5950
rect 3210 5940 3250 5950
rect 3870 5940 3880 5950
rect 4140 5940 4150 5950
rect 5340 5940 5350 5950
rect 6790 5940 6830 5950
rect 6940 5940 7000 5950
rect 8380 5940 8390 5950
rect 8580 5940 8590 5950
rect 8950 5940 8960 5950
rect 9020 5940 9030 5950
rect 9150 5940 9170 5950
rect 9180 5940 9200 5950
rect 9450 5940 9460 5950
rect 720 5930 730 5940
rect 750 5930 760 5940
rect 780 5930 790 5940
rect 800 5930 840 5940
rect 930 5930 970 5940
rect 1690 5930 1700 5940
rect 2520 5930 2540 5940
rect 2550 5930 2560 5940
rect 3140 5930 3170 5940
rect 3210 5930 3250 5940
rect 3880 5930 3890 5940
rect 5340 5930 5350 5940
rect 6790 5930 6820 5940
rect 6950 5930 7000 5940
rect 8130 5930 8150 5940
rect 8540 5930 8570 5940
rect 8900 5930 8920 5940
rect 8950 5930 8970 5940
rect 9020 5930 9030 5940
rect 9150 5930 9200 5940
rect 9250 5930 9260 5940
rect 9460 5930 9470 5940
rect 710 5920 730 5930
rect 740 5920 750 5930
rect 760 5920 790 5930
rect 810 5920 840 5930
rect 940 5920 950 5930
rect 1700 5920 1720 5930
rect 2540 5920 2550 5930
rect 3120 5920 3160 5930
rect 3210 5920 3260 5930
rect 3890 5920 3900 5930
rect 4170 5920 4180 5930
rect 4330 5920 4340 5930
rect 6800 5920 6830 5930
rect 6950 5920 7000 5930
rect 8100 5920 8150 5930
rect 8520 5920 8540 5930
rect 8940 5920 8970 5930
rect 9160 5920 9200 5930
rect 9370 5920 9380 5930
rect 9420 5920 9430 5930
rect 9480 5920 9500 5930
rect 700 5910 720 5920
rect 740 5910 750 5920
rect 760 5910 770 5920
rect 940 5910 950 5920
rect 1710 5910 1740 5920
rect 2560 5910 2590 5920
rect 3120 5910 3150 5920
rect 3220 5910 3260 5920
rect 3910 5910 3920 5920
rect 5130 5910 5140 5920
rect 5330 5910 5340 5920
rect 6800 5910 6830 5920
rect 6960 5910 7000 5920
rect 8090 5910 8100 5920
rect 8120 5910 8150 5920
rect 8480 5910 8530 5920
rect 8810 5910 8820 5920
rect 8940 5910 8980 5920
rect 9170 5910 9200 5920
rect 9250 5910 9260 5920
rect 9370 5910 9380 5920
rect 9420 5910 9430 5920
rect 700 5900 720 5910
rect 750 5900 770 5910
rect 810 5900 820 5910
rect 950 5900 960 5910
rect 1720 5900 1740 5910
rect 2560 5900 2600 5910
rect 3100 5900 3150 5910
rect 3220 5900 3260 5910
rect 3750 5900 3760 5910
rect 4300 5900 4310 5910
rect 5330 5900 5340 5910
rect 6800 5900 6820 5910
rect 6960 5900 7000 5910
rect 8090 5900 8100 5910
rect 8120 5900 8150 5910
rect 8360 5900 8370 5910
rect 8450 5900 8460 5910
rect 8500 5900 8510 5910
rect 8800 5900 8810 5910
rect 8940 5900 8980 5910
rect 9180 5900 9210 5910
rect 9250 5900 9260 5910
rect 9300 5900 9320 5910
rect 9330 5900 9340 5910
rect 9900 5900 9910 5910
rect 690 5890 710 5900
rect 730 5890 740 5900
rect 790 5890 820 5900
rect 950 5890 970 5900
rect 1730 5890 1740 5900
rect 2570 5890 2610 5900
rect 3100 5890 3140 5900
rect 3220 5890 3250 5900
rect 3750 5890 3770 5900
rect 4260 5890 4280 5900
rect 5120 5890 5130 5900
rect 5330 5890 5340 5900
rect 6800 5890 6830 5900
rect 6960 5890 7000 5900
rect 8090 5890 8100 5900
rect 8130 5890 8150 5900
rect 8420 5890 8440 5900
rect 8700 5890 8720 5900
rect 8750 5890 8760 5900
rect 8850 5890 8860 5900
rect 8870 5890 8900 5900
rect 8950 5890 8980 5900
rect 9070 5890 9080 5900
rect 9170 5890 9190 5900
rect 9200 5890 9210 5900
rect 9260 5890 9280 5900
rect 9390 5890 9410 5900
rect 9900 5890 9910 5900
rect 710 5880 800 5890
rect 940 5880 980 5890
rect 1740 5880 1770 5890
rect 1780 5880 1790 5890
rect 1830 5880 1850 5890
rect 2590 5880 2610 5890
rect 3080 5880 3110 5890
rect 3230 5880 3250 5890
rect 3920 5880 3940 5890
rect 5120 5880 5150 5890
rect 5330 5880 5340 5890
rect 6800 5880 6830 5890
rect 6960 5880 7010 5890
rect 8090 5880 8100 5890
rect 8390 5880 8400 5890
rect 8680 5880 8690 5890
rect 8790 5880 8800 5890
rect 8840 5880 8850 5890
rect 8870 5880 8900 5890
rect 8960 5880 8990 5890
rect 9070 5880 9080 5890
rect 9160 5880 9210 5890
rect 690 5870 710 5880
rect 720 5870 770 5880
rect 780 5870 790 5880
rect 980 5870 990 5880
rect 1780 5870 1810 5880
rect 1840 5870 1850 5880
rect 2600 5870 2620 5880
rect 3060 5870 3100 5880
rect 3230 5870 3250 5880
rect 3740 5870 3760 5880
rect 5120 5870 5140 5880
rect 6800 5870 6830 5880
rect 6960 5870 6990 5880
rect 7000 5870 7010 5880
rect 8350 5870 8360 5880
rect 8650 5870 8660 5880
rect 8790 5870 8800 5880
rect 8880 5870 8900 5880
rect 8950 5870 8990 5880
rect 9070 5870 9090 5880
rect 9160 5870 9210 5880
rect 9330 5870 9340 5880
rect 670 5860 710 5870
rect 720 5860 770 5870
rect 870 5860 890 5870
rect 1840 5860 1850 5870
rect 2590 5860 2630 5870
rect 3040 5860 3080 5870
rect 3240 5860 3260 5870
rect 3930 5860 3940 5870
rect 5120 5860 5130 5870
rect 5320 5860 5330 5870
rect 6780 5860 6830 5870
rect 6970 5860 6990 5870
rect 7910 5860 7920 5870
rect 7940 5860 7960 5870
rect 8140 5860 8150 5870
rect 8320 5860 8330 5870
rect 8620 5860 8630 5870
rect 8790 5860 8800 5870
rect 8890 5860 8910 5870
rect 8950 5860 8960 5870
rect 8970 5860 8990 5870
rect 9070 5860 9100 5870
rect 9190 5860 9210 5870
rect 9310 5860 9320 5870
rect 650 5850 670 5860
rect 690 5850 700 5860
rect 720 5850 770 5860
rect 790 5850 800 5860
rect 820 5850 830 5860
rect 870 5850 880 5860
rect 2600 5850 2650 5860
rect 3000 5850 3060 5860
rect 3230 5850 3270 5860
rect 3740 5850 3750 5860
rect 5320 5850 5330 5860
rect 6780 5850 6830 5860
rect 7890 5850 7910 5860
rect 7950 5850 7960 5860
rect 8090 5850 8100 5860
rect 8140 5850 8150 5860
rect 8280 5850 8300 5860
rect 8790 5850 8800 5860
rect 8900 5850 8910 5860
rect 8980 5850 9000 5860
rect 9080 5850 9100 5860
rect 9200 5850 9220 5860
rect 9270 5850 9280 5860
rect 630 5840 660 5850
rect 720 5840 730 5850
rect 740 5840 770 5850
rect 780 5840 790 5850
rect 810 5840 830 5850
rect 880 5840 890 5850
rect 1850 5840 1860 5850
rect 2310 5840 2360 5850
rect 2610 5840 2660 5850
rect 2980 5840 3050 5850
rect 3230 5840 3260 5850
rect 3730 5840 3750 5850
rect 3790 5840 3800 5850
rect 3940 5840 3960 5850
rect 5320 5840 5330 5850
rect 6790 5840 6830 5850
rect 6990 5840 7000 5850
rect 7880 5840 7890 5850
rect 7950 5840 7960 5850
rect 8130 5840 8140 5850
rect 8250 5840 8260 5850
rect 8790 5840 8800 5850
rect 8840 5840 8850 5850
rect 8900 5840 8910 5850
rect 8980 5840 9000 5850
rect 9090 5840 9110 5850
rect 9210 5840 9220 5850
rect 9240 5840 9250 5850
rect 9910 5840 9920 5850
rect 600 5830 660 5840
rect 740 5830 760 5840
rect 2300 5830 2360 5840
rect 2620 5830 2670 5840
rect 2980 5830 3030 5840
rect 3230 5830 3260 5840
rect 3730 5830 3740 5840
rect 3800 5830 3830 5840
rect 5320 5830 5330 5840
rect 6800 5830 6830 5840
rect 6980 5830 6990 5840
rect 7890 5830 7900 5840
rect 7960 5830 7970 5840
rect 8230 5830 8240 5840
rect 8620 5830 8630 5840
rect 8640 5830 8670 5840
rect 8840 5830 8850 5840
rect 8900 5830 8920 5840
rect 8990 5830 9000 5840
rect 9100 5830 9120 5840
rect 590 5820 660 5830
rect 740 5820 750 5830
rect 2300 5820 2360 5830
rect 2620 5820 2670 5830
rect 2880 5820 2930 5830
rect 2950 5820 3020 5830
rect 3230 5820 3260 5830
rect 3730 5820 3740 5830
rect 3760 5820 3770 5830
rect 3800 5820 3880 5830
rect 5100 5820 5110 5830
rect 5320 5820 5330 5830
rect 6800 5820 6830 5830
rect 6980 5820 6990 5830
rect 7890 5820 7900 5830
rect 7970 5820 7980 5830
rect 8200 5820 8210 5830
rect 8660 5820 8680 5830
rect 8800 5820 8810 5830
rect 8910 5820 8920 5830
rect 8960 5820 8970 5830
rect 8990 5820 9010 5830
rect 9110 5820 9120 5830
rect 9940 5820 9960 5830
rect 580 5810 630 5820
rect 650 5810 660 5820
rect 730 5810 740 5820
rect 2290 5810 2350 5820
rect 2620 5810 2690 5820
rect 2870 5810 3000 5820
rect 3230 5810 3260 5820
rect 3720 5810 3750 5820
rect 3760 5810 3780 5820
rect 3830 5810 3850 5820
rect 3950 5810 3970 5820
rect 5100 5810 5110 5820
rect 5320 5810 5330 5820
rect 6800 5810 6830 5820
rect 6970 5810 7000 5820
rect 7890 5810 7900 5820
rect 7970 5810 8010 5820
rect 8170 5810 8180 5820
rect 8670 5810 8680 5820
rect 8720 5810 8730 5820
rect 8790 5810 8810 5820
rect 8910 5810 8920 5820
rect 8960 5810 8970 5820
rect 8990 5810 9010 5820
rect 9940 5810 9950 5820
rect 570 5800 580 5810
rect 590 5800 610 5810
rect 650 5800 660 5810
rect 730 5800 740 5810
rect 880 5800 890 5810
rect 2270 5800 2350 5810
rect 2610 5800 2700 5810
rect 2850 5800 3000 5810
rect 3230 5800 3260 5810
rect 3770 5800 3780 5810
rect 3790 5800 3800 5810
rect 3820 5800 3840 5810
rect 5320 5800 5330 5810
rect 6800 5800 6830 5810
rect 6970 5800 7000 5810
rect 7890 5800 7930 5810
rect 7940 5800 7950 5810
rect 7990 5800 8010 5810
rect 8140 5800 8150 5810
rect 8670 5800 8680 5810
rect 8800 5800 8810 5810
rect 8850 5800 8860 5810
rect 8900 5800 8920 5810
rect 8960 5800 8970 5810
rect 9000 5800 9020 5810
rect 9060 5800 9070 5810
rect 9940 5800 9950 5810
rect 560 5790 580 5800
rect 600 5790 610 5800
rect 650 5790 660 5800
rect 700 5790 720 5800
rect 880 5790 900 5800
rect 1850 5790 1870 5800
rect 2260 5790 2350 5800
rect 2610 5790 2690 5800
rect 2830 5790 2970 5800
rect 3240 5790 3260 5800
rect 3800 5790 3810 5800
rect 3880 5790 3890 5800
rect 3920 5790 3930 5800
rect 4060 5790 4070 5800
rect 5310 5790 5330 5800
rect 6810 5790 6830 5800
rect 6980 5790 7000 5800
rect 7900 5790 7910 5800
rect 7940 5790 7990 5800
rect 8110 5790 8120 5800
rect 8390 5790 8410 5800
rect 8670 5790 8690 5800
rect 8900 5790 8910 5800
rect 8960 5790 8970 5800
rect 9010 5790 9030 5800
rect 550 5780 570 5790
rect 590 5780 610 5790
rect 650 5780 700 5790
rect 810 5780 820 5790
rect 1850 5780 1870 5790
rect 2250 5780 2300 5790
rect 2320 5780 2340 5790
rect 2600 5780 2670 5790
rect 2830 5780 2960 5790
rect 3240 5780 3260 5790
rect 3920 5780 3930 5790
rect 3960 5780 3970 5790
rect 4070 5780 4080 5790
rect 5090 5780 5100 5790
rect 5310 5780 5330 5790
rect 6810 5780 6830 5790
rect 6980 5780 6990 5790
rect 7740 5780 7780 5790
rect 8070 5780 8080 5790
rect 8380 5780 8390 5790
rect 8680 5780 8690 5790
rect 8810 5780 8820 5790
rect 8860 5780 8870 5790
rect 8890 5780 8900 5790
rect 570 5770 600 5780
rect 650 5770 690 5780
rect 780 5770 790 5780
rect 810 5770 820 5780
rect 870 5770 900 5780
rect 1870 5770 1880 5780
rect 2230 5770 2280 5780
rect 2310 5770 2330 5780
rect 2600 5770 2670 5780
rect 2810 5770 2960 5780
rect 3240 5770 3260 5780
rect 3800 5770 3830 5780
rect 3850 5770 3870 5780
rect 5090 5770 5100 5780
rect 5310 5770 5320 5780
rect 6810 5770 6840 5780
rect 6980 5770 6990 5780
rect 8030 5770 8050 5780
rect 8680 5770 8690 5780
rect 8810 5770 8820 5780
rect 9940 5770 9950 5780
rect 660 5760 680 5770
rect 780 5760 790 5770
rect 860 5760 880 5770
rect 1870 5760 1880 5770
rect 2240 5760 2270 5770
rect 2310 5760 2320 5770
rect 2590 5760 2650 5770
rect 2800 5760 2960 5770
rect 3240 5760 3260 5770
rect 3790 5760 3850 5770
rect 3890 5760 3900 5770
rect 3920 5760 3930 5770
rect 5090 5760 5100 5770
rect 5300 5760 5320 5770
rect 6820 5760 6840 5770
rect 6980 5760 6990 5770
rect 7990 5760 8020 5770
rect 8420 5760 8430 5770
rect 8730 5760 8740 5770
rect 8820 5760 8830 5770
rect 9940 5760 9950 5770
rect 790 5750 800 5760
rect 870 5750 880 5760
rect 1870 5750 1880 5760
rect 2220 5750 2260 5760
rect 2300 5750 2320 5760
rect 2560 5750 2570 5760
rect 2580 5750 2640 5760
rect 2790 5750 2970 5760
rect 3230 5750 3260 5760
rect 3740 5750 3760 5760
rect 3820 5750 3830 5760
rect 3840 5750 3860 5760
rect 5300 5750 5310 5760
rect 6810 5750 6840 5760
rect 6970 5750 6990 5760
rect 7970 5750 7990 5760
rect 8380 5750 8390 5760
rect 8690 5750 8700 5760
rect 8830 5750 8840 5760
rect 9940 5750 9950 5760
rect 630 5740 700 5750
rect 770 5740 780 5750
rect 800 5740 820 5750
rect 870 5740 880 5750
rect 1870 5740 1890 5750
rect 2220 5740 2250 5750
rect 2290 5740 2310 5750
rect 2550 5740 2620 5750
rect 2780 5740 2960 5750
rect 3230 5740 3260 5750
rect 3730 5740 3760 5750
rect 3770 5740 3790 5750
rect 5080 5740 5090 5750
rect 5290 5740 5310 5750
rect 6820 5740 6840 5750
rect 6970 5740 6980 5750
rect 7930 5740 7960 5750
rect 8380 5740 8390 5750
rect 8690 5740 8700 5750
rect 8840 5740 8860 5750
rect 9950 5740 9960 5750
rect 610 5730 660 5740
rect 680 5730 720 5740
rect 820 5730 850 5740
rect 1860 5730 1900 5740
rect 2220 5730 2250 5740
rect 2290 5730 2300 5740
rect 2530 5730 2610 5740
rect 2760 5730 2960 5740
rect 3230 5730 3260 5740
rect 3700 5730 3710 5740
rect 3740 5730 3750 5740
rect 3800 5730 3810 5740
rect 3940 5730 3950 5740
rect 3960 5730 3970 5740
rect 5290 5730 5300 5740
rect 6820 5730 6840 5740
rect 6970 5730 6980 5740
rect 7910 5730 7920 5740
rect 8380 5730 8390 5740
rect 8690 5730 8700 5740
rect 8740 5730 8750 5740
rect 9950 5730 9960 5740
rect 760 5720 770 5730
rect 1860 5720 1910 5730
rect 2210 5720 2240 5730
rect 2280 5720 2290 5730
rect 2530 5720 2580 5730
rect 2770 5720 2830 5730
rect 2840 5720 2950 5730
rect 3230 5720 3260 5730
rect 3760 5720 3770 5730
rect 3820 5720 3830 5730
rect 4010 5720 4020 5730
rect 4390 5720 4400 5730
rect 5290 5720 5300 5730
rect 6820 5720 6840 5730
rect 6910 5720 6930 5730
rect 6970 5720 6980 5730
rect 7800 5720 7820 5730
rect 7890 5720 7910 5730
rect 8210 5720 8220 5730
rect 8230 5720 8240 5730
rect 8280 5720 8290 5730
rect 8430 5720 8440 5730
rect 9950 5720 9960 5730
rect 1210 5710 1230 5720
rect 1860 5710 1910 5720
rect 2210 5710 2240 5720
rect 2530 5710 2570 5720
rect 2760 5710 2820 5720
rect 2930 5710 2940 5720
rect 3230 5710 3260 5720
rect 3750 5710 3770 5720
rect 3780 5710 3790 5720
rect 3840 5710 3850 5720
rect 5280 5710 5300 5720
rect 6830 5710 6850 5720
rect 6900 5710 6920 5720
rect 6930 5710 6950 5720
rect 6960 5710 6980 5720
rect 7770 5710 7790 5720
rect 7840 5710 7860 5720
rect 7890 5710 7910 5720
rect 8170 5710 8180 5720
rect 8240 5710 8250 5720
rect 8390 5710 8400 5720
rect 9950 5710 9960 5720
rect 1170 5700 1180 5710
rect 1210 5700 1220 5710
rect 1860 5700 1930 5710
rect 2210 5700 2230 5710
rect 2510 5700 2560 5710
rect 2720 5700 2750 5710
rect 2760 5700 2810 5710
rect 3230 5700 3260 5710
rect 3750 5700 3770 5710
rect 3840 5700 3870 5710
rect 5070 5700 5080 5710
rect 5110 5700 5120 5710
rect 5290 5700 5300 5710
rect 6840 5700 6850 5710
rect 6930 5700 6960 5710
rect 7740 5700 7750 5710
rect 7800 5700 7920 5710
rect 8150 5700 8180 5710
rect 8220 5700 8250 5710
rect 8390 5700 8400 5710
rect 8700 5700 8710 5710
rect 8740 5700 8750 5710
rect 9960 5700 9970 5710
rect 810 5690 820 5700
rect 1180 5690 1200 5700
rect 1870 5690 1940 5700
rect 2200 5690 2220 5700
rect 2480 5690 2550 5700
rect 2710 5690 2750 5700
rect 2760 5690 2800 5700
rect 3240 5690 3260 5700
rect 3750 5690 3760 5700
rect 3800 5690 3810 5700
rect 3860 5690 3900 5700
rect 4260 5690 4270 5700
rect 5070 5690 5080 5700
rect 5100 5690 5120 5700
rect 5280 5690 5290 5700
rect 6840 5690 6860 5700
rect 6940 5690 6980 5700
rect 7750 5690 7800 5700
rect 7810 5690 7920 5700
rect 8150 5690 8180 5700
rect 8220 5690 8250 5700
rect 8390 5690 8400 5700
rect 8720 5690 8740 5700
rect 810 5680 820 5690
rect 1070 5680 1080 5690
rect 1140 5680 1180 5690
rect 1860 5680 1930 5690
rect 2210 5680 2220 5690
rect 2260 5680 2270 5690
rect 2470 5680 2540 5690
rect 2690 5680 2750 5690
rect 2770 5680 2800 5690
rect 3210 5680 3220 5690
rect 3240 5680 3270 5690
rect 3790 5680 3800 5690
rect 3910 5680 3930 5690
rect 5070 5680 5080 5690
rect 5090 5680 5120 5690
rect 5280 5680 5300 5690
rect 6840 5680 6860 5690
rect 6910 5680 6980 5690
rect 7740 5680 7750 5690
rect 7810 5680 7880 5690
rect 7900 5680 7920 5690
rect 8030 5680 8040 5690
rect 8050 5680 8060 5690
rect 8100 5680 8110 5690
rect 8150 5680 8180 5690
rect 8230 5680 8250 5690
rect 8390 5680 8400 5690
rect 8440 5680 8450 5690
rect 800 5670 810 5680
rect 1870 5670 1930 5680
rect 2200 5670 2220 5680
rect 2260 5670 2270 5680
rect 2470 5670 2530 5680
rect 2680 5670 2800 5680
rect 3210 5670 3220 5680
rect 3250 5670 3270 5680
rect 3790 5670 3800 5680
rect 3820 5670 3830 5680
rect 3910 5670 3920 5680
rect 5070 5670 5100 5680
rect 5110 5670 5130 5680
rect 5280 5670 5290 5680
rect 6850 5670 6860 5680
rect 6910 5670 6950 5680
rect 6960 5670 6970 5680
rect 7710 5670 7730 5680
rect 7820 5670 7880 5680
rect 7900 5670 7920 5680
rect 8020 5670 8030 5680
rect 8060 5670 8070 5680
rect 8090 5670 8110 5680
rect 8160 5670 8190 5680
rect 8230 5670 8250 5680
rect 8290 5670 8300 5680
rect 800 5660 810 5670
rect 1870 5660 1940 5670
rect 2190 5660 2210 5670
rect 2250 5660 2260 5670
rect 2470 5660 2530 5670
rect 2650 5660 2800 5670
rect 3250 5660 3260 5670
rect 4220 5660 4240 5670
rect 4400 5660 4410 5670
rect 5070 5660 5100 5670
rect 5130 5660 5140 5670
rect 5280 5660 5290 5670
rect 6850 5660 6860 5670
rect 6930 5660 6940 5670
rect 7690 5660 7720 5670
rect 7820 5660 7890 5670
rect 7900 5660 7920 5670
rect 8010 5660 8020 5670
rect 8070 5660 8080 5670
rect 8090 5660 8120 5670
rect 8160 5660 8190 5670
rect 8230 5660 8260 5670
rect 8400 5660 8410 5670
rect 8500 5660 8520 5670
rect 780 5650 810 5660
rect 1880 5650 1960 5660
rect 2190 5650 2210 5660
rect 2250 5650 2260 5660
rect 2480 5650 2520 5660
rect 2660 5650 2800 5660
rect 3250 5650 3260 5660
rect 3690 5650 3700 5660
rect 3730 5650 3750 5660
rect 3790 5650 3800 5660
rect 3910 5650 3920 5660
rect 3980 5650 3990 5660
rect 4220 5650 4240 5660
rect 5070 5650 5100 5660
rect 5280 5650 5290 5660
rect 6850 5650 6870 5660
rect 6940 5650 6950 5660
rect 7650 5650 7710 5660
rect 7820 5650 7890 5660
rect 7900 5650 7920 5660
rect 8010 5650 8030 5660
rect 8090 5650 8120 5660
rect 8160 5650 8190 5660
rect 8230 5650 8260 5660
rect 8400 5650 8410 5660
rect 760 5640 800 5650
rect 1880 5640 1960 5650
rect 2180 5640 2210 5650
rect 2470 5640 2500 5650
rect 2640 5640 2730 5650
rect 2760 5640 2810 5650
rect 3250 5640 3260 5650
rect 3720 5640 3740 5650
rect 6850 5640 6870 5650
rect 6950 5640 6970 5650
rect 7620 5640 7690 5650
rect 7820 5640 7920 5650
rect 8010 5640 8030 5650
rect 8070 5640 8080 5650
rect 8090 5640 8120 5650
rect 8170 5640 8190 5650
rect 8230 5640 8260 5650
rect 8390 5640 8410 5650
rect 620 5630 630 5640
rect 750 5630 770 5640
rect 1890 5630 1940 5640
rect 1950 5630 1960 5640
rect 2180 5630 2200 5640
rect 2240 5630 2250 5640
rect 2470 5630 2500 5640
rect 2640 5630 2730 5640
rect 2790 5630 2810 5640
rect 3250 5630 3270 5640
rect 3730 5630 3740 5640
rect 3790 5630 3800 5640
rect 3810 5630 3820 5640
rect 3840 5630 3850 5640
rect 5720 5630 5760 5640
rect 6860 5630 6870 5640
rect 6960 5630 6970 5640
rect 7580 5630 7700 5640
rect 7830 5630 7920 5640
rect 8000 5630 8030 5640
rect 8070 5630 8120 5640
rect 8170 5630 8190 5640
rect 8240 5630 8260 5640
rect 8300 5630 8310 5640
rect 8400 5630 8410 5640
rect 8520 5630 8530 5640
rect 9980 5630 9990 5640
rect 620 5620 630 5630
rect 740 5620 750 5630
rect 1890 5620 1900 5630
rect 1930 5620 1940 5630
rect 1950 5620 1960 5630
rect 2180 5620 2190 5630
rect 2240 5620 2250 5630
rect 2470 5620 2480 5630
rect 2640 5620 2720 5630
rect 2800 5620 2820 5630
rect 3250 5620 3260 5630
rect 4190 5620 4220 5630
rect 5080 5620 5100 5630
rect 5270 5620 5280 5630
rect 5600 5620 5780 5630
rect 6860 5620 6880 5630
rect 7530 5620 7690 5630
rect 7820 5620 7840 5630
rect 7900 5620 7930 5630
rect 8010 5620 8030 5630
rect 8070 5620 8100 5630
rect 8170 5620 8200 5630
rect 8240 5620 8260 5630
rect 8300 5620 8310 5630
rect 8400 5620 8410 5630
rect 8500 5620 8510 5630
rect 9980 5620 9990 5630
rect 720 5610 730 5620
rect 1930 5610 1950 5620
rect 2180 5610 2190 5620
rect 2240 5610 2250 5620
rect 2460 5610 2470 5620
rect 2630 5610 2720 5620
rect 2810 5610 2840 5620
rect 3240 5610 3270 5620
rect 3790 5610 3800 5620
rect 5110 5610 5120 5620
rect 5270 5610 5280 5620
rect 5580 5610 5640 5620
rect 5740 5610 5820 5620
rect 6870 5610 6880 5620
rect 6950 5610 6960 5620
rect 7480 5610 7490 5620
rect 7500 5610 7680 5620
rect 7800 5610 7810 5620
rect 7910 5610 7930 5620
rect 8010 5610 8030 5620
rect 8170 5610 8200 5620
rect 8240 5610 8270 5620
rect 8340 5610 8350 5620
rect 8400 5610 8420 5620
rect 9970 5610 9990 5620
rect 710 5600 720 5610
rect 1940 5600 1950 5610
rect 2180 5600 2190 5610
rect 2450 5600 2470 5610
rect 2640 5600 2720 5610
rect 2820 5600 2870 5610
rect 3250 5600 3270 5610
rect 3670 5600 3680 5610
rect 3790 5600 3800 5610
rect 5270 5600 5280 5610
rect 5560 5600 5590 5610
rect 5770 5600 5840 5610
rect 6950 5600 6970 5610
rect 7450 5600 7500 5610
rect 7510 5600 7520 5610
rect 7530 5600 7570 5610
rect 7590 5600 7680 5610
rect 7790 5600 7800 5610
rect 7920 5600 7930 5610
rect 8010 5600 8030 5610
rect 8170 5600 8200 5610
rect 8240 5600 8270 5610
rect 8310 5600 8320 5610
rect 8390 5600 8400 5610
rect 9050 5600 9060 5610
rect 9980 5600 9990 5610
rect 1940 5590 1950 5600
rect 2180 5590 2190 5600
rect 2440 5590 2470 5600
rect 2610 5590 2660 5600
rect 2680 5590 2710 5600
rect 2840 5590 2860 5600
rect 3250 5590 3270 5600
rect 3430 5590 3440 5600
rect 3660 5590 3670 5600
rect 3870 5590 3880 5600
rect 4190 5590 4210 5600
rect 5100 5590 5110 5600
rect 5520 5590 5580 5600
rect 5840 5590 5870 5600
rect 6320 5590 6420 5600
rect 6880 5590 6890 5600
rect 6950 5590 6960 5600
rect 7430 5590 7460 5600
rect 7540 5590 7570 5600
rect 7600 5590 7680 5600
rect 7780 5590 7790 5600
rect 7920 5590 7940 5600
rect 8010 5590 8040 5600
rect 8180 5590 8200 5600
rect 8250 5590 8270 5600
rect 8980 5590 8990 5600
rect 9070 5590 9080 5600
rect 9980 5590 9990 5600
rect 600 5580 610 5590
rect 670 5580 680 5590
rect 1940 5580 1950 5590
rect 2180 5580 2190 5590
rect 2230 5580 2240 5590
rect 2430 5580 2450 5590
rect 2620 5580 2690 5590
rect 2850 5580 2870 5590
rect 2890 5580 2900 5590
rect 3250 5580 3270 5590
rect 3670 5580 3680 5590
rect 3700 5580 3710 5590
rect 3860 5580 3870 5590
rect 4160 5580 4190 5590
rect 4200 5580 4210 5590
rect 5100 5580 5110 5590
rect 5490 5580 5580 5590
rect 5850 5580 5880 5590
rect 6300 5580 6460 5590
rect 6880 5580 6890 5590
rect 6950 5580 6960 5590
rect 7310 5580 7320 5590
rect 7410 5580 7430 5590
rect 7610 5580 7690 5590
rect 7700 5580 7720 5590
rect 7780 5580 7790 5590
rect 7930 5580 7940 5590
rect 8010 5580 8040 5590
rect 8100 5580 8140 5590
rect 8180 5580 8210 5590
rect 8250 5580 8270 5590
rect 8370 5580 8380 5590
rect 9080 5580 9090 5590
rect 600 5570 610 5580
rect 660 5570 670 5580
rect 1940 5570 1950 5580
rect 2170 5570 2190 5580
rect 2230 5570 2240 5580
rect 2420 5570 2450 5580
rect 2620 5570 2690 5580
rect 2860 5570 2880 5580
rect 2910 5570 2920 5580
rect 3240 5570 3270 5580
rect 3450 5570 3460 5580
rect 3660 5570 3680 5580
rect 3690 5570 3700 5580
rect 3770 5570 3780 5580
rect 3850 5570 3860 5580
rect 4170 5570 4190 5580
rect 4210 5570 4220 5580
rect 5100 5570 5110 5580
rect 5260 5570 5270 5580
rect 5490 5570 5590 5580
rect 5870 5570 5900 5580
rect 6240 5570 6250 5580
rect 6270 5570 6330 5580
rect 6420 5570 6530 5580
rect 6540 5570 6550 5580
rect 6880 5570 6890 5580
rect 6950 5570 6970 5580
rect 7370 5570 7390 5580
rect 7540 5570 7550 5580
rect 7610 5570 7680 5580
rect 7760 5570 7770 5580
rect 7830 5570 7880 5580
rect 7930 5570 7950 5580
rect 8020 5570 8040 5580
rect 8100 5570 8110 5580
rect 8120 5570 8140 5580
rect 8180 5570 8210 5580
rect 8250 5570 8280 5580
rect 8340 5570 8350 5580
rect 580 5560 610 5570
rect 650 5560 660 5570
rect 1930 5560 1960 5570
rect 2170 5560 2190 5570
rect 2230 5560 2240 5570
rect 2400 5560 2430 5570
rect 2620 5560 2680 5570
rect 2690 5560 2700 5570
rect 2870 5560 2900 5570
rect 2920 5560 2930 5570
rect 3240 5560 3260 5570
rect 3660 5560 3670 5570
rect 3740 5560 3750 5570
rect 3770 5560 3780 5570
rect 4100 5560 4110 5570
rect 5090 5560 5110 5570
rect 5260 5560 5270 5570
rect 5510 5560 5590 5570
rect 5880 5560 5940 5570
rect 6220 5560 6290 5570
rect 6450 5560 6580 5570
rect 6880 5560 6890 5570
rect 6950 5560 6960 5570
rect 7610 5560 7660 5570
rect 7830 5560 7880 5570
rect 7930 5560 7940 5570
rect 8020 5560 8040 5570
rect 8090 5560 8140 5570
rect 8180 5560 8210 5570
rect 8280 5560 8320 5570
rect 8890 5560 8900 5570
rect 8950 5560 8960 5570
rect 9010 5560 9030 5570
rect 9040 5560 9050 5570
rect 580 5550 600 5560
rect 1940 5550 1970 5560
rect 2170 5550 2190 5560
rect 2230 5550 2240 5560
rect 2400 5550 2430 5560
rect 2600 5550 2700 5560
rect 2870 5550 2920 5560
rect 2940 5550 2950 5560
rect 3230 5550 3260 5560
rect 3680 5550 3690 5560
rect 3700 5550 3710 5560
rect 3720 5550 3730 5560
rect 3760 5550 3770 5560
rect 3780 5550 3790 5560
rect 4100 5550 4110 5560
rect 4150 5550 4160 5560
rect 4200 5550 4210 5560
rect 5100 5550 5110 5560
rect 5500 5550 5630 5560
rect 5900 5550 5940 5560
rect 6200 5550 6270 5560
rect 6500 5550 6590 5560
rect 6890 5550 6900 5560
rect 7370 5550 7380 5560
rect 7620 5550 7650 5560
rect 7740 5550 7750 5560
rect 7840 5550 7880 5560
rect 7930 5550 7950 5560
rect 8020 5550 8050 5560
rect 8090 5550 8140 5560
rect 8180 5550 8190 5560
rect 8200 5550 8210 5560
rect 8860 5550 8870 5560
rect 9060 5550 9080 5560
rect 570 5540 580 5550
rect 650 5540 660 5550
rect 1940 5540 1960 5550
rect 2160 5540 2190 5550
rect 2230 5540 2240 5550
rect 2410 5540 2430 5550
rect 2590 5540 2690 5550
rect 2870 5540 2930 5550
rect 2950 5540 2960 5550
rect 3230 5540 3260 5550
rect 3660 5540 3680 5550
rect 3750 5540 3760 5550
rect 3820 5540 3830 5550
rect 4100 5540 4110 5550
rect 4140 5540 4150 5550
rect 4190 5540 4210 5550
rect 5490 5540 5550 5550
rect 5600 5540 5650 5550
rect 5900 5540 5950 5550
rect 6180 5540 6260 5550
rect 6540 5540 6600 5550
rect 6890 5540 6900 5550
rect 6950 5540 6960 5550
rect 7310 5540 7330 5550
rect 7370 5540 7380 5550
rect 7620 5540 7650 5550
rect 7790 5540 7800 5550
rect 7840 5540 7880 5550
rect 7940 5540 7950 5550
rect 8020 5540 8050 5550
rect 8090 5540 8110 5550
rect 8120 5540 8140 5550
rect 8180 5540 8190 5550
rect 8210 5540 8240 5550
rect 8940 5540 8950 5550
rect 8990 5540 9000 5550
rect 520 5530 540 5540
rect 560 5530 570 5540
rect 620 5530 630 5540
rect 930 5530 950 5540
rect 1940 5530 1970 5540
rect 2160 5530 2190 5540
rect 2230 5530 2240 5540
rect 2390 5530 2420 5540
rect 2600 5530 2690 5540
rect 2850 5530 2860 5540
rect 2870 5530 2900 5540
rect 2920 5530 2940 5540
rect 2960 5530 2970 5540
rect 3220 5530 3250 5540
rect 3480 5530 3490 5540
rect 3500 5530 3510 5540
rect 3660 5530 3670 5540
rect 3800 5530 3810 5540
rect 4190 5530 4210 5540
rect 5110 5530 5120 5540
rect 5480 5530 5510 5540
rect 5610 5530 5690 5540
rect 5910 5530 5970 5540
rect 6170 5530 6240 5540
rect 6550 5530 6600 5540
rect 6610 5530 6620 5540
rect 6890 5530 6900 5540
rect 6950 5530 6970 5540
rect 7300 5530 7330 5540
rect 7370 5530 7380 5540
rect 7530 5530 7550 5540
rect 7610 5530 7650 5540
rect 7700 5530 7710 5540
rect 7790 5530 7800 5540
rect 7840 5530 7880 5540
rect 7940 5530 7960 5540
rect 8030 5530 8050 5540
rect 8100 5530 8110 5540
rect 8130 5530 8150 5540
rect 8770 5530 8780 5540
rect 8940 5530 8950 5540
rect 8990 5530 9000 5540
rect 510 5520 530 5530
rect 550 5520 570 5530
rect 590 5520 600 5530
rect 620 5520 640 5530
rect 1940 5520 1970 5530
rect 2160 5520 2190 5530
rect 2230 5520 2240 5530
rect 2390 5520 2420 5530
rect 2610 5520 2700 5530
rect 2840 5520 2900 5530
rect 2940 5520 2950 5530
rect 2970 5520 2980 5530
rect 3200 5520 3210 5530
rect 3220 5520 3250 5530
rect 3510 5520 3520 5530
rect 4160 5520 4170 5530
rect 4190 5520 4200 5530
rect 5110 5520 5130 5530
rect 5250 5520 5260 5530
rect 5470 5520 5480 5530
rect 5630 5520 5740 5530
rect 5920 5520 5960 5530
rect 6160 5520 6210 5530
rect 6550 5520 6600 5530
rect 6890 5520 6900 5530
rect 6950 5520 6970 5530
rect 7310 5520 7330 5530
rect 7350 5520 7360 5530
rect 7510 5520 7520 5530
rect 7620 5520 7650 5530
rect 7700 5520 7710 5530
rect 7840 5520 7880 5530
rect 7940 5520 7950 5530
rect 8030 5520 8050 5530
rect 8150 5520 8170 5530
rect 8860 5520 8870 5530
rect 8940 5520 8950 5530
rect 8990 5520 9000 5530
rect 480 5510 490 5520
rect 500 5510 540 5520
rect 590 5510 600 5520
rect 620 5510 640 5520
rect 930 5510 940 5520
rect 950 5510 960 5520
rect 1960 5510 1970 5520
rect 2160 5510 2190 5520
rect 2230 5510 2240 5520
rect 2270 5510 2280 5520
rect 2370 5510 2410 5520
rect 2600 5510 2620 5520
rect 2630 5510 2640 5520
rect 2650 5510 2700 5520
rect 2840 5510 2910 5520
rect 2940 5510 2990 5520
rect 3200 5510 3210 5520
rect 3220 5510 3250 5520
rect 3650 5510 3660 5520
rect 3730 5510 3740 5520
rect 3770 5510 3780 5520
rect 4150 5510 4160 5520
rect 4180 5510 4190 5520
rect 5100 5510 5110 5520
rect 5120 5510 5130 5520
rect 5250 5510 5260 5520
rect 5670 5510 5730 5520
rect 5920 5510 5960 5520
rect 6160 5510 6210 5520
rect 6540 5510 6600 5520
rect 6890 5510 6900 5520
rect 6940 5510 6960 5520
rect 7350 5510 7360 5520
rect 7380 5510 7390 5520
rect 7500 5510 7510 5520
rect 7640 5510 7650 5520
rect 7700 5510 7710 5520
rect 7840 5510 7880 5520
rect 7940 5510 7960 5520
rect 8040 5510 8060 5520
rect 8700 5510 8720 5520
rect 8750 5510 8760 5520
rect 8860 5510 8870 5520
rect 8910 5510 8920 5520
rect 8940 5510 8950 5520
rect 9060 5510 9080 5520
rect 430 5500 490 5510
rect 610 5500 620 5510
rect 2160 5500 2190 5510
rect 2230 5500 2240 5510
rect 2280 5500 2290 5510
rect 2370 5500 2410 5510
rect 2590 5500 2610 5510
rect 2660 5500 2690 5510
rect 2790 5500 2860 5510
rect 2870 5500 2910 5510
rect 2940 5500 3000 5510
rect 3200 5500 3210 5510
rect 3220 5500 3240 5510
rect 3650 5500 3660 5510
rect 3700 5500 3710 5510
rect 4150 5500 4160 5510
rect 4170 5500 4180 5510
rect 5680 5500 5730 5510
rect 5930 5500 5960 5510
rect 6160 5500 6200 5510
rect 6510 5500 6590 5510
rect 6920 5500 6930 5510
rect 6950 5500 6960 5510
rect 7380 5500 7390 5510
rect 7640 5500 7660 5510
rect 7700 5500 7720 5510
rect 7850 5500 7890 5510
rect 7940 5500 7960 5510
rect 8040 5500 8060 5510
rect 8740 5500 8760 5510
rect 8830 5500 8840 5510
rect 8850 5500 8870 5510
rect 400 5490 420 5500
rect 590 5490 610 5500
rect 1970 5490 1980 5500
rect 2160 5490 2180 5500
rect 2230 5490 2240 5500
rect 2290 5490 2300 5500
rect 2370 5490 2400 5500
rect 2590 5490 2600 5500
rect 2670 5490 2690 5500
rect 2730 5490 2740 5500
rect 2750 5490 2920 5500
rect 2940 5490 3010 5500
rect 3200 5490 3240 5500
rect 3290 5490 3300 5500
rect 3670 5490 3680 5500
rect 3730 5490 3750 5500
rect 4110 5490 4120 5500
rect 5520 5490 5540 5500
rect 5670 5490 5730 5500
rect 5760 5490 5790 5500
rect 5820 5490 5840 5500
rect 5930 5490 5960 5500
rect 6160 5490 6190 5500
rect 6460 5490 6540 5500
rect 6900 5490 6950 5500
rect 7260 5490 7270 5500
rect 7310 5490 7330 5500
rect 7550 5490 7590 5500
rect 7640 5490 7660 5500
rect 7750 5490 7760 5500
rect 7800 5490 7810 5500
rect 7850 5490 7890 5500
rect 7940 5490 7960 5500
rect 8630 5490 8650 5500
rect 8730 5490 8760 5500
rect 8840 5490 8870 5500
rect 8950 5490 8960 5500
rect 420 5480 430 5490
rect 550 5480 560 5490
rect 570 5480 580 5490
rect 600 5480 610 5490
rect 1970 5480 1980 5490
rect 2160 5480 2190 5490
rect 2230 5480 2240 5490
rect 2340 5480 2400 5490
rect 2490 5480 2500 5490
rect 2580 5480 2590 5490
rect 2680 5480 2690 5490
rect 2730 5480 3020 5490
rect 3200 5480 3240 5490
rect 3290 5480 3300 5490
rect 3620 5480 3650 5490
rect 4090 5480 4130 5490
rect 5100 5480 5120 5490
rect 5240 5480 5250 5490
rect 5520 5480 5760 5490
rect 5790 5480 5810 5490
rect 5820 5480 5840 5490
rect 5920 5480 5960 5490
rect 6150 5480 6180 5490
rect 6450 5480 6530 5490
rect 6900 5480 6960 5490
rect 7300 5480 7310 5490
rect 7320 5480 7340 5490
rect 7500 5480 7510 5490
rect 7560 5480 7590 5490
rect 7630 5480 7660 5490
rect 7800 5480 7810 5490
rect 7850 5480 7880 5490
rect 7940 5480 7960 5490
rect 8650 5480 8660 5490
rect 8680 5480 8690 5490
rect 8730 5480 8770 5490
rect 8850 5480 8870 5490
rect 8920 5480 8930 5490
rect 8940 5480 8960 5490
rect 9040 5480 9050 5490
rect 440 5470 460 5480
rect 570 5470 580 5480
rect 1970 5470 1980 5480
rect 2160 5470 2180 5480
rect 2230 5470 2240 5480
rect 2340 5470 2400 5480
rect 2570 5470 2600 5480
rect 2730 5470 3040 5480
rect 3190 5470 3240 5480
rect 3290 5470 3300 5480
rect 3570 5470 3580 5480
rect 3640 5470 3650 5480
rect 4090 5470 4130 5480
rect 4170 5470 4190 5480
rect 5090 5470 5110 5480
rect 5240 5470 5250 5480
rect 5500 5470 5540 5480
rect 5800 5470 5850 5480
rect 5930 5470 5960 5480
rect 6150 5470 6180 5480
rect 6440 5470 6530 5480
rect 6900 5470 6950 5480
rect 7260 5470 7280 5480
rect 7300 5470 7340 5480
rect 7390 5470 7400 5480
rect 7500 5470 7510 5480
rect 7550 5470 7580 5480
rect 7630 5470 7660 5480
rect 7740 5470 7750 5480
rect 7800 5470 7810 5480
rect 7850 5470 7870 5480
rect 7930 5470 7960 5480
rect 8610 5470 8620 5480
rect 8680 5470 8690 5480
rect 8730 5470 8740 5480
rect 8750 5470 8770 5480
rect 8860 5470 8880 5480
rect 8920 5470 8930 5480
rect 8940 5470 8960 5480
rect 9050 5470 9080 5480
rect 9120 5470 9130 5480
rect 1970 5460 1990 5470
rect 2160 5460 2190 5470
rect 2230 5460 2240 5470
rect 2350 5460 2390 5470
rect 2440 5460 2460 5470
rect 2570 5460 2600 5470
rect 2740 5460 2910 5470
rect 2930 5460 3040 5470
rect 3170 5460 3230 5470
rect 3280 5460 3300 5470
rect 3580 5460 3590 5470
rect 4110 5460 4120 5470
rect 5100 5460 5110 5470
rect 5240 5460 5250 5470
rect 5490 5460 5520 5470
rect 5930 5460 5960 5470
rect 6160 5460 6180 5470
rect 6440 5460 6530 5470
rect 6910 5460 6930 5470
rect 7250 5460 7280 5470
rect 7300 5460 7340 5470
rect 7500 5460 7510 5470
rect 7550 5460 7570 5470
rect 7630 5460 7670 5470
rect 7720 5460 7730 5470
rect 7930 5460 7960 5470
rect 8530 5460 8550 5470
rect 8610 5460 8620 5470
rect 8660 5460 8690 5470
rect 8740 5460 8770 5470
rect 8870 5460 8880 5470
rect 8950 5460 8960 5470
rect 9070 5460 9080 5470
rect 9120 5460 9130 5470
rect 440 5450 450 5460
rect 530 5450 540 5460
rect 580 5450 590 5460
rect 1970 5450 2010 5460
rect 2160 5450 2190 5460
rect 2230 5450 2240 5460
rect 2360 5450 2430 5460
rect 2590 5450 2630 5460
rect 2760 5450 2850 5460
rect 2910 5450 3010 5460
rect 3160 5450 3230 5460
rect 3280 5450 3300 5460
rect 4100 5450 4120 5460
rect 5470 5450 5500 5460
rect 5590 5450 5600 5460
rect 5650 5450 5670 5460
rect 5920 5450 5960 5460
rect 6160 5450 6180 5460
rect 6450 5450 6520 5460
rect 6900 5450 6940 5460
rect 7250 5450 7290 5460
rect 7300 5450 7340 5460
rect 7370 5450 7390 5460
rect 7620 5450 7670 5460
rect 7710 5450 7720 5460
rect 7920 5450 7960 5460
rect 8560 5450 8570 5460
rect 8610 5450 8620 5460
rect 8660 5450 8670 5460
rect 8680 5450 8700 5460
rect 8740 5450 8770 5460
rect 8950 5450 8970 5460
rect 9070 5450 9080 5460
rect 450 5440 460 5450
rect 1970 5440 2010 5450
rect 2160 5440 2190 5450
rect 2220 5440 2240 5450
rect 2360 5440 2390 5450
rect 2590 5440 2600 5450
rect 2780 5440 2860 5450
rect 2930 5440 3020 5450
rect 3160 5440 3230 5450
rect 3270 5440 3290 5450
rect 4100 5440 4110 5450
rect 5120 5440 5130 5450
rect 5450 5440 5480 5450
rect 5550 5440 5580 5450
rect 5650 5440 5680 5450
rect 5920 5440 5950 5450
rect 6160 5440 6180 5450
rect 6480 5440 6530 5450
rect 6900 5440 6920 5450
rect 7200 5440 7220 5450
rect 7240 5440 7290 5450
rect 7300 5440 7390 5450
rect 7510 5440 7520 5450
rect 7610 5440 7670 5450
rect 7810 5440 7820 5450
rect 7900 5440 7960 5450
rect 8510 5440 8520 5450
rect 8570 5440 8580 5450
rect 8680 5440 8700 5450
rect 8740 5440 8770 5450
rect 8820 5440 8830 5450
rect 8930 5440 8940 5450
rect 8960 5440 8970 5450
rect 450 5430 460 5440
rect 1970 5430 2020 5440
rect 2160 5430 2190 5440
rect 2230 5430 2240 5440
rect 2360 5430 2390 5440
rect 2620 5430 2640 5440
rect 2650 5430 2680 5440
rect 2730 5430 2740 5440
rect 2760 5430 2770 5440
rect 2790 5430 2820 5440
rect 2830 5430 2860 5440
rect 2950 5430 3000 5440
rect 3020 5430 3030 5440
rect 3050 5430 3060 5440
rect 3150 5430 3220 5440
rect 3270 5430 3290 5440
rect 3580 5430 3590 5440
rect 4100 5430 4110 5440
rect 4470 5430 4480 5440
rect 5120 5430 5130 5440
rect 5450 5430 5470 5440
rect 5530 5430 5570 5440
rect 5580 5430 5640 5440
rect 5920 5430 5950 5440
rect 6150 5430 6180 5440
rect 6510 5430 6600 5440
rect 6910 5430 6920 5440
rect 6940 5430 6950 5440
rect 7190 5430 7210 5440
rect 7250 5430 7290 5440
rect 7300 5430 7390 5440
rect 7510 5430 7520 5440
rect 7600 5430 7630 5440
rect 7640 5430 7670 5440
rect 7720 5430 7740 5440
rect 7810 5430 7820 5440
rect 7880 5430 7960 5440
rect 8510 5430 8520 5440
rect 8580 5430 8590 5440
rect 8620 5430 8630 5440
rect 8670 5430 8700 5440
rect 8750 5430 8780 5440
rect 8820 5430 8840 5440
rect 570 5420 580 5430
rect 1970 5420 2020 5430
rect 2050 5420 2060 5430
rect 2160 5420 2200 5430
rect 2230 5420 2240 5430
rect 2370 5420 2390 5430
rect 2660 5420 2700 5430
rect 2720 5420 2740 5430
rect 2770 5420 2820 5430
rect 2830 5420 2860 5430
rect 3030 5420 3040 5430
rect 3070 5420 3200 5430
rect 3580 5420 3590 5430
rect 4090 5420 4110 5430
rect 4320 5420 4340 5430
rect 4480 5420 4490 5430
rect 5090 5420 5110 5430
rect 5440 5420 5460 5430
rect 5510 5420 5550 5430
rect 5920 5420 5950 5430
rect 6160 5420 6180 5430
rect 6540 5420 6610 5430
rect 6910 5420 6930 5430
rect 6940 5420 6950 5430
rect 7260 5420 7290 5430
rect 7310 5420 7390 5430
rect 7510 5420 7520 5430
rect 7610 5420 7630 5430
rect 7640 5420 7670 5430
rect 7820 5420 7850 5430
rect 7860 5420 7870 5430
rect 7880 5420 7960 5430
rect 8390 5420 8400 5430
rect 8510 5420 8520 5430
rect 8590 5420 8600 5430
rect 8620 5420 8630 5430
rect 8670 5420 8700 5430
rect 8750 5420 8780 5430
rect 8830 5420 8850 5430
rect 440 5410 450 5420
rect 1970 5410 2020 5420
rect 2040 5410 2050 5420
rect 2160 5410 2200 5420
rect 2220 5410 2240 5420
rect 2360 5410 2390 5420
rect 2660 5410 2720 5420
rect 2730 5410 2810 5420
rect 2830 5410 2860 5420
rect 3040 5410 3050 5420
rect 3070 5410 3200 5420
rect 3580 5410 3590 5420
rect 5090 5410 5100 5420
rect 5110 5410 5120 5420
rect 5440 5410 5450 5420
rect 5500 5410 5530 5420
rect 5920 5410 5940 5420
rect 6160 5410 6180 5420
rect 6600 5410 6630 5420
rect 6910 5410 6960 5420
rect 7260 5410 7280 5420
rect 7300 5410 7400 5420
rect 7620 5410 7630 5420
rect 7640 5410 7680 5420
rect 7880 5410 7950 5420
rect 8360 5410 8370 5420
rect 8510 5410 8520 5420
rect 8600 5410 8610 5420
rect 8620 5410 8630 5420
rect 8670 5410 8700 5420
rect 8750 5410 8780 5420
rect 8830 5410 8860 5420
rect 490 5400 500 5410
rect 910 5400 920 5410
rect 1980 5400 2020 5410
rect 2040 5400 2060 5410
rect 2170 5400 2200 5410
rect 2220 5400 2240 5410
rect 2360 5400 2390 5410
rect 2660 5400 2720 5410
rect 2730 5400 2800 5410
rect 2820 5400 2870 5410
rect 3050 5400 3160 5410
rect 4500 5400 4520 5410
rect 5230 5400 5240 5410
rect 5430 5400 5440 5410
rect 5490 5400 5520 5410
rect 5920 5400 5940 5410
rect 6160 5400 6180 5410
rect 6620 5400 6660 5410
rect 6910 5400 6930 5410
rect 7300 5400 7400 5410
rect 7630 5400 7680 5410
rect 7890 5400 7960 5410
rect 8510 5400 8520 5410
rect 8610 5400 8640 5410
rect 8680 5400 8710 5410
rect 8750 5400 8790 5410
rect 8840 5400 8870 5410
rect 8940 5400 8950 5410
rect 9000 5400 9010 5410
rect 9510 5400 9520 5410
rect 500 5390 510 5400
rect 1990 5390 2040 5400
rect 2050 5390 2060 5400
rect 2170 5390 2200 5400
rect 2220 5390 2240 5400
rect 2360 5390 2380 5400
rect 2610 5390 2620 5400
rect 2680 5390 2760 5400
rect 2790 5390 2890 5400
rect 3090 5390 3130 5400
rect 4090 5390 4100 5400
rect 4500 5390 4510 5400
rect 4530 5390 4540 5400
rect 5090 5390 5100 5400
rect 5230 5390 5240 5400
rect 5400 5390 5430 5400
rect 5910 5390 5940 5400
rect 6160 5390 6180 5400
rect 6640 5390 6670 5400
rect 6910 5390 6930 5400
rect 7250 5390 7260 5400
rect 7300 5390 7410 5400
rect 7570 5390 7580 5400
rect 7650 5390 7680 5400
rect 7740 5390 7750 5400
rect 7890 5390 7900 5400
rect 7910 5390 7960 5400
rect 8490 5390 8500 5400
rect 8520 5390 8530 5400
rect 8620 5390 8640 5400
rect 8680 5390 8710 5400
rect 8760 5390 8790 5400
rect 8830 5390 8840 5400
rect 8860 5390 8880 5400
rect 9410 5390 9430 5400
rect 9540 5390 9550 5400
rect 470 5380 480 5390
rect 560 5380 570 5390
rect 1990 5380 2030 5390
rect 2080 5380 2090 5390
rect 2160 5380 2200 5390
rect 2220 5380 2240 5390
rect 2370 5380 2380 5390
rect 2610 5380 2640 5390
rect 2690 5380 2740 5390
rect 2840 5380 2870 5390
rect 2880 5380 2900 5390
rect 2910 5380 2920 5390
rect 3570 5380 3580 5390
rect 4530 5380 4540 5390
rect 5080 5380 5090 5390
rect 5230 5380 5240 5390
rect 5380 5380 5410 5390
rect 5450 5380 5460 5390
rect 5920 5380 5940 5390
rect 6160 5380 6180 5390
rect 6670 5380 6690 5390
rect 6910 5380 6930 5390
rect 7260 5380 7280 5390
rect 7300 5380 7410 5390
rect 7520 5380 7530 5390
rect 7570 5380 7590 5390
rect 7650 5380 7700 5390
rect 7710 5380 7720 5390
rect 7890 5380 7960 5390
rect 8490 5380 8500 5390
rect 8520 5380 8530 5390
rect 8570 5380 8580 5390
rect 8630 5380 8640 5390
rect 8680 5380 8710 5390
rect 8760 5380 8790 5390
rect 8830 5380 8840 5390
rect 8880 5380 8890 5390
rect 500 5370 530 5380
rect 1990 5370 2020 5380
rect 2080 5370 2110 5380
rect 2170 5370 2250 5380
rect 2360 5370 2380 5380
rect 2610 5370 2680 5380
rect 2710 5370 2720 5380
rect 2740 5370 2750 5380
rect 2880 5370 2940 5380
rect 4530 5370 4540 5380
rect 5390 5370 5400 5380
rect 5410 5370 5440 5380
rect 5910 5370 5940 5380
rect 6160 5370 6180 5380
rect 6670 5370 6700 5380
rect 6910 5370 6920 5380
rect 7260 5370 7280 5380
rect 7300 5370 7310 5380
rect 7330 5370 7410 5380
rect 7510 5370 7530 5380
rect 7570 5370 7600 5380
rect 7900 5370 7970 5380
rect 8230 5370 8240 5380
rect 8270 5370 8280 5380
rect 8390 5370 8400 5380
rect 8440 5370 8450 5380
rect 8490 5370 8500 5380
rect 8680 5370 8710 5380
rect 8760 5370 8800 5380
rect 8880 5370 8890 5380
rect 9570 5370 9580 5380
rect 340 5360 350 5370
rect 530 5360 540 5370
rect 1990 5360 2020 5370
rect 2030 5360 2040 5370
rect 2080 5360 2110 5370
rect 2170 5360 2250 5370
rect 2360 5360 2390 5370
rect 2610 5360 2710 5370
rect 2910 5360 2930 5370
rect 4080 5360 4100 5370
rect 5420 5360 5430 5370
rect 5720 5360 5750 5370
rect 5900 5360 5930 5370
rect 6160 5360 6180 5370
rect 6680 5360 6720 5370
rect 6910 5360 6930 5370
rect 7320 5360 7420 5370
rect 7520 5360 7530 5370
rect 7570 5360 7620 5370
rect 7920 5360 7970 5370
rect 8440 5360 8450 5370
rect 8580 5360 8600 5370
rect 8690 5360 8720 5370
rect 8760 5360 8800 5370
rect 8910 5360 8930 5370
rect 9310 5360 9350 5370
rect 440 5350 450 5360
rect 540 5350 550 5360
rect 2000 5350 2050 5360
rect 2060 5350 2080 5360
rect 2110 5350 2120 5360
rect 2170 5350 2250 5360
rect 2360 5350 2390 5360
rect 2620 5350 2720 5360
rect 4080 5350 4100 5360
rect 5390 5350 5410 5360
rect 5470 5350 5520 5360
rect 5530 5350 5550 5360
rect 5860 5350 5930 5360
rect 6160 5350 6180 5360
rect 6700 5350 6720 5360
rect 6910 5350 6930 5360
rect 7330 5350 7400 5360
rect 7520 5350 7530 5360
rect 7570 5350 7580 5360
rect 7900 5350 7970 5360
rect 8140 5350 8150 5360
rect 8350 5350 8360 5360
rect 8420 5350 8430 5360
rect 8580 5350 8600 5360
rect 8690 5350 8720 5360
rect 8780 5350 8800 5360
rect 270 5340 300 5350
rect 380 5340 410 5350
rect 540 5340 560 5350
rect 2000 5340 2090 5350
rect 2120 5340 2130 5350
rect 2170 5340 2250 5350
rect 2370 5340 2390 5350
rect 2600 5340 2610 5350
rect 2620 5340 2720 5350
rect 4110 5340 4120 5350
rect 5370 5340 5400 5350
rect 5420 5340 5440 5350
rect 5580 5340 5590 5350
rect 5620 5340 5670 5350
rect 5850 5340 5930 5350
rect 6170 5340 6200 5350
rect 6380 5340 6390 5350
rect 6710 5340 6730 5350
rect 7250 5340 7260 5350
rect 7310 5340 7320 5350
rect 7340 5340 7370 5350
rect 7530 5340 7540 5350
rect 7560 5340 7570 5350
rect 7900 5340 7970 5350
rect 8130 5340 8140 5350
rect 8220 5340 8230 5350
rect 8290 5340 8300 5350
rect 8480 5340 8490 5350
rect 8530 5340 8540 5350
rect 8580 5340 8600 5350
rect 8700 5340 8720 5350
rect 9370 5340 9380 5350
rect 9410 5340 9420 5350
rect 9570 5340 9580 5350
rect 260 5330 270 5340
rect 330 5330 350 5340
rect 2000 5330 2090 5340
rect 2110 5330 2130 5340
rect 2170 5330 2250 5340
rect 2360 5330 2390 5340
rect 2480 5330 2520 5340
rect 2600 5330 2720 5340
rect 5110 5330 5130 5340
rect 5610 5330 5700 5340
rect 5860 5330 5870 5340
rect 5900 5330 5920 5340
rect 6170 5330 6190 5340
rect 6370 5330 6400 5340
rect 6720 5330 6740 5340
rect 7290 5330 7360 5340
rect 7900 5330 7980 5340
rect 8080 5330 8100 5340
rect 8110 5330 8130 5340
rect 8220 5330 8230 5340
rect 8470 5330 8480 5340
rect 8530 5330 8540 5340
rect 8580 5330 8590 5340
rect 8610 5330 8620 5340
rect 8690 5330 8730 5340
rect 9260 5330 9270 5340
rect 9330 5330 9340 5340
rect 9450 5330 9460 5340
rect 240 5320 250 5330
rect 300 5320 310 5330
rect 2000 5320 2060 5330
rect 2080 5320 2090 5330
rect 2110 5320 2130 5330
rect 2170 5320 2250 5330
rect 2370 5320 2390 5330
rect 2480 5320 2520 5330
rect 2600 5320 2650 5330
rect 2660 5320 2730 5330
rect 3550 5320 3560 5330
rect 4650 5320 4680 5330
rect 5150 5320 5160 5330
rect 5220 5320 5230 5330
rect 5660 5320 5750 5330
rect 5860 5320 5870 5330
rect 6170 5320 6190 5330
rect 6730 5320 6750 5330
rect 7280 5320 7310 5330
rect 7320 5320 7360 5330
rect 7890 5320 7980 5330
rect 8060 5320 8070 5330
rect 8110 5320 8130 5330
rect 8170 5320 8180 5330
rect 8220 5320 8230 5330
rect 8300 5320 8310 5330
rect 8360 5320 8370 5330
rect 8530 5320 8540 5330
rect 8580 5320 8590 5330
rect 8620 5320 8630 5330
rect 8690 5320 8710 5330
rect 8720 5320 8730 5330
rect 8760 5320 8770 5330
rect 9300 5320 9310 5330
rect 230 5310 240 5320
rect 290 5310 300 5320
rect 570 5310 580 5320
rect 2000 5310 2070 5320
rect 2100 5310 2130 5320
rect 2170 5310 2250 5320
rect 2370 5310 2390 5320
rect 2470 5310 2530 5320
rect 2600 5310 2630 5320
rect 2680 5310 2740 5320
rect 4590 5310 4600 5320
rect 4650 5310 4680 5320
rect 4700 5310 4720 5320
rect 5130 5310 5150 5320
rect 5700 5310 5770 5320
rect 5790 5310 5800 5320
rect 5810 5310 5860 5320
rect 6170 5310 6200 5320
rect 6460 5310 6490 5320
rect 6590 5310 6640 5320
rect 6740 5310 6790 5320
rect 7270 5310 7360 5320
rect 7900 5310 7980 5320
rect 8010 5310 8030 5320
rect 8120 5310 8130 5320
rect 8170 5310 8180 5320
rect 8220 5310 8230 5320
rect 8470 5310 8480 5320
rect 8540 5310 8550 5320
rect 8630 5310 8640 5320
rect 8740 5310 8750 5320
rect 9420 5310 9430 5320
rect 9520 5310 9530 5320
rect 9600 5310 9610 5320
rect 220 5300 230 5310
rect 240 5300 260 5310
rect 560 5300 570 5310
rect 2010 5300 2080 5310
rect 2090 5300 2140 5310
rect 2180 5300 2250 5310
rect 2370 5300 2390 5310
rect 2460 5300 2530 5310
rect 2600 5300 2630 5310
rect 2660 5300 2740 5310
rect 3540 5300 3550 5310
rect 4680 5300 4700 5310
rect 5130 5300 5150 5310
rect 5170 5300 5180 5310
rect 5210 5300 5220 5310
rect 5700 5300 5840 5310
rect 6180 5300 6200 5310
rect 6390 5300 6400 5310
rect 6430 5300 6480 5310
rect 6540 5300 6570 5310
rect 6640 5300 6680 5310
rect 6770 5300 6790 5310
rect 7270 5300 7350 5310
rect 7910 5300 7980 5310
rect 8040 5300 8060 5310
rect 8120 5300 8130 5310
rect 8170 5300 8180 5310
rect 8200 5300 8230 5310
rect 8310 5300 8320 5310
rect 8410 5300 8420 5310
rect 8540 5300 8550 5310
rect 8640 5300 8650 5310
rect 9330 5300 9340 5310
rect 9350 5300 9360 5310
rect 9610 5300 9620 5310
rect 230 5290 240 5300
rect 300 5290 320 5300
rect 2010 5290 2080 5300
rect 2090 5290 2150 5300
rect 2180 5290 2250 5300
rect 2370 5290 2400 5300
rect 2460 5290 2490 5300
rect 2520 5290 2570 5300
rect 2600 5290 2610 5300
rect 2630 5290 2640 5300
rect 2660 5290 2680 5300
rect 2700 5290 2760 5300
rect 5100 5290 5120 5300
rect 5140 5290 5150 5300
rect 5160 5290 5180 5300
rect 5210 5290 5220 5300
rect 5700 5290 5850 5300
rect 6180 5290 6210 5300
rect 6380 5290 6400 5300
rect 6460 5290 6480 5300
rect 6490 5290 6520 5300
rect 6640 5290 6670 5300
rect 6680 5290 6700 5300
rect 6770 5290 6780 5300
rect 7260 5290 7340 5300
rect 7910 5290 7990 5300
rect 8040 5290 8060 5300
rect 8180 5290 8200 5300
rect 8210 5290 8230 5300
rect 8410 5290 8430 5300
rect 8640 5290 8660 5300
rect 8670 5290 8680 5300
rect 9260 5290 9270 5300
rect 9370 5290 9380 5300
rect 9460 5290 9470 5300
rect 9570 5290 9580 5300
rect 200 5280 220 5290
rect 310 5280 330 5290
rect 2010 5280 2080 5290
rect 2090 5280 2150 5290
rect 2190 5280 2250 5290
rect 2370 5280 2400 5290
rect 2460 5280 2480 5290
rect 2530 5280 2580 5290
rect 2640 5280 2680 5290
rect 2700 5280 2800 5290
rect 3530 5280 3540 5290
rect 5080 5280 5100 5290
rect 5150 5280 5180 5290
rect 5690 5280 5850 5290
rect 6190 5280 6220 5290
rect 6290 5280 6300 5290
rect 6380 5280 6460 5290
rect 6630 5280 6670 5290
rect 6730 5280 6740 5290
rect 6760 5280 6780 5290
rect 7250 5280 7330 5290
rect 7910 5280 8000 5290
rect 8050 5280 8060 5290
rect 8180 5280 8190 5290
rect 8200 5280 8230 5290
rect 8270 5280 8280 5290
rect 8320 5280 8330 5290
rect 8420 5280 8430 5290
rect 8440 5280 8450 5290
rect 8500 5280 8510 5290
rect 9120 5280 9130 5290
rect 9160 5280 9170 5290
rect 9380 5280 9390 5290
rect 9430 5280 9440 5290
rect 9550 5280 9560 5290
rect 9610 5280 9620 5290
rect 190 5270 200 5280
rect 300 5270 340 5280
rect 2010 5270 2160 5280
rect 2190 5270 2250 5280
rect 2370 5270 2410 5280
rect 2450 5270 2480 5280
rect 2560 5270 2590 5280
rect 2650 5270 2680 5280
rect 2700 5270 2810 5280
rect 5090 5270 5160 5280
rect 5170 5270 5180 5280
rect 5210 5270 5220 5280
rect 5630 5270 5660 5280
rect 5680 5270 5860 5280
rect 6190 5270 6310 5280
rect 6330 5270 6430 5280
rect 6620 5270 6660 5280
rect 6760 5270 6780 5280
rect 7260 5270 7330 5280
rect 7910 5270 8000 5280
rect 8050 5270 8060 5280
rect 8180 5270 8190 5280
rect 8200 5270 8230 5280
rect 8270 5270 8280 5280
rect 8370 5270 8380 5280
rect 8580 5270 8590 5280
rect 9080 5270 9090 5280
rect 9280 5270 9290 5280
rect 9340 5270 9350 5280
rect 9430 5270 9440 5280
rect 9850 5270 9860 5280
rect 9870 5270 9880 5280
rect 320 5260 350 5270
rect 2020 5260 2160 5270
rect 2180 5260 2240 5270
rect 2380 5260 2410 5270
rect 2440 5260 2470 5270
rect 2570 5260 2600 5270
rect 2700 5260 2730 5270
rect 2750 5260 2820 5270
rect 2860 5260 2870 5270
rect 5070 5260 5080 5270
rect 5100 5260 5180 5270
rect 5210 5260 5220 5270
rect 5630 5260 5840 5270
rect 6200 5260 6300 5270
rect 6330 5260 6430 5270
rect 6560 5260 6570 5270
rect 6590 5260 6620 5270
rect 7230 5260 7250 5270
rect 7270 5260 7340 5270
rect 7430 5260 7440 5270
rect 7940 5260 8010 5270
rect 8050 5260 8060 5270
rect 8180 5260 8190 5270
rect 8200 5260 8230 5270
rect 8270 5260 8290 5270
rect 8330 5260 8340 5270
rect 8370 5260 8380 5270
rect 8450 5260 8470 5270
rect 8510 5260 8520 5270
rect 8940 5260 8950 5270
rect 9090 5260 9100 5270
rect 9390 5260 9400 5270
rect 9520 5260 9540 5270
rect 340 5250 350 5260
rect 360 5250 370 5260
rect 2020 5250 2170 5260
rect 2180 5250 2250 5260
rect 2380 5250 2470 5260
rect 2590 5250 2610 5260
rect 2700 5250 2730 5260
rect 2740 5250 2750 5260
rect 2790 5250 2820 5260
rect 2850 5250 2890 5260
rect 5070 5250 5080 5260
rect 5100 5250 5180 5260
rect 5190 5250 5220 5260
rect 5550 5250 5600 5260
rect 5630 5250 5730 5260
rect 5750 5250 5810 5260
rect 6210 5250 6230 5260
rect 6240 5250 6340 5260
rect 6370 5250 6450 5260
rect 6530 5250 6600 5260
rect 7270 5250 7340 5260
rect 7930 5250 8010 5260
rect 8180 5250 8190 5260
rect 8220 5250 8230 5260
rect 8270 5250 8280 5260
rect 8370 5250 8380 5260
rect 8420 5250 8430 5260
rect 8470 5250 8480 5260
rect 8510 5250 8520 5260
rect 9130 5250 9140 5260
rect 9170 5250 9180 5260
rect 9470 5250 9480 5260
rect 370 5240 380 5250
rect 600 5240 620 5250
rect 2020 5240 2160 5250
rect 2180 5240 2250 5250
rect 2380 5240 2470 5250
rect 2610 5240 2620 5250
rect 2690 5240 2740 5250
rect 2790 5240 2830 5250
rect 2840 5240 2890 5250
rect 3510 5240 3520 5250
rect 5070 5240 5080 5250
rect 5140 5240 5220 5250
rect 5590 5240 5700 5250
rect 5750 5240 5780 5250
rect 6240 5240 6250 5250
rect 6270 5240 6370 5250
rect 6380 5240 6390 5250
rect 6410 5240 6420 5250
rect 6430 5240 6580 5250
rect 7270 5240 7330 5250
rect 7940 5240 8010 5250
rect 8180 5240 8190 5250
rect 8220 5240 8230 5250
rect 8420 5240 8430 5250
rect 8930 5240 8940 5250
rect 9040 5240 9050 5250
rect 9740 5240 9750 5250
rect 9800 5240 9810 5250
rect 9910 5240 9920 5250
rect 430 5230 440 5240
rect 2030 5230 2160 5240
rect 2190 5230 2250 5240
rect 2380 5230 2470 5240
rect 2630 5230 2640 5240
rect 2650 5230 2660 5240
rect 2690 5230 2730 5240
rect 2790 5230 2810 5240
rect 2830 5230 2840 5240
rect 2870 5230 2900 5240
rect 5060 5230 5210 5240
rect 5620 5230 5730 5240
rect 6300 5230 6310 5240
rect 6330 5230 6380 5240
rect 6450 5230 6460 5240
rect 6480 5230 6540 5240
rect 6560 5230 6600 5240
rect 7280 5230 7340 5240
rect 7930 5230 8020 5240
rect 8180 5230 8190 5240
rect 8220 5230 8230 5240
rect 8370 5230 8390 5240
rect 8420 5230 8430 5240
rect 8930 5230 8940 5240
rect 9130 5230 9150 5240
rect 9330 5230 9350 5240
rect 9850 5230 9860 5240
rect 9920 5230 9930 5240
rect 430 5220 450 5230
rect 2030 5220 2110 5230
rect 2120 5220 2160 5230
rect 2190 5220 2250 5230
rect 2380 5220 2470 5230
rect 2650 5220 2660 5230
rect 2690 5220 2720 5230
rect 2790 5220 2810 5230
rect 2820 5220 2830 5230
rect 2880 5220 2900 5230
rect 5060 5220 5070 5230
rect 5110 5220 5130 5230
rect 5140 5220 5210 5230
rect 6340 5220 6390 5230
rect 6550 5220 6590 5230
rect 7310 5220 7340 5230
rect 7420 5220 7430 5230
rect 7930 5220 8020 5230
rect 8100 5220 8110 5230
rect 8180 5220 8190 5230
rect 8200 5220 8220 5230
rect 8350 5220 8360 5230
rect 8380 5220 8400 5230
rect 8930 5220 8940 5230
rect 9380 5220 9390 5230
rect 9820 5220 9830 5230
rect 9960 5220 9970 5230
rect 650 5210 670 5220
rect 2030 5210 2100 5220
rect 2120 5210 2180 5220
rect 2210 5210 2250 5220
rect 2380 5210 2460 5220
rect 2670 5210 2710 5220
rect 2800 5210 2820 5220
rect 2890 5210 2910 5220
rect 5060 5210 5080 5220
rect 5110 5210 5120 5220
rect 5140 5210 5200 5220
rect 6360 5210 6470 5220
rect 6480 5210 6560 5220
rect 7260 5210 7290 5220
rect 7330 5210 7340 5220
rect 7420 5210 7430 5220
rect 7940 5210 8020 5220
rect 8100 5210 8120 5220
rect 8180 5210 8190 5220
rect 8200 5210 8220 5220
rect 8280 5210 8290 5220
rect 8300 5210 8310 5220
rect 8350 5210 8360 5220
rect 8930 5210 8940 5220
rect 9050 5210 9060 5220
rect 9090 5210 9100 5220
rect 9750 5210 9760 5220
rect 9970 5210 9980 5220
rect 2030 5200 2090 5210
rect 2120 5200 2190 5210
rect 2210 5200 2250 5210
rect 2380 5200 2460 5210
rect 2790 5200 2810 5210
rect 2890 5200 2910 5210
rect 5060 5200 5080 5210
rect 5100 5200 5120 5210
rect 5140 5200 5160 5210
rect 5170 5200 5200 5210
rect 6440 5200 6460 5210
rect 6510 5200 6520 5210
rect 7230 5200 7280 5210
rect 7290 5200 7320 5210
rect 7330 5200 7350 5210
rect 7950 5200 8010 5210
rect 8020 5200 8030 5210
rect 8100 5200 8120 5210
rect 8200 5200 8220 5210
rect 8260 5200 8270 5210
rect 8310 5200 8320 5210
rect 8830 5200 8840 5210
rect 8930 5200 8940 5210
rect 9000 5200 9010 5210
rect 9110 5200 9120 5210
rect 9320 5200 9330 5210
rect 9340 5200 9350 5210
rect 9990 5200 9990 5210
rect 640 5190 660 5200
rect 680 5190 690 5200
rect 2030 5190 2090 5200
rect 2130 5190 2250 5200
rect 2390 5190 2460 5200
rect 2670 5190 2680 5200
rect 2790 5190 2810 5200
rect 2890 5190 2910 5200
rect 5070 5190 5080 5200
rect 5100 5190 5120 5200
rect 5140 5190 5160 5200
rect 5170 5190 5190 5200
rect 7260 5190 7280 5200
rect 7290 5190 7350 5200
rect 7950 5190 8010 5200
rect 8100 5190 8120 5200
rect 8190 5190 8220 5200
rect 8260 5190 8270 5200
rect 8690 5190 8700 5200
rect 8710 5190 8720 5200
rect 8870 5190 8880 5200
rect 8930 5190 8940 5200
rect 9560 5190 9590 5200
rect 9930 5190 9940 5200
rect 660 5180 670 5190
rect 2040 5180 2100 5190
rect 2110 5180 2120 5190
rect 2130 5180 2250 5190
rect 2380 5180 2460 5190
rect 2680 5180 2700 5190
rect 2780 5180 2810 5190
rect 2880 5180 2910 5190
rect 2940 5180 2990 5190
rect 5170 5180 5200 5190
rect 7290 5180 7350 5190
rect 7960 5180 8010 5190
rect 8100 5180 8130 5190
rect 8190 5180 8230 5190
rect 8660 5180 8670 5190
rect 8840 5180 8850 5190
rect 8930 5180 8940 5190
rect 8970 5180 8980 5190
rect 9060 5180 9070 5190
rect 9520 5180 9530 5190
rect 9600 5180 9610 5190
rect 9800 5180 9810 5190
rect 9870 5180 9880 5190
rect 640 5170 660 5180
rect 2040 5170 2100 5180
rect 2110 5170 2190 5180
rect 2210 5170 2250 5180
rect 2390 5170 2460 5180
rect 2690 5170 2700 5180
rect 2760 5170 2790 5180
rect 2860 5170 2910 5180
rect 2930 5170 2990 5180
rect 5070 5170 5080 5180
rect 5170 5170 5200 5180
rect 7290 5170 7340 5180
rect 7950 5170 8010 5180
rect 8030 5170 8040 5180
rect 8110 5170 8130 5180
rect 8230 5170 8250 5180
rect 8750 5170 8760 5180
rect 8840 5170 8850 5180
rect 9150 5170 9160 5180
rect 9610 5170 9620 5180
rect 130 5160 140 5170
rect 610 5160 620 5170
rect 650 5160 690 5170
rect 2040 5160 2180 5170
rect 2230 5160 2260 5170
rect 2390 5160 2420 5170
rect 2430 5160 2460 5170
rect 2700 5160 2720 5170
rect 2850 5160 2900 5170
rect 2920 5160 2990 5170
rect 5170 5160 5200 5170
rect 7290 5160 7330 5170
rect 7960 5160 8010 5170
rect 8030 5160 8040 5170
rect 8120 5160 8140 5170
rect 8180 5160 8190 5170
rect 8790 5160 8810 5170
rect 8880 5160 8890 5170
rect 8970 5160 8980 5170
rect 9450 5160 9460 5170
rect 9500 5160 9510 5170
rect 9570 5160 9580 5170
rect 9710 5160 9720 5170
rect 9750 5160 9760 5170
rect 9810 5160 9820 5170
rect 9970 5160 9980 5170
rect 130 5150 140 5160
rect 580 5150 590 5160
rect 610 5150 620 5160
rect 660 5150 680 5160
rect 2050 5150 2190 5160
rect 2230 5150 2260 5160
rect 2400 5150 2410 5160
rect 2430 5150 2460 5160
rect 2710 5150 2730 5160
rect 2850 5150 2900 5160
rect 2920 5150 3000 5160
rect 3460 5150 3470 5160
rect 5160 5150 5200 5160
rect 7310 5150 7340 5160
rect 7960 5150 8010 5160
rect 8090 5150 8100 5160
rect 8140 5150 8150 5160
rect 8170 5150 8180 5160
rect 9070 5150 9080 5160
rect 9410 5150 9420 5160
rect 9540 5150 9550 5160
rect 9620 5150 9630 5160
rect 9810 5150 9820 5160
rect 9840 5150 9850 5160
rect 9880 5150 9890 5160
rect 130 5140 140 5150
rect 570 5140 610 5150
rect 2040 5140 2200 5150
rect 2220 5140 2260 5150
rect 2430 5140 2460 5150
rect 2730 5140 2740 5150
rect 2810 5140 2820 5150
rect 2850 5140 2890 5150
rect 2910 5140 2990 5150
rect 5100 5140 5110 5150
rect 5150 5140 5180 5150
rect 5190 5140 5200 5150
rect 7310 5140 7340 5150
rect 7970 5140 8000 5150
rect 8040 5140 8050 5150
rect 8090 5140 8100 5150
rect 8640 5140 8660 5150
rect 9540 5140 9550 5150
rect 9720 5140 9730 5150
rect 9810 5140 9820 5150
rect 9880 5140 9890 5150
rect 530 5130 540 5140
rect 570 5130 610 5140
rect 2060 5130 2110 5140
rect 2120 5130 2200 5140
rect 2220 5130 2260 5140
rect 2420 5130 2460 5140
rect 2840 5130 2890 5140
rect 2910 5130 2980 5140
rect 3470 5130 3480 5140
rect 5110 5130 5120 5140
rect 5150 5130 5170 5140
rect 5190 5130 5210 5140
rect 7310 5130 7330 5140
rect 7970 5130 8010 5140
rect 8510 5130 8520 5140
rect 8760 5130 8770 5140
rect 8810 5130 8820 5140
rect 8850 5130 8860 5140
rect 9450 5130 9460 5140
rect 9590 5130 9600 5140
rect 9810 5130 9820 5140
rect 130 5120 150 5130
rect 520 5120 560 5130
rect 570 5120 580 5130
rect 590 5120 610 5130
rect 2060 5120 2110 5130
rect 2130 5120 2200 5130
rect 2230 5120 2260 5130
rect 2420 5120 2460 5130
rect 2750 5120 2770 5130
rect 2910 5120 2960 5130
rect 3440 5120 3450 5130
rect 5140 5120 5180 5130
rect 5200 5120 5210 5130
rect 7310 5120 7330 5130
rect 7970 5120 8010 5130
rect 8440 5120 8450 5130
rect 8660 5120 8670 5130
rect 8920 5120 8930 5130
rect 9020 5120 9040 5130
rect 9290 5120 9300 5130
rect 9330 5120 9340 5130
rect 9420 5120 9430 5130
rect 9510 5120 9520 5130
rect 9760 5120 9770 5130
rect 9910 5120 9920 5130
rect 130 5110 150 5120
rect 520 5110 580 5120
rect 600 5110 620 5120
rect 2070 5110 2130 5120
rect 2140 5110 2200 5120
rect 2230 5110 2260 5120
rect 2410 5110 2420 5120
rect 2430 5110 2470 5120
rect 2770 5110 2780 5120
rect 2910 5110 2960 5120
rect 3460 5110 3490 5120
rect 5130 5110 5140 5120
rect 5150 5110 5180 5120
rect 5200 5110 5210 5120
rect 7310 5110 7320 5120
rect 7970 5110 8010 5120
rect 8420 5110 8430 5120
rect 8660 5110 8670 5120
rect 8800 5110 8810 5120
rect 8890 5110 8900 5120
rect 9260 5110 9270 5120
rect 9630 5110 9640 5120
rect 9770 5110 9800 5120
rect 9840 5110 9850 5120
rect 140 5100 150 5110
rect 520 5100 580 5110
rect 2080 5100 2140 5110
rect 2150 5100 2200 5110
rect 2230 5100 2260 5110
rect 2410 5100 2460 5110
rect 2730 5100 2750 5110
rect 2780 5100 2810 5110
rect 2940 5100 2970 5110
rect 3450 5100 3460 5110
rect 5150 5100 5170 5110
rect 5200 5100 5210 5110
rect 7300 5100 7310 5110
rect 7970 5100 8010 5110
rect 8480 5100 8490 5110
rect 8770 5100 8780 5110
rect 8800 5100 8810 5110
rect 8930 5100 8940 5110
rect 8950 5100 8960 5110
rect 9230 5100 9240 5110
rect 9330 5100 9340 5110
rect 9600 5100 9610 5110
rect 140 5090 160 5100
rect 470 5090 540 5100
rect 550 5090 580 5100
rect 2090 5090 2140 5100
rect 2150 5090 2220 5100
rect 2230 5090 2270 5100
rect 2410 5090 2420 5100
rect 2430 5090 2470 5100
rect 2720 5090 2750 5100
rect 2790 5090 2830 5100
rect 3420 5090 3430 5100
rect 5150 5090 5170 5100
rect 7300 5090 7320 5100
rect 7980 5090 8010 5100
rect 8330 5090 8370 5100
rect 9310 5090 9320 5100
rect 9370 5090 9380 5100
rect 9420 5090 9430 5100
rect 9470 5090 9480 5100
rect 9520 5090 9530 5100
rect 9550 5090 9560 5100
rect 9600 5090 9610 5100
rect 140 5080 160 5090
rect 480 5080 500 5090
rect 520 5080 590 5090
rect 2100 5080 2220 5090
rect 2230 5080 2270 5090
rect 2430 5080 2460 5090
rect 2710 5080 2720 5090
rect 2790 5080 2860 5090
rect 5160 5080 5170 5090
rect 7300 5080 7310 5090
rect 7990 5080 8020 5090
rect 8290 5080 8300 5090
rect 8420 5080 8430 5090
rect 8670 5080 8680 5090
rect 8810 5080 8820 5090
rect 8880 5080 8890 5090
rect 9140 5080 9150 5090
rect 9230 5080 9240 5090
rect 9790 5080 9800 5090
rect 140 5070 170 5080
rect 450 5070 480 5080
rect 540 5070 600 5080
rect 2080 5070 2280 5080
rect 2430 5070 2480 5080
rect 2680 5070 2710 5080
rect 2790 5070 2860 5080
rect 5150 5070 5170 5080
rect 5200 5070 5220 5080
rect 7300 5070 7310 5080
rect 7990 5070 8030 5080
rect 8280 5070 8290 5080
rect 8460 5070 8470 5080
rect 8810 5070 8820 5080
rect 9270 5070 9280 5080
rect 40 5060 70 5070
rect 150 5060 170 5070
rect 370 5060 430 5070
rect 480 5060 490 5070
rect 500 5060 610 5070
rect 2080 5060 2230 5070
rect 2240 5060 2280 5070
rect 2420 5060 2500 5070
rect 2670 5060 2700 5070
rect 2740 5060 2870 5070
rect 5150 5060 5180 5070
rect 5200 5060 5220 5070
rect 7300 5060 7310 5070
rect 7990 5060 8030 5070
rect 8400 5060 8410 5070
rect 9190 5060 9200 5070
rect 9270 5060 9280 5070
rect 9310 5060 9320 5070
rect 9560 5060 9570 5070
rect 9590 5060 9600 5070
rect 30 5050 50 5060
rect 160 5050 170 5060
rect 310 5050 320 5060
rect 360 5050 380 5060
rect 2090 5050 2230 5060
rect 2240 5050 2270 5060
rect 2430 5050 2520 5060
rect 2650 5050 2700 5060
rect 2720 5050 2890 5060
rect 3310 5050 3320 5060
rect 3390 5050 3400 5060
rect 5160 5050 5180 5060
rect 5200 5050 5220 5060
rect 7990 5050 8030 5060
rect 8240 5050 8250 5060
rect 8280 5050 8290 5060
rect 8320 5050 8330 5060
rect 8400 5050 8410 5060
rect 8430 5050 8440 5060
rect 8510 5050 8520 5060
rect 8710 5050 8720 5060
rect 9050 5050 9060 5060
rect 9170 5050 9180 5060
rect 9530 5050 9540 5060
rect 40 5040 50 5050
rect 300 5040 320 5050
rect 360 5040 380 5050
rect 2100 5040 2270 5050
rect 2430 5040 2520 5050
rect 2600 5040 2630 5050
rect 2640 5040 2860 5050
rect 2870 5040 2890 5050
rect 2940 5040 2960 5050
rect 3390 5040 3410 5050
rect 5160 5040 5180 5050
rect 5200 5040 5220 5050
rect 7300 5040 7310 5050
rect 7360 5040 7370 5050
rect 7980 5040 8030 5050
rect 8160 5040 8170 5050
rect 8250 5040 8260 5050
rect 8280 5040 8290 5050
rect 8320 5040 8330 5050
rect 8400 5040 8410 5050
rect 8430 5040 8440 5050
rect 8490 5040 8500 5050
rect 9030 5040 9040 5050
rect 9110 5040 9140 5050
rect 170 5030 180 5040
rect 340 5030 380 5040
rect 2110 5030 2280 5040
rect 2440 5030 2520 5040
rect 2650 5030 2830 5040
rect 2870 5030 2890 5040
rect 2940 5030 2960 5040
rect 3400 5030 3410 5040
rect 5160 5030 5180 5040
rect 5210 5030 5230 5040
rect 7350 5030 7400 5040
rect 7980 5030 8030 5040
rect 8150 5030 8160 5040
rect 8260 5030 8270 5040
rect 8280 5030 8290 5040
rect 8320 5030 8330 5040
rect 8470 5030 8480 5040
rect 8690 5030 8700 5040
rect 8970 5030 8980 5040
rect 9030 5030 9040 5040
rect 9280 5030 9290 5040
rect 9390 5030 9400 5040
rect 9420 5030 9430 5040
rect 9480 5030 9490 5040
rect 9590 5030 9600 5040
rect 170 5020 180 5030
rect 190 5020 200 5030
rect 350 5020 380 5030
rect 2110 5020 2280 5030
rect 2440 5020 2540 5030
rect 2580 5020 2620 5030
rect 2650 5020 2830 5030
rect 2940 5020 2960 5030
rect 5160 5020 5180 5030
rect 5200 5020 5230 5030
rect 7310 5020 7320 5030
rect 7400 5020 7440 5030
rect 7990 5020 8030 5030
rect 8140 5020 8150 5030
rect 8200 5020 8230 5030
rect 8260 5020 8270 5030
rect 8330 5020 8340 5030
rect 8470 5020 8480 5030
rect 9030 5020 9040 5030
rect 9320 5020 9330 5030
rect 9430 5020 9450 5030
rect 9500 5020 9510 5030
rect 170 5010 200 5020
rect 380 5010 400 5020
rect 2120 5010 2300 5020
rect 2450 5010 2500 5020
rect 2510 5010 2550 5020
rect 2570 5010 2820 5020
rect 2940 5010 2950 5020
rect 3360 5010 3370 5020
rect 3390 5010 3400 5020
rect 5160 5010 5180 5020
rect 5740 5010 5780 5020
rect 7450 5010 7460 5020
rect 7990 5010 8040 5020
rect 8140 5010 8150 5020
rect 8440 5010 8450 5020
rect 8490 5010 8500 5020
rect 8910 5010 8920 5020
rect 9070 5010 9080 5020
rect 9140 5010 9150 5020
rect 180 5000 190 5010
rect 210 5000 220 5010
rect 370 5000 410 5010
rect 2120 5000 2300 5010
rect 2450 5000 2760 5010
rect 3360 5000 3370 5010
rect 3390 5000 3410 5010
rect 4160 5000 4170 5010
rect 4180 5000 4190 5010
rect 5170 5000 5180 5010
rect 5710 5000 5780 5010
rect 6330 5000 6340 5010
rect 6350 5000 6360 5010
rect 7310 5000 7320 5010
rect 7990 5000 8000 5010
rect 8030 5000 8050 5010
rect 8130 5000 8150 5010
rect 8220 5000 8230 5010
rect 8290 5000 8300 5010
rect 8440 5000 8450 5010
rect 9290 5000 9300 5010
rect 200 4990 210 5000
rect 220 4990 230 5000
rect 370 4990 410 5000
rect 2120 4990 2310 5000
rect 2440 4990 2590 5000
rect 2600 4990 2760 5000
rect 3360 4990 3370 5000
rect 3390 4990 3400 5000
rect 5180 4990 5190 5000
rect 5700 4990 5750 5000
rect 5760 4990 5780 5000
rect 6340 4990 6370 5000
rect 7310 4990 7320 5000
rect 7990 4990 8000 5000
rect 8070 4990 8080 5000
rect 8120 4990 8130 5000
rect 8270 4990 8280 5000
rect 210 4980 240 4990
rect 370 4980 420 4990
rect 2130 4980 2310 4990
rect 2450 4980 2760 4990
rect 3360 4980 3390 4990
rect 4210 4980 4220 4990
rect 4290 4980 4330 4990
rect 4510 4980 4560 4990
rect 5200 4980 5220 4990
rect 5660 4980 5670 4990
rect 5690 4980 5720 4990
rect 5760 4980 5770 4990
rect 6340 4980 6390 4990
rect 7310 4980 7320 4990
rect 7990 4980 8000 4990
rect 8050 4980 8070 4990
rect 8120 4980 8150 4990
rect 8270 4980 8280 4990
rect 8340 4980 8350 4990
rect 8400 4980 8410 4990
rect 8510 4980 8520 4990
rect 8760 4980 8770 4990
rect 9040 4980 9050 4990
rect 9150 4980 9160 4990
rect 220 4970 260 4980
rect 370 4970 420 4980
rect 2140 4970 2320 4980
rect 2460 4970 2680 4980
rect 2690 4970 2760 4980
rect 3340 4970 3350 4980
rect 3370 4970 3390 4980
rect 4020 4970 4030 4980
rect 4040 4970 4050 4980
rect 4060 4970 4070 4980
rect 4270 4970 4280 4980
rect 4310 4970 4320 4980
rect 4520 4970 4530 4980
rect 4560 4970 4570 4980
rect 4580 4970 4590 4980
rect 5200 4970 5230 4980
rect 5640 4970 5720 4980
rect 5750 4970 5770 4980
rect 6340 4970 6400 4980
rect 7990 4970 8000 4980
rect 8060 4970 8070 4980
rect 8140 4970 8150 4980
rect 8190 4970 8200 4980
rect 8230 4970 8240 4980
rect 8270 4970 8280 4980
rect 8300 4970 8310 4980
rect 8340 4970 8360 4980
rect 8460 4970 8480 4980
rect 8840 4970 8850 4980
rect 8880 4970 8890 4980
rect 8940 4970 8950 4980
rect 9300 4970 9310 4980
rect 9660 4970 9670 4980
rect 240 4960 280 4970
rect 380 4960 420 4970
rect 2150 4960 2330 4970
rect 2460 4960 2640 4970
rect 2690 4960 2700 4970
rect 2710 4960 2760 4970
rect 3350 4960 3360 4970
rect 3380 4960 3390 4970
rect 4000 4960 4010 4970
rect 4060 4960 4070 4970
rect 4090 4960 4100 4970
rect 4310 4960 4340 4970
rect 5200 4960 5230 4970
rect 5620 4960 5700 4970
rect 5740 4960 5770 4970
rect 6340 4960 6350 4970
rect 6370 4960 6410 4970
rect 7320 4960 7330 4970
rect 7850 4960 7860 4970
rect 7990 4960 8000 4970
rect 8060 4960 8070 4970
rect 8130 4960 8160 4970
rect 8200 4960 8210 4970
rect 8230 4960 8240 4970
rect 8300 4960 8310 4970
rect 8850 4960 8860 4970
rect 8880 4960 8890 4970
rect 8950 4960 8960 4970
rect 9080 4960 9090 4970
rect 9190 4960 9200 4970
rect 9630 4960 9640 4970
rect 260 4950 270 4960
rect 280 4950 300 4960
rect 390 4950 420 4960
rect 2160 4950 2340 4960
rect 2460 4950 2640 4960
rect 3350 4950 3360 4960
rect 3370 4950 3380 4960
rect 4060 4950 4070 4960
rect 4350 4950 4360 4960
rect 4380 4950 4390 4960
rect 4600 4950 4610 4960
rect 4620 4950 4650 4960
rect 5200 4950 5230 4960
rect 5610 4950 5690 4960
rect 5730 4950 5760 4960
rect 6340 4950 6350 4960
rect 6380 4950 6430 4960
rect 7320 4950 7330 4960
rect 7840 4950 7850 4960
rect 7930 4950 7940 4960
rect 7990 4950 8000 4960
rect 8150 4950 8160 4960
rect 8230 4950 8240 4960
rect 8340 4950 8350 4960
rect 8380 4950 8390 4960
rect 8400 4950 8410 4960
rect 9050 4950 9060 4960
rect 9160 4950 9170 4960
rect 9610 4950 9620 4960
rect 180 4940 190 4950
rect 220 4940 250 4950
rect 260 4940 280 4950
rect 330 4940 400 4950
rect 2170 4940 2270 4950
rect 2320 4940 2340 4950
rect 2460 4940 2650 4950
rect 3230 4940 3240 4950
rect 3360 4940 3380 4950
rect 4000 4940 4010 4950
rect 4420 4940 4430 4950
rect 4490 4940 4520 4950
rect 4660 4940 4670 4950
rect 4700 4940 4710 4950
rect 5200 4940 5240 4950
rect 5600 4940 5670 4950
rect 5730 4940 5750 4950
rect 6140 4940 6190 4950
rect 6340 4940 6350 4950
rect 6400 4940 6440 4950
rect 7320 4940 7330 4950
rect 7830 4940 7840 4950
rect 7990 4940 8010 4950
rect 8130 4940 8140 4950
rect 8220 4940 8230 4950
rect 8620 4940 8630 4950
rect 8820 4940 8830 4950
rect 8890 4940 8900 4950
rect 9160 4940 9170 4950
rect 9660 4940 9670 4950
rect 110 4930 260 4940
rect 320 4930 360 4940
rect 2170 4930 2190 4940
rect 2210 4930 2260 4940
rect 2320 4930 2340 4940
rect 2470 4930 2640 4940
rect 3330 4930 3340 4940
rect 3360 4930 3370 4940
rect 4060 4930 4070 4940
rect 4360 4930 4370 4940
rect 4440 4930 4450 4940
rect 4510 4930 4520 4940
rect 4540 4930 4550 4940
rect 4740 4930 4760 4940
rect 5060 4930 5070 4940
rect 5210 4930 5240 4940
rect 5590 4930 5650 4940
rect 5720 4930 5740 4940
rect 5790 4930 5860 4940
rect 5880 4930 5900 4940
rect 5930 4930 5940 4940
rect 6140 4930 6200 4940
rect 6230 4930 6300 4940
rect 6330 4930 6350 4940
rect 6400 4930 6450 4940
rect 7880 4930 7900 4940
rect 7940 4930 7950 4940
rect 7990 4930 8010 4940
rect 8130 4930 8140 4940
rect 8160 4930 8170 4940
rect 8270 4930 8280 4940
rect 8320 4930 8340 4940
rect 8600 4930 8610 4940
rect 8700 4930 8710 4940
rect 8740 4930 8750 4940
rect 8820 4930 8830 4940
rect 8930 4930 8940 4940
rect 8980 4930 9000 4940
rect 9020 4930 9030 4940
rect 9140 4930 9150 4940
rect 9610 4930 9620 4940
rect 80 4920 220 4930
rect 320 4920 380 4930
rect 2210 4920 2250 4930
rect 2330 4920 2350 4930
rect 2470 4920 2660 4930
rect 3330 4920 3340 4930
rect 3360 4920 3370 4930
rect 3990 4920 4000 4930
rect 4050 4920 4070 4930
rect 4120 4920 4140 4930
rect 4190 4920 4200 4930
rect 4350 4920 4360 4930
rect 4390 4920 4400 4930
rect 4470 4920 4480 4930
rect 4580 4920 4600 4930
rect 4790 4920 4810 4930
rect 5050 4920 5060 4930
rect 5210 4920 5240 4930
rect 5580 4920 5650 4930
rect 5720 4920 5740 4930
rect 5790 4920 5830 4930
rect 5910 4920 5930 4930
rect 5960 4920 5970 4930
rect 6130 4920 6280 4930
rect 6290 4920 6340 4930
rect 6410 4920 6450 4930
rect 7820 4920 7830 4930
rect 7890 4920 7900 4930
rect 7940 4920 7950 4930
rect 8000 4920 8010 4930
rect 8160 4920 8170 4930
rect 8260 4920 8270 4930
rect 8740 4920 8750 4930
rect 8810 4920 8820 4930
rect 8930 4920 8940 4930
rect 8980 4920 8990 4930
rect 9130 4920 9140 4930
rect 9460 4920 9470 4930
rect 9650 4920 9660 4930
rect 60 4910 90 4920
rect 150 4910 190 4920
rect 330 4910 410 4920
rect 2240 4910 2250 4920
rect 2330 4910 2370 4920
rect 2480 4910 2490 4920
rect 2500 4910 2650 4920
rect 3300 4910 3310 4920
rect 3920 4910 3930 4920
rect 3970 4910 3980 4920
rect 3990 4910 4000 4920
rect 4010 4910 4020 4920
rect 4110 4910 4120 4920
rect 4180 4910 4190 4920
rect 4490 4910 4500 4920
rect 4580 4910 4590 4920
rect 4630 4910 4660 4920
rect 5040 4910 5060 4920
rect 5210 4910 5240 4920
rect 5570 4910 5630 4920
rect 5710 4910 5740 4920
rect 5790 4910 5820 4920
rect 5930 4910 5980 4920
rect 6060 4910 6080 4920
rect 6090 4910 6220 4920
rect 6420 4910 6470 4920
rect 7320 4910 7330 4920
rect 7690 4910 7700 4920
rect 7710 4910 7720 4920
rect 7820 4910 7830 4920
rect 7860 4910 7870 4920
rect 7890 4910 7900 4920
rect 7940 4910 7950 4920
rect 8000 4910 8010 4920
rect 8170 4910 8180 4920
rect 8250 4910 8260 4920
rect 8510 4910 8520 4920
rect 8600 4910 8610 4920
rect 8640 4910 8650 4920
rect 8900 4910 8910 4920
rect 9060 4910 9070 4920
rect 9450 4910 9460 4920
rect 9680 4910 9690 4920
rect 9710 4910 9720 4920
rect 40 4900 70 4910
rect 380 4900 420 4910
rect 2200 4900 2220 4910
rect 2330 4900 2370 4910
rect 2510 4900 2640 4910
rect 3300 4900 3310 4910
rect 3320 4900 3330 4910
rect 3350 4900 3370 4910
rect 3480 4900 3490 4910
rect 3900 4900 3910 4910
rect 3970 4900 3980 4910
rect 3990 4900 4000 4910
rect 4080 4900 4090 4910
rect 4520 4900 4540 4910
rect 4550 4900 4570 4910
rect 4620 4900 4630 4910
rect 4710 4900 4720 4910
rect 5020 4900 5050 4910
rect 5210 4900 5240 4910
rect 5550 4900 5610 4910
rect 5700 4900 5730 4910
rect 5790 4900 5820 4910
rect 5950 4900 6140 4910
rect 6170 4900 6200 4910
rect 6430 4900 6470 4910
rect 7760 4900 7770 4910
rect 7800 4900 7810 4910
rect 7820 4900 7830 4910
rect 7900 4900 7910 4910
rect 8000 4900 8010 4910
rect 8100 4900 8110 4910
rect 8140 4900 8150 4910
rect 8180 4900 8200 4910
rect 8220 4900 8230 4910
rect 8640 4900 8650 4910
rect 8970 4900 8980 4910
rect 9070 4900 9080 4910
rect 9390 4900 9410 4910
rect 9490 4900 9500 4910
rect 9530 4900 9540 4910
rect 30 4890 50 4900
rect 2200 4890 2220 4900
rect 2240 4890 2250 4900
rect 2340 4890 2380 4900
rect 2520 4890 2580 4900
rect 2590 4890 2640 4900
rect 3320 4890 3330 4900
rect 3350 4890 3370 4900
rect 3910 4890 3920 4900
rect 3930 4890 3940 4900
rect 3960 4890 3980 4900
rect 4010 4890 4020 4900
rect 4060 4890 4070 4900
rect 4490 4890 4500 4900
rect 4540 4890 4550 4900
rect 4600 4890 4670 4900
rect 4750 4890 4780 4900
rect 4830 4890 4840 4900
rect 5210 4890 5240 4900
rect 5540 4890 5600 4900
rect 5690 4890 5730 4900
rect 5790 4890 5820 4900
rect 5960 4890 6130 4900
rect 6440 4890 6480 4900
rect 7800 4890 7810 4900
rect 7900 4890 7910 4900
rect 8000 4890 8020 4900
rect 8060 4890 8070 4900
rect 8100 4890 8110 4900
rect 8140 4890 8150 4900
rect 8660 4890 8670 4900
rect 8750 4890 8760 4900
rect 8940 4890 8950 4900
rect 9000 4890 9010 4900
rect 9380 4890 9390 4900
rect 9450 4890 9460 4900
rect 9530 4890 9540 4900
rect 9620 4890 9630 4900
rect 10 4880 40 4890
rect 490 4880 500 4890
rect 2240 4880 2250 4890
rect 2360 4880 2370 4890
rect 2520 4880 2660 4890
rect 3320 4880 3330 4890
rect 3360 4880 3370 4890
rect 3740 4880 3750 4890
rect 3930 4880 3940 4890
rect 3960 4880 3970 4890
rect 4040 4880 4050 4890
rect 4180 4880 4190 4890
rect 4550 4880 4580 4890
rect 4790 4880 4800 4890
rect 4810 4880 4830 4890
rect 4870 4880 4880 4890
rect 5210 4880 5220 4890
rect 5520 4880 5590 4890
rect 5680 4880 5740 4890
rect 5800 4880 5830 4890
rect 5970 4880 6050 4890
rect 6090 4880 6120 4890
rect 6440 4880 6500 4890
rect 7330 4880 7350 4890
rect 7900 4880 7910 4890
rect 8000 4880 8020 4890
rect 8060 4880 8070 4890
rect 8520 4880 8540 4890
rect 8580 4880 8590 4890
rect 8790 4880 8800 4890
rect 9310 4880 9330 4890
rect 9350 4880 9360 4890
rect 9380 4880 9390 4890
rect 0 4870 30 4880
rect 2240 4870 2250 4880
rect 2350 4870 2370 4880
rect 2530 4870 2540 4880
rect 2550 4870 2660 4880
rect 3320 4870 3330 4880
rect 3360 4870 3370 4880
rect 3700 4870 3710 4880
rect 3920 4870 3940 4880
rect 4020 4870 4030 4880
rect 4830 4870 4840 4880
rect 5210 4870 5220 4880
rect 5230 4870 5240 4880
rect 5510 4870 5590 4880
rect 5680 4870 5750 4880
rect 5800 4870 5850 4880
rect 5980 4870 6030 4880
rect 6450 4870 6510 4880
rect 7220 4870 7240 4880
rect 7330 4870 7340 4880
rect 7760 4870 7770 4880
rect 7870 4870 7880 4880
rect 7950 4870 7960 4880
rect 8000 4870 8020 4880
rect 8060 4870 8070 4880
rect 8580 4870 8590 4880
rect 8610 4870 8620 4880
rect 8940 4870 8950 4880
rect 9520 4870 9530 4880
rect 0 4860 30 4870
rect 40 4860 70 4870
rect 2350 4860 2370 4870
rect 2570 4860 2580 4870
rect 2610 4860 2660 4870
rect 3320 4860 3330 4870
rect 3340 4860 3350 4870
rect 3370 4860 3380 4870
rect 3840 4860 3850 4870
rect 3860 4860 3870 4870
rect 5500 4860 5580 4870
rect 5680 4860 5750 4870
rect 5810 4860 5850 4870
rect 5910 4860 5920 4870
rect 5980 4860 6010 4870
rect 6370 4860 6380 4870
rect 6460 4860 6520 4870
rect 7330 4860 7360 4870
rect 7690 4860 7700 4870
rect 7770 4860 7780 4870
rect 7810 4860 7820 4870
rect 7830 4860 7840 4870
rect 7870 4860 7880 4870
rect 7900 4860 7910 4870
rect 7950 4860 7960 4870
rect 8010 4860 8030 4870
rect 8060 4860 8070 4870
rect 8340 4860 8350 4870
rect 8540 4860 8550 4870
rect 8580 4860 8590 4870
rect 8670 4860 8680 4870
rect 8760 4860 8770 4870
rect 8790 4860 8800 4870
rect 8820 4860 8830 4870
rect 8930 4860 8940 4870
rect 9080 4860 9090 4870
rect 9460 4860 9470 4870
rect 0 4850 80 4860
rect 350 4850 370 4860
rect 2350 4850 2380 4860
rect 2610 4850 2670 4860
rect 3340 4850 3360 4860
rect 3370 4850 3380 4860
rect 3750 4850 3770 4860
rect 3820 4850 3830 4860
rect 3990 4850 4000 4860
rect 4930 4850 4940 4860
rect 4950 4850 4960 4860
rect 5480 4850 5570 4860
rect 5670 4850 5740 4860
rect 5830 4850 5960 4860
rect 6360 4850 6370 4860
rect 6460 4850 6530 4860
rect 7330 4850 7360 4860
rect 7380 4850 7390 4860
rect 7810 4850 7820 4860
rect 7830 4850 7840 4860
rect 7890 4850 7910 4860
rect 8020 4850 8040 4860
rect 8050 4850 8060 4860
rect 8290 4850 8300 4860
rect 8470 4850 8480 4860
rect 8540 4850 8550 4860
rect 8760 4850 8770 4860
rect 8870 4850 8880 4860
rect 9390 4850 9400 4860
rect 9460 4850 9470 4860
rect 9560 4850 9570 4860
rect 9630 4850 9640 4860
rect 9670 4850 9680 4860
rect 9740 4850 9750 4860
rect 0 4840 80 4850
rect 90 4840 100 4850
rect 2350 4840 2380 4850
rect 2630 4840 2680 4850
rect 3160 4840 3170 4850
rect 3250 4840 3260 4850
rect 3330 4840 3340 4850
rect 3370 4840 3380 4850
rect 3710 4840 3720 4850
rect 3730 4840 3770 4850
rect 3800 4840 3820 4850
rect 4910 4840 4940 4850
rect 4960 4840 4970 4850
rect 5190 4840 5200 4850
rect 5470 4840 5560 4850
rect 5670 4840 5740 4850
rect 5840 4840 5990 4850
rect 6470 4840 6530 4850
rect 7830 4840 7840 4850
rect 7940 4840 7950 4850
rect 8050 4840 8060 4850
rect 8620 4840 8630 4850
rect 8650 4840 8660 4850
rect 9070 4840 9080 4850
rect 9500 4840 9510 4850
rect 9550 4840 9560 4850
rect 9690 4840 9710 4850
rect 0 4830 170 4840
rect 2350 4830 2390 4840
rect 2630 4830 2690 4840
rect 3150 4830 3160 4840
rect 3240 4830 3260 4840
rect 3360 4830 3370 4840
rect 3380 4830 3390 4840
rect 3710 4830 3720 4840
rect 3750 4830 3810 4840
rect 3940 4830 3950 4840
rect 3970 4830 3980 4840
rect 5190 4830 5220 4840
rect 5460 4830 5550 4840
rect 5660 4830 5730 4840
rect 5850 4830 5980 4840
rect 6370 4830 6380 4840
rect 6480 4830 6530 4840
rect 7280 4830 7290 4840
rect 7700 4830 7710 4840
rect 7830 4830 7840 4840
rect 8200 4830 8210 4840
rect 8620 4830 8630 4840
rect 8730 4830 8740 4840
rect 8790 4830 8800 4840
rect 9060 4830 9070 4840
rect 9500 4830 9520 4840
rect 9550 4830 9560 4840
rect 9600 4830 9610 4840
rect 40 4820 200 4830
rect 2360 4820 2390 4830
rect 2650 4820 2670 4830
rect 2680 4820 2710 4830
rect 3150 4820 3160 4830
rect 3250 4820 3270 4830
rect 3360 4820 3370 4830
rect 3380 4820 3390 4830
rect 3570 4820 3580 4830
rect 3750 4820 3770 4830
rect 3780 4820 3800 4830
rect 3930 4820 3940 4830
rect 4920 4820 4930 4830
rect 4990 4820 5000 4830
rect 5190 4820 5240 4830
rect 5450 4820 5550 4830
rect 5670 4820 5730 4830
rect 5870 4820 5980 4830
rect 6370 4820 6380 4830
rect 6480 4820 6550 4830
rect 7340 4820 7350 4830
rect 7740 4820 7750 4830
rect 7760 4820 7770 4830
rect 7820 4820 7830 4830
rect 7920 4820 7930 4830
rect 8310 4820 8320 4830
rect 9470 4820 9480 4830
rect 9730 4820 9740 4830
rect 0 4810 220 4820
rect 280 4810 290 4820
rect 2360 4810 2390 4820
rect 2670 4810 2710 4820
rect 3140 4810 3150 4820
rect 3220 4810 3260 4820
rect 3360 4810 3380 4820
rect 3560 4810 3570 4820
rect 3740 4810 3760 4820
rect 3790 4810 3800 4820
rect 3940 4810 3950 4820
rect 4960 4810 4970 4820
rect 5000 4810 5010 4820
rect 5170 4810 5210 4820
rect 5460 4810 5520 4820
rect 5660 4810 5700 4820
rect 5890 4810 5980 4820
rect 6490 4810 6580 4820
rect 7740 4810 7750 4820
rect 7820 4810 7830 4820
rect 7860 4810 7870 4820
rect 8130 4810 8150 4820
rect 8230 4810 8240 4820
rect 8480 4810 8490 4820
rect 8520 4810 8530 4820
rect 8730 4810 8740 4820
rect 9050 4810 9060 4820
rect 9400 4810 9410 4820
rect 9570 4810 9580 4820
rect 9640 4810 9650 4820
rect 9700 4810 9710 4820
rect 0 4800 130 4810
rect 150 4800 230 4810
rect 2370 4800 2390 4810
rect 2430 4800 2450 4810
rect 2670 4800 2750 4810
rect 3130 4800 3140 4810
rect 3270 4800 3280 4810
rect 3370 4800 3380 4810
rect 3550 4800 3560 4810
rect 3910 4800 3930 4810
rect 4960 4800 4970 4810
rect 5180 4800 5210 4810
rect 5430 4800 5510 4810
rect 5660 4800 5700 4810
rect 5910 4800 5920 4810
rect 5940 4800 5980 4810
rect 6250 4800 6290 4810
rect 6320 4800 6360 4810
rect 6510 4800 6580 4810
rect 7780 4800 7790 4810
rect 7820 4800 7830 4810
rect 9000 4800 9010 4810
rect 9040 4800 9050 4810
rect 9330 4800 9340 4810
rect 9510 4800 9520 4810
rect 0 4790 110 4800
rect 140 4790 150 4800
rect 160 4790 170 4800
rect 180 4790 210 4800
rect 2390 4790 2420 4800
rect 2430 4790 2440 4800
rect 2680 4790 2760 4800
rect 3130 4790 3140 4800
rect 3360 4790 3370 4800
rect 3550 4790 3560 4800
rect 3890 4790 3910 4800
rect 4940 4790 4950 4800
rect 5420 4790 5500 4800
rect 5650 4790 5690 4800
rect 5950 4790 5990 4800
rect 6230 4790 6360 4800
rect 6510 4790 6580 4800
rect 8030 4790 8070 4800
rect 8240 4790 8250 4800
rect 8270 4790 8280 4800
rect 8370 4790 8380 4800
rect 9030 4790 9050 4800
rect 9440 4790 9450 4800
rect 0 4780 110 4790
rect 130 4780 180 4790
rect 2390 4780 2420 4790
rect 2690 4780 2800 4790
rect 3120 4780 3130 4790
rect 3340 4780 3350 4790
rect 3540 4780 3550 4790
rect 5030 4780 5040 4790
rect 5410 4780 5490 4790
rect 5640 4780 5690 4790
rect 5960 4780 5990 4790
rect 6210 4780 6380 4790
rect 6520 4780 6590 4790
rect 7710 4780 7720 4790
rect 8010 4780 8020 4790
rect 8200 4780 8210 4790
rect 8240 4780 8250 4790
rect 8490 4780 8500 4790
rect 8930 4780 8940 4790
rect 0 4770 140 4780
rect 2420 4770 2430 4780
rect 2440 4770 2450 4780
rect 2690 4770 2820 4780
rect 3110 4770 3120 4780
rect 3240 4770 3250 4780
rect 3270 4770 3280 4780
rect 3340 4770 3350 4780
rect 3530 4770 3550 4780
rect 3590 4770 3600 4780
rect 3860 4770 3880 4780
rect 5410 4770 5480 4780
rect 5630 4770 5670 4780
rect 5970 4770 6010 4780
rect 6130 4770 6140 4780
rect 6190 4770 6390 4780
rect 6530 4770 6620 4780
rect 6630 4770 6640 4780
rect 7720 4770 7740 4780
rect 8100 4770 8110 4780
rect 8190 4770 8210 4780
rect 8390 4770 8400 4780
rect 8910 4770 8920 4780
rect 9000 4770 9010 4780
rect 9340 4770 9350 4780
rect 0 4760 160 4770
rect 2420 4760 2430 4770
rect 2450 4760 2460 4770
rect 2500 4760 2510 4770
rect 2720 4760 2830 4770
rect 3100 4760 3110 4770
rect 3340 4760 3350 4770
rect 3530 4760 3540 4770
rect 3840 4760 3870 4770
rect 5070 4760 5080 4770
rect 5410 4760 5470 4770
rect 5620 4760 5670 4770
rect 5970 4760 6030 4770
rect 6110 4760 6400 4770
rect 6540 4760 6640 4770
rect 7350 4760 7360 4770
rect 7990 4760 8000 4770
rect 8100 4760 8130 4770
rect 8200 4760 8210 4770
rect 8830 4760 8850 4770
rect 0 4750 150 4760
rect 2450 4750 2480 4760
rect 2490 4750 2510 4760
rect 2730 4750 2830 4760
rect 3100 4750 3120 4760
rect 3340 4750 3350 4760
rect 3520 4750 3550 4760
rect 3860 4750 3870 4760
rect 5080 4750 5090 4760
rect 5410 4750 5470 4760
rect 5610 4750 5660 4760
rect 5980 4750 6410 4760
rect 6550 4750 6640 4760
rect 7380 4750 7390 4760
rect 7900 4750 7940 4760
rect 8110 4750 8130 4760
rect 8870 4750 8880 4760
rect 9310 4750 9320 4760
rect 0 4740 150 4750
rect 2450 4740 2470 4750
rect 2480 4740 2510 4750
rect 2720 4740 2850 4750
rect 3090 4740 3110 4750
rect 3350 4740 3360 4750
rect 3530 4740 3550 4750
rect 3830 4740 3840 4750
rect 5090 4740 5100 4750
rect 5400 4740 5470 4750
rect 5600 4740 5650 4750
rect 5990 4740 6420 4750
rect 6560 4740 6640 4750
rect 7360 4740 7380 4750
rect 7950 4740 7960 4750
rect 7980 4740 7990 4750
rect 8030 4740 8060 4750
rect 8110 4740 8130 4750
rect 8250 4740 8260 4750
rect 8290 4740 8300 4750
rect 8350 4740 8360 4750
rect 8790 4740 8800 4750
rect 8880 4740 8890 4750
rect 9990 4740 9990 4750
rect 0 4730 160 4740
rect 2450 4730 2480 4740
rect 2500 4730 2550 4740
rect 2710 4730 2850 4740
rect 3260 4730 3270 4740
rect 3530 4730 3540 4740
rect 3560 4730 3580 4740
rect 5110 4730 5120 4740
rect 5400 4730 5470 4740
rect 5600 4730 5640 4740
rect 6020 4730 6310 4740
rect 6320 4730 6430 4740
rect 6570 4730 6640 4740
rect 7980 4730 7990 4740
rect 8030 4730 8060 4740
rect 8170 4730 8180 4740
rect 8840 4730 8850 4740
rect 8990 4730 9000 4740
rect 0 4720 150 4730
rect 2450 4720 2480 4730
rect 2500 4720 2550 4730
rect 2710 4720 2860 4730
rect 2990 4720 3010 4730
rect 3060 4720 3080 4730
rect 3530 4720 3540 4730
rect 3550 4720 3560 4730
rect 5120 4720 5130 4730
rect 5400 4720 5470 4730
rect 5600 4720 5640 4730
rect 6030 4720 6240 4730
rect 6250 4720 6270 4730
rect 6300 4720 6440 4730
rect 6570 4720 6640 4730
rect 7980 4720 7990 4730
rect 8030 4720 8070 4730
rect 8130 4720 8140 4730
rect 8170 4720 8180 4730
rect 8190 4720 8200 4730
rect 8780 4720 8790 4730
rect 8920 4720 8930 4730
rect 9000 4720 9010 4730
rect 0 4710 150 4720
rect 2460 4710 2470 4720
rect 2530 4710 2560 4720
rect 2620 4710 2650 4720
rect 2710 4710 2850 4720
rect 2980 4710 3010 4720
rect 3060 4710 3070 4720
rect 3350 4710 3360 4720
rect 3530 4710 3550 4720
rect 5130 4710 5140 4720
rect 5210 4710 5220 4720
rect 5400 4710 5460 4720
rect 5600 4710 5650 4720
rect 6030 4710 6070 4720
rect 6080 4710 6230 4720
rect 6320 4710 6440 4720
rect 6580 4710 6640 4720
rect 7360 4710 7370 4720
rect 7740 4710 7750 4720
rect 7850 4710 7860 4720
rect 7980 4710 7990 4720
rect 8030 4710 8070 4720
rect 8200 4710 8210 4720
rect 8260 4710 8270 4720
rect 8290 4710 8300 4720
rect 8360 4710 8370 4720
rect 8640 4710 8650 4720
rect 8660 4710 8670 4720
rect 8960 4710 8970 4720
rect 0 4700 160 4710
rect 2540 4700 2580 4710
rect 2640 4700 2840 4710
rect 2850 4700 2890 4710
rect 2960 4700 3020 4710
rect 3060 4700 3090 4710
rect 3350 4700 3360 4710
rect 3520 4700 3540 4710
rect 5100 4700 5110 4710
rect 5140 4700 5150 4710
rect 5200 4700 5220 4710
rect 5400 4700 5460 4710
rect 5610 4700 5650 4710
rect 6040 4700 6050 4710
rect 6100 4700 6200 4710
rect 6320 4700 6460 4710
rect 6580 4700 6650 4710
rect 7820 4700 7830 4710
rect 7890 4700 7900 4710
rect 8030 4700 8040 4710
rect 8060 4700 8080 4710
rect 8110 4700 8120 4710
rect 8210 4700 8220 4710
rect 8260 4700 8270 4710
rect 8310 4700 8340 4710
rect 8780 4700 8790 4710
rect 8960 4700 8970 4710
rect 9280 4700 9290 4710
rect 0 4690 150 4700
rect 2450 4690 2460 4700
rect 2540 4690 2630 4700
rect 2670 4690 2720 4700
rect 2730 4690 2750 4700
rect 2780 4690 2830 4700
rect 2860 4690 2880 4700
rect 2960 4690 3000 4700
rect 3350 4690 3360 4700
rect 5390 4690 5470 4700
rect 5630 4690 5660 4700
rect 6140 4690 6180 4700
rect 6320 4690 6460 4700
rect 6570 4690 6640 4700
rect 7370 4690 7380 4700
rect 7850 4690 7860 4700
rect 7900 4690 7920 4700
rect 7940 4690 7950 4700
rect 8060 4690 8080 4700
rect 8140 4690 8150 4700
rect 8220 4690 8230 4700
rect 8570 4690 8580 4700
rect 8780 4690 8790 4700
rect 8860 4690 8870 4700
rect 9820 4690 9830 4700
rect 0 4680 140 4690
rect 2450 4680 2470 4690
rect 2550 4680 2600 4690
rect 2800 4680 2820 4690
rect 2960 4680 3000 4690
rect 3150 4680 3160 4690
rect 3350 4680 3370 4690
rect 5390 4680 5470 4690
rect 5630 4680 5680 4690
rect 6320 4680 6460 4690
rect 6570 4680 6640 4690
rect 7380 4680 7390 4690
rect 7630 4680 7650 4690
rect 7690 4680 7700 4690
rect 7770 4680 7790 4690
rect 7830 4680 7860 4690
rect 7960 4680 7970 4690
rect 7990 4680 8000 4690
rect 8030 4680 8040 4690
rect 8060 4680 8080 4690
rect 8180 4680 8190 4690
rect 8900 4680 8910 4690
rect 8930 4680 8940 4690
rect 9270 4680 9280 4690
rect 9810 4680 9820 4690
rect 0 4670 130 4680
rect 2620 4670 2630 4680
rect 2670 4670 2680 4680
rect 2970 4670 2990 4680
rect 3100 4670 3110 4680
rect 3140 4670 3150 4680
rect 3480 4670 3500 4680
rect 5120 4670 5130 4680
rect 5140 4670 5150 4680
rect 5240 4670 5250 4680
rect 5390 4670 5480 4680
rect 5650 4670 5780 4680
rect 6330 4670 6430 4680
rect 6570 4670 6640 4680
rect 7690 4670 7700 4680
rect 7720 4670 7730 4680
rect 7760 4670 7770 4680
rect 7780 4670 7800 4680
rect 7830 4670 7840 4680
rect 7860 4670 7870 4680
rect 7970 4670 7980 4680
rect 8050 4670 8070 4680
rect 8500 4670 8510 4680
rect 8990 4670 9000 4680
rect 0 4660 90 4670
rect 100 4660 110 4670
rect 2620 4660 2640 4670
rect 3030 4660 3050 4670
rect 3100 4660 3110 4670
rect 3130 4660 3140 4670
rect 3260 4660 3270 4670
rect 3410 4660 3420 4670
rect 3490 4660 3500 4670
rect 5230 4660 5250 4670
rect 5390 4660 5490 4670
rect 5740 4660 5790 4670
rect 5940 4660 5990 4670
rect 6080 4660 6190 4670
rect 6230 4660 6250 4670
rect 6300 4660 6420 4670
rect 6580 4660 6640 4670
rect 7680 4660 7690 4670
rect 7720 4660 7730 4670
rect 7790 4660 7800 4670
rect 7830 4660 7840 4670
rect 8000 4660 8010 4670
rect 8870 4660 8880 4670
rect 8970 4660 8980 4670
rect 0 4650 90 4660
rect 2500 4650 2510 4660
rect 3010 4650 3050 4660
rect 3100 4650 3110 4660
rect 3130 4650 3150 4660
rect 3160 4650 3170 4660
rect 5140 4650 5150 4660
rect 5240 4650 5250 4660
rect 5390 4650 5500 4660
rect 5770 4650 6260 4660
rect 6300 4650 6420 4660
rect 6580 4650 6640 4660
rect 7380 4650 7390 4660
rect 7520 4650 7560 4660
rect 7660 4650 7670 4660
rect 7770 4650 7780 4660
rect 8540 4650 8550 4660
rect 8640 4650 8650 4660
rect 8790 4650 8800 4660
rect 30 4640 40 4650
rect 3010 4640 3030 4650
rect 3090 4640 3110 4650
rect 3130 4640 3150 4650
rect 3320 4640 3330 4650
rect 5150 4640 5170 4650
rect 5400 4640 5500 4650
rect 5830 4640 6080 4650
rect 6190 4640 6200 4650
rect 6230 4640 6410 4650
rect 6580 4640 6630 4650
rect 6650 4640 6660 4650
rect 7490 4640 7500 4650
rect 7820 4640 7830 4650
rect 8010 4640 8020 4650
rect 8090 4640 8100 4650
rect 8870 4640 8880 4650
rect 8940 4640 8950 4650
rect 8980 4640 8990 4650
rect 3010 4630 3020 4640
rect 3090 4630 3100 4640
rect 3340 4630 3360 4640
rect 5160 4630 5170 4640
rect 5200 4630 5210 4640
rect 5400 4630 5510 4640
rect 5860 4630 5870 4640
rect 5960 4630 6050 4640
rect 6240 4630 6410 4640
rect 6580 4630 6630 4640
rect 7600 4630 7610 4640
rect 7730 4630 7740 4640
rect 7810 4630 7820 4640
rect 7880 4630 7910 4640
rect 8020 4630 8030 4640
rect 8070 4630 8080 4640
rect 8310 4630 8320 4640
rect 8350 4630 8360 4640
rect 8550 4630 8560 4640
rect 8610 4630 8620 4640
rect 8840 4630 8850 4640
rect 8860 4630 8870 4640
rect 9250 4630 9260 4640
rect 2890 4620 2910 4630
rect 2970 4620 2980 4630
rect 3300 4620 3310 4630
rect 3340 4620 3350 4630
rect 3370 4620 3390 4630
rect 5170 4620 5180 4630
rect 5380 4620 5520 4630
rect 5970 4620 5980 4630
rect 5990 4620 6020 4630
rect 6570 4620 6620 4630
rect 7600 4620 7610 4630
rect 7730 4620 7740 4630
rect 7810 4620 7820 4630
rect 7870 4620 7880 4630
rect 8280 4620 8290 4630
rect 9750 4620 9760 4630
rect 2890 4610 2920 4620
rect 3000 4610 3010 4620
rect 3350 4610 3400 4620
rect 3450 4610 3460 4620
rect 5170 4610 5180 4620
rect 5380 4610 5520 4620
rect 5800 4610 5810 4620
rect 5890 4610 5900 4620
rect 6570 4610 6590 4620
rect 6600 4610 6610 4620
rect 7870 4610 7880 4620
rect 8810 4610 8820 4620
rect 8970 4610 8980 4620
rect 9740 4610 9750 4620
rect 3000 4600 3010 4610
rect 3280 4600 3290 4610
rect 3350 4600 3360 4610
rect 3370 4600 3390 4610
rect 5210 4600 5230 4610
rect 5390 4600 5530 4610
rect 5610 4600 5640 4610
rect 5790 4600 5800 4610
rect 5820 4600 6000 4610
rect 6560 4600 6580 4610
rect 7880 4600 7890 4610
rect 8210 4600 8220 4610
rect 8250 4600 8260 4610
rect 8330 4600 8340 4610
rect 8570 4600 8580 4610
rect 8830 4600 8840 4610
rect 8860 4600 8870 4610
rect 3220 4590 3230 4600
rect 3280 4590 3290 4600
rect 3350 4590 3360 4600
rect 3370 4590 3380 4600
rect 3440 4590 3450 4600
rect 3460 4590 3470 4600
rect 5220 4590 5230 4600
rect 5390 4590 5530 4600
rect 5600 4590 5650 4600
rect 5780 4590 5790 4600
rect 5830 4590 5870 4600
rect 5890 4590 5910 4600
rect 6010 4590 6030 4600
rect 6080 4590 6110 4600
rect 6560 4590 6580 4600
rect 7580 4590 7590 4600
rect 7610 4590 7620 4600
rect 7660 4590 7670 4600
rect 7780 4590 7800 4600
rect 7840 4590 7850 4600
rect 8170 4590 8180 4600
rect 8250 4590 8260 4600
rect 8620 4590 8630 4600
rect 3220 4580 3230 4590
rect 3340 4580 3370 4590
rect 3440 4580 3450 4590
rect 5230 4580 5240 4590
rect 5390 4580 5530 4590
rect 5600 4580 5650 4590
rect 5780 4580 5790 4590
rect 5840 4580 5860 4590
rect 6030 4580 6070 4590
rect 6080 4580 6100 4590
rect 6110 4580 6170 4590
rect 6550 4580 6580 4590
rect 7330 4580 7340 4590
rect 7380 4580 7390 4590
rect 7480 4580 7490 4590
rect 7740 4580 7750 4590
rect 7780 4580 7790 4590
rect 7800 4580 7810 4590
rect 8580 4580 8590 4590
rect 8660 4580 8670 4590
rect 8960 4580 8970 4590
rect 3200 4570 3220 4580
rect 3260 4570 3270 4580
rect 3340 4570 3360 4580
rect 5230 4570 5240 4580
rect 5290 4570 5300 4580
rect 5410 4570 5430 4580
rect 5450 4570 5530 4580
rect 5600 4570 5610 4580
rect 5630 4570 5660 4580
rect 5780 4570 5790 4580
rect 6130 4570 6210 4580
rect 6530 4570 6570 4580
rect 7650 4570 7660 4580
rect 7700 4570 7710 4580
rect 7740 4570 7750 4580
rect 8090 4570 8100 4580
rect 8120 4570 8130 4580
rect 8150 4570 8160 4580
rect 8220 4570 8230 4580
rect 8280 4570 8290 4580
rect 8320 4570 8330 4580
rect 8340 4570 8350 4580
rect 8660 4570 8670 4580
rect 3130 4560 3140 4570
rect 3170 4560 3180 4570
rect 3200 4560 3220 4570
rect 3330 4560 3350 4570
rect 3380 4560 3390 4570
rect 3440 4560 3450 4570
rect 5230 4560 5240 4570
rect 5290 4560 5300 4570
rect 5410 4560 5430 4570
rect 5460 4560 5540 4570
rect 5600 4560 5610 4570
rect 5640 4560 5650 4570
rect 5660 4560 5670 4570
rect 5780 4560 5800 4570
rect 6140 4560 6210 4570
rect 6240 4560 6280 4570
rect 6520 4560 6560 4570
rect 7370 4560 7380 4570
rect 7650 4560 7670 4570
rect 7750 4560 7760 4570
rect 8090 4560 8100 4570
rect 8130 4560 8140 4570
rect 8190 4560 8200 4570
rect 8660 4560 8670 4570
rect 2810 4550 2820 4560
rect 3040 4550 3050 4560
rect 3140 4550 3150 4560
rect 3170 4550 3190 4560
rect 3200 4550 3210 4560
rect 3330 4550 3340 4560
rect 5240 4550 5250 4560
rect 5470 4550 5540 4560
rect 5580 4550 5610 4560
rect 5790 4550 5800 4560
rect 6130 4550 6210 4560
rect 6230 4550 6240 4560
rect 6270 4550 6280 4560
rect 6520 4550 6550 4560
rect 7330 4550 7360 4560
rect 7380 4550 7390 4560
rect 7540 4550 7550 4560
rect 8010 4550 8020 4560
rect 8030 4550 8040 4560
rect 8080 4550 8100 4560
rect 8130 4550 8140 4560
rect 8640 4550 8650 4560
rect 2810 4540 2820 4550
rect 3040 4540 3050 4550
rect 3180 4540 3200 4550
rect 3250 4540 3260 4550
rect 5300 4540 5310 4550
rect 5460 4540 5540 4550
rect 5580 4540 5610 4550
rect 5670 4540 5680 4550
rect 6140 4540 6160 4550
rect 6200 4540 6210 4550
rect 6220 4540 6230 4550
rect 6270 4540 6280 4550
rect 6520 4540 6550 4550
rect 7380 4540 7390 4550
rect 8040 4540 8050 4550
rect 8090 4540 8100 4550
rect 8200 4540 8220 4550
rect 8540 4540 8550 4550
rect 9680 4540 9690 4550
rect 9990 4540 9990 4550
rect 2980 4530 2990 4540
rect 3240 4530 3250 4540
rect 5250 4530 5260 4540
rect 5300 4530 5320 4540
rect 5400 4530 5410 4540
rect 5450 4530 5540 4540
rect 5580 4530 5620 4540
rect 6140 4530 6150 4540
rect 6200 4530 6230 4540
rect 6260 4530 6270 4540
rect 6280 4530 6290 4540
rect 6510 4530 6540 4540
rect 7340 4530 7360 4540
rect 7490 4530 7500 4540
rect 7530 4530 7540 4540
rect 7620 4530 7630 4540
rect 7680 4530 7690 4540
rect 8050 4530 8060 4540
rect 9990 4530 9990 4540
rect 3010 4520 3020 4530
rect 3210 4520 3220 4530
rect 3240 4520 3250 4530
rect 3420 4520 3430 4530
rect 5260 4520 5270 4530
rect 5300 4520 5320 4530
rect 5460 4520 5540 4530
rect 5580 4520 5620 4530
rect 6260 4520 6270 4530
rect 6510 4520 6540 4530
rect 7330 4520 7350 4530
rect 7900 4520 7910 4530
rect 7980 4520 7990 4530
rect 8050 4520 8060 4530
rect 8160 4520 8170 4530
rect 8330 4520 8340 4530
rect 9980 4520 9990 4530
rect 3020 4510 3030 4520
rect 3040 4510 3050 4520
rect 3220 4510 3240 4520
rect 3410 4510 3420 4520
rect 5300 4510 5340 4520
rect 5460 4510 5540 4520
rect 5580 4510 5610 4520
rect 5690 4510 5700 4520
rect 5810 4510 5820 4520
rect 5860 4510 5870 4520
rect 6250 4510 6260 4520
rect 6510 4510 6530 4520
rect 7990 4510 8000 4520
rect 8010 4510 8020 4520
rect 8160 4510 8170 4520
rect 8230 4510 8240 4520
rect 8340 4510 8350 4520
rect 9220 4510 9230 4520
rect 9970 4510 9990 4520
rect 3240 4500 3250 4510
rect 5270 4500 5280 4510
rect 5310 4500 5350 4510
rect 5470 4500 5540 4510
rect 5570 4500 5610 4510
rect 5700 4500 5710 4510
rect 5810 4500 5840 4510
rect 5860 4500 5870 4510
rect 6250 4500 6260 4510
rect 6510 4500 6530 4510
rect 7330 4500 7340 4510
rect 7530 4500 7540 4510
rect 7800 4500 7810 4510
rect 7990 4500 8000 4510
rect 8010 4500 8020 4510
rect 8140 4500 8150 4510
rect 8340 4500 8350 4510
rect 8400 4500 8410 4510
rect 8930 4500 8940 4510
rect 9960 4500 9980 4510
rect 3400 4490 3410 4500
rect 3910 4490 3930 4500
rect 5310 4490 5360 4500
rect 5390 4490 5420 4500
rect 5480 4490 5540 4500
rect 5570 4490 5600 4500
rect 5710 4490 5720 4500
rect 5800 4490 5820 4500
rect 5830 4490 5840 4500
rect 5850 4490 5870 4500
rect 6240 4490 6250 4500
rect 6510 4490 6530 4500
rect 7350 4490 7360 4500
rect 7410 4490 7420 4500
rect 7510 4490 7520 4500
rect 7880 4490 7890 4500
rect 7950 4490 7960 4500
rect 8140 4490 8150 4500
rect 9950 4490 9980 4500
rect 3070 4480 3080 4490
rect 3090 4480 3100 4490
rect 3910 4480 3930 4490
rect 5280 4480 5290 4490
rect 5310 4480 5360 4490
rect 5400 4480 5420 4490
rect 5490 4480 5590 4490
rect 5720 4480 5730 4490
rect 5800 4480 5810 4490
rect 5840 4480 5860 4490
rect 6190 4480 6210 4490
rect 6230 4480 6240 4490
rect 6410 4480 6420 4490
rect 6510 4480 6530 4490
rect 7340 4480 7360 4490
rect 7950 4480 7960 4490
rect 8020 4480 8030 4490
rect 8140 4480 8150 4490
rect 8170 4480 8180 4490
rect 8240 4480 8250 4490
rect 8270 4480 8280 4490
rect 8920 4480 8930 4490
rect 9940 4480 9970 4490
rect 3270 4470 3280 4480
rect 3890 4470 3950 4480
rect 5280 4470 5300 4480
rect 5330 4470 5350 4480
rect 5400 4470 5430 4480
rect 5500 4470 5590 4480
rect 5730 4470 5740 4480
rect 5790 4470 5800 4480
rect 5840 4470 5860 4480
rect 5890 4470 5920 4480
rect 6180 4470 6190 4480
rect 6200 4470 6210 4480
rect 6220 4470 6230 4480
rect 6400 4470 6430 4480
rect 6510 4470 6530 4480
rect 7350 4470 7360 4480
rect 7830 4470 7840 4480
rect 7880 4470 7890 4480
rect 7920 4470 7930 4480
rect 8000 4470 8010 4480
rect 8140 4470 8150 4480
rect 8170 4470 8180 4480
rect 8280 4470 8290 4480
rect 8330 4470 8340 4480
rect 9930 4470 9960 4480
rect 3030 4460 3040 4470
rect 3110 4460 3120 4470
rect 3160 4460 3170 4470
rect 3280 4460 3290 4470
rect 3940 4460 3950 4470
rect 5280 4460 5290 4470
rect 5320 4460 5350 4470
rect 5410 4460 5430 4470
rect 5500 4460 5590 4470
rect 5740 4460 5750 4470
rect 5830 4460 5850 4470
rect 5890 4460 5920 4470
rect 6390 4460 6430 4470
rect 6500 4460 6520 4470
rect 7830 4460 7840 4470
rect 7880 4460 7890 4470
rect 7920 4460 7930 4470
rect 8000 4460 8010 4470
rect 8030 4460 8040 4470
rect 8140 4460 8150 4470
rect 9920 4460 9950 4470
rect 3110 4450 3120 4460
rect 3160 4450 3170 4460
rect 5300 4450 5310 4460
rect 5330 4450 5360 4460
rect 5420 4450 5430 4460
rect 5500 4450 5600 4460
rect 5750 4450 5760 4460
rect 5830 4450 5850 4460
rect 5890 4450 5930 4460
rect 6140 4450 6180 4460
rect 6380 4450 6430 4460
rect 6500 4450 6530 4460
rect 7410 4450 7420 4460
rect 7960 4450 7970 4460
rect 8090 4450 8100 4460
rect 8140 4450 8150 4460
rect 9910 4450 9940 4460
rect 3100 4440 3110 4450
rect 3250 4440 3260 4450
rect 3280 4440 3290 4450
rect 5290 4440 5300 4450
rect 5340 4440 5370 4450
rect 5420 4440 5430 4450
rect 5500 4440 5600 4450
rect 5760 4440 5770 4450
rect 5780 4440 5790 4450
rect 5820 4440 5850 4450
rect 5900 4440 5920 4450
rect 5940 4440 5980 4450
rect 6010 4440 6030 4450
rect 6120 4440 6140 4450
rect 6170 4440 6200 4450
rect 6370 4440 6430 4450
rect 6500 4440 6520 4450
rect 7410 4440 7420 4450
rect 7960 4440 7970 4450
rect 8090 4440 8100 4450
rect 8220 4440 8230 4450
rect 8900 4440 8910 4450
rect 9890 4440 9930 4450
rect 2990 4430 3020 4440
rect 3140 4430 3150 4440
rect 3170 4430 3180 4440
rect 3250 4430 3260 4440
rect 3270 4430 3280 4440
rect 3300 4430 3310 4440
rect 3910 4430 3940 4440
rect 5300 4430 5320 4440
rect 5340 4430 5370 4440
rect 5410 4430 5430 4440
rect 5510 4430 5600 4440
rect 5780 4430 5800 4440
rect 5820 4430 5840 4440
rect 5940 4430 6090 4440
rect 6100 4430 6180 4440
rect 6190 4430 6200 4440
rect 6360 4430 6440 4440
rect 6490 4430 6530 4440
rect 7410 4430 7420 4440
rect 8080 4430 8090 4440
rect 8100 4430 8110 4440
rect 8140 4430 8150 4440
rect 9880 4430 9920 4440
rect 3100 4420 3130 4430
rect 3150 4420 3160 4430
rect 3250 4420 3260 4430
rect 3280 4420 3290 4430
rect 3920 4420 3940 4430
rect 5310 4420 5320 4430
rect 5350 4420 5380 4430
rect 5410 4420 5440 4430
rect 5510 4420 5600 4430
rect 5790 4420 5840 4430
rect 5960 4420 5970 4430
rect 6010 4420 6090 4430
rect 6100 4420 6170 4430
rect 6340 4420 6350 4430
rect 6360 4420 6440 4430
rect 6490 4420 6520 4430
rect 7350 4420 7370 4430
rect 7800 4420 7810 4430
rect 7840 4420 7850 4430
rect 7890 4420 7900 4430
rect 7930 4420 7940 4430
rect 8130 4420 8140 4430
rect 9200 4420 9210 4430
rect 9860 4420 9900 4430
rect 2750 4410 2760 4420
rect 2970 4410 2980 4420
rect 2990 4410 3000 4420
rect 3010 4410 3020 4420
rect 3050 4410 3060 4420
rect 3110 4410 3130 4420
rect 3180 4410 3190 4420
rect 3290 4410 3300 4420
rect 3310 4410 3320 4420
rect 3920 4410 3940 4420
rect 4620 4410 4660 4420
rect 5320 4410 5330 4420
rect 5350 4410 5380 4420
rect 5410 4410 5450 4420
rect 5520 4410 5590 4420
rect 5810 4410 5860 4420
rect 6010 4410 6060 4420
rect 6070 4410 6110 4420
rect 6130 4410 6210 4420
rect 6330 4410 6440 4420
rect 6490 4410 6520 4420
rect 7840 4410 7850 4420
rect 7940 4410 7960 4420
rect 8050 4410 8060 4420
rect 9850 4410 9890 4420
rect 2660 4400 2670 4410
rect 2960 4400 2970 4410
rect 3050 4400 3060 4410
rect 3110 4400 3130 4410
rect 3180 4400 3190 4410
rect 4610 4400 4700 4410
rect 5310 4400 5330 4410
rect 5360 4400 5390 4410
rect 5400 4400 5460 4410
rect 5520 4400 5570 4410
rect 5840 4400 5910 4410
rect 5950 4400 5970 4410
rect 6020 4400 6050 4410
rect 6070 4400 6100 4410
rect 6140 4400 6200 4410
rect 6300 4400 6440 4410
rect 6480 4400 6520 4410
rect 7420 4400 7430 4410
rect 9540 4400 9550 4410
rect 9860 4400 9870 4410
rect 2830 4390 2840 4400
rect 2960 4390 2970 4400
rect 3050 4390 3070 4400
rect 3180 4390 3200 4400
rect 3260 4390 3270 4400
rect 3280 4390 3300 4400
rect 4610 4390 4650 4400
rect 4680 4390 4710 4400
rect 5370 4390 5390 4400
rect 5440 4390 5460 4400
rect 5520 4390 5570 4400
rect 5860 4390 5970 4400
rect 6010 4390 6040 4400
rect 6080 4390 6110 4400
rect 6130 4390 6200 4400
rect 6290 4390 6450 4400
rect 6470 4390 6510 4400
rect 7990 4390 8000 4400
rect 8680 4390 8710 4400
rect 9860 4390 9870 4400
rect 2640 4380 2650 4390
rect 2800 4380 2820 4390
rect 2860 4380 2870 4390
rect 3050 4380 3060 4390
rect 3070 4380 3080 4390
rect 3190 4380 3210 4390
rect 3230 4380 3240 4390
rect 3280 4380 3300 4390
rect 3320 4380 3330 4390
rect 4600 4380 4630 4390
rect 4700 4380 4730 4390
rect 5320 4380 5330 4390
rect 5370 4380 5400 4390
rect 5420 4380 5460 4390
rect 5520 4380 5570 4390
rect 5890 4380 5950 4390
rect 5960 4380 5980 4390
rect 6000 4380 6050 4390
rect 6070 4380 6080 4390
rect 6100 4380 6150 4390
rect 6160 4380 6190 4390
rect 6280 4380 6500 4390
rect 7850 4380 7860 4390
rect 7920 4380 7930 4390
rect 8660 4380 8670 4390
rect 9860 4380 9870 4390
rect 2640 4370 2650 4380
rect 2700 4370 2710 4380
rect 2850 4370 2860 4380
rect 2970 4370 2980 4380
rect 3040 4370 3060 4380
rect 3080 4370 3090 4380
rect 3200 4370 3240 4380
rect 3260 4370 3270 4380
rect 3280 4370 3300 4380
rect 4590 4370 4610 4380
rect 4720 4370 4740 4380
rect 4840 4370 4850 4380
rect 5380 4370 5410 4380
rect 5430 4370 5470 4380
rect 5520 4370 5560 4380
rect 5930 4370 5960 4380
rect 5980 4370 5990 4380
rect 6050 4370 6070 4380
rect 6260 4370 6500 4380
rect 7330 4370 7340 4380
rect 7420 4370 7430 4380
rect 7810 4370 7820 4380
rect 7850 4370 7860 4380
rect 8650 4370 8660 4380
rect 9850 4370 9870 4380
rect 2830 4360 2840 4370
rect 2950 4360 2960 4370
rect 2970 4360 2980 4370
rect 3040 4360 3060 4370
rect 3070 4360 3080 4370
rect 3230 4360 3240 4370
rect 3260 4360 3270 4370
rect 3290 4360 3300 4370
rect 4580 4360 4610 4370
rect 4750 4360 4820 4370
rect 5380 4360 5410 4370
rect 5420 4360 5470 4370
rect 5540 4360 5560 4370
rect 5950 4360 5980 4370
rect 6240 4360 6500 4370
rect 7360 4360 7370 4370
rect 7420 4360 7430 4370
rect 7850 4360 7860 4370
rect 8550 4360 8560 4370
rect 8670 4360 8680 4370
rect 9490 4360 9500 4370
rect 9850 4360 9860 4370
rect 2820 4350 2830 4360
rect 2940 4350 2960 4360
rect 2970 4350 2980 4360
rect 3060 4350 3070 4360
rect 3250 4350 3280 4360
rect 3300 4350 3310 4360
rect 3340 4350 3350 4360
rect 4310 4350 4320 4360
rect 4580 4350 4600 4360
rect 4780 4350 4800 4360
rect 4810 4350 4840 4360
rect 4860 4350 4890 4360
rect 5390 4350 5470 4360
rect 6000 4350 6080 4360
rect 6150 4350 6490 4360
rect 7350 4350 7360 4360
rect 7420 4350 7430 4360
rect 7820 4350 7830 4360
rect 8590 4350 8600 4360
rect 8670 4350 8680 4360
rect 9180 4350 9190 4360
rect 9480 4350 9490 4360
rect 9840 4350 9850 4360
rect 2830 4340 2840 4350
rect 2950 4340 2970 4350
rect 2980 4340 2990 4350
rect 3040 4340 3050 4350
rect 3270 4340 3280 4350
rect 4310 4340 4320 4350
rect 4570 4340 4590 4350
rect 4830 4340 4890 4350
rect 5340 4340 5350 4350
rect 5400 4340 5430 4350
rect 5450 4340 5470 4350
rect 6060 4340 6480 4350
rect 7350 4340 7380 4350
rect 7420 4340 7430 4350
rect 8540 4340 8550 4350
rect 8650 4340 8660 4350
rect 8720 4340 8730 4350
rect 8860 4340 8870 4350
rect 9470 4340 9480 4350
rect 9830 4340 9840 4350
rect 9900 4340 9910 4350
rect 9960 4340 9980 4350
rect 2840 4330 2850 4340
rect 2950 4330 2960 4340
rect 3270 4330 3280 4340
rect 4570 4330 4590 4340
rect 4840 4330 4900 4340
rect 5410 4330 5480 4340
rect 6190 4330 6200 4340
rect 6220 4330 6480 4340
rect 7360 4330 7370 4340
rect 8450 4330 8460 4340
rect 8730 4330 8740 4340
rect 9180 4330 9190 4340
rect 9460 4330 9470 4340
rect 9820 4330 9840 4340
rect 9880 4330 9890 4340
rect 3010 4320 3020 4330
rect 3140 4320 3160 4330
rect 3170 4320 3190 4330
rect 3260 4320 3270 4330
rect 4230 4320 4240 4330
rect 4320 4320 4330 4330
rect 4560 4320 4590 4330
rect 4860 4320 4910 4330
rect 5410 4320 5490 4330
rect 6180 4320 6470 4330
rect 6580 4320 6590 4330
rect 8510 4320 8520 4330
rect 8710 4320 8720 4330
rect 9180 4320 9190 4330
rect 9450 4320 9460 4330
rect 9880 4320 9900 4330
rect 9920 4320 9940 4330
rect 2810 4310 2820 4320
rect 2840 4310 2850 4320
rect 3000 4310 3010 4320
rect 3140 4310 3160 4320
rect 3180 4310 3200 4320
rect 3230 4310 3250 4320
rect 4220 4310 4250 4320
rect 4550 4310 4580 4320
rect 4880 4310 4910 4320
rect 5420 4310 5500 4320
rect 5940 4310 5950 4320
rect 5970 4310 5980 4320
rect 5990 4310 6010 4320
rect 6140 4310 6460 4320
rect 6570 4310 6590 4320
rect 7290 4310 7310 4320
rect 7320 4310 7330 4320
rect 8470 4310 8480 4320
rect 8600 4310 8610 4320
rect 8670 4310 8680 4320
rect 8860 4310 8870 4320
rect 9180 4310 9190 4320
rect 9880 4310 9890 4320
rect 9910 4310 9920 4320
rect 9950 4310 9970 4320
rect 2560 4300 2570 4310
rect 2810 4300 2820 4310
rect 2910 4300 2930 4310
rect 2940 4300 2950 4310
rect 2960 4300 3000 4310
rect 3130 4300 3160 4310
rect 3170 4300 3180 4310
rect 3190 4300 3200 4310
rect 3210 4300 3220 4310
rect 3240 4300 3250 4310
rect 3290 4300 3300 4310
rect 4200 4300 4270 4310
rect 4550 4300 4570 4310
rect 4890 4300 4920 4310
rect 5420 4300 5500 4310
rect 5920 4300 6450 4310
rect 6550 4300 6580 4310
rect 8480 4300 8500 4310
rect 8600 4300 8610 4310
rect 8660 4300 8670 4310
rect 8690 4300 8710 4310
rect 9940 4300 9950 4310
rect 9960 4300 9970 4310
rect 2840 4290 2850 4300
rect 2910 4290 2920 4300
rect 2940 4290 2950 4300
rect 2970 4290 2990 4300
rect 3050 4290 3060 4300
rect 3140 4290 3150 4300
rect 3160 4290 3170 4300
rect 3180 4290 3200 4300
rect 3290 4290 3300 4300
rect 4180 4290 4290 4300
rect 4550 4290 4570 4300
rect 4890 4290 4920 4300
rect 5430 4290 5510 4300
rect 5930 4290 6090 4300
rect 6100 4290 6150 4300
rect 6170 4290 6450 4300
rect 6550 4290 6580 4300
rect 7220 4290 7230 4300
rect 8490 4290 8500 4300
rect 9920 4290 9930 4300
rect 2880 4280 2900 4290
rect 2940 4280 2960 4290
rect 2980 4280 2990 4290
rect 3040 4280 3060 4290
rect 3080 4280 3090 4290
rect 3140 4280 3150 4290
rect 3170 4280 3190 4290
rect 3280 4280 3290 4290
rect 4180 4280 4300 4290
rect 4540 4280 4570 4290
rect 4910 4280 4940 4290
rect 5440 4280 5510 4290
rect 5940 4280 6080 4290
rect 6180 4280 6440 4290
rect 6540 4280 6570 4290
rect 7180 4280 7200 4290
rect 8440 4280 8450 4290
rect 8520 4280 8530 4290
rect 8580 4280 8590 4290
rect 9420 4280 9430 4290
rect 9770 4280 9790 4290
rect 9870 4280 9880 4290
rect 9920 4280 9930 4290
rect 9940 4280 9950 4290
rect 2880 4270 2890 4280
rect 2920 4270 2960 4280
rect 2970 4270 2980 4280
rect 3030 4270 3040 4280
rect 3090 4270 3110 4280
rect 3140 4270 3160 4280
rect 3180 4270 3190 4280
rect 3280 4270 3290 4280
rect 4170 4270 4210 4280
rect 4230 4270 4310 4280
rect 4540 4270 4560 4280
rect 4910 4270 4950 4280
rect 5440 4270 5510 4280
rect 5950 4270 6430 4280
rect 6540 4270 6570 4280
rect 7150 4270 7160 4280
rect 8440 4270 8450 4280
rect 8470 4270 8480 4280
rect 9410 4270 9420 4280
rect 9760 4270 9810 4280
rect 9820 4270 9830 4280
rect 9860 4270 9880 4280
rect 9910 4270 9920 4280
rect 9930 4270 9940 4280
rect 2830 4260 2850 4270
rect 2890 4260 2930 4270
rect 2940 4260 2950 4270
rect 2960 4260 2980 4270
rect 3030 4260 3040 4270
rect 3050 4260 3060 4270
rect 3090 4260 3100 4270
rect 3160 4260 3170 4270
rect 3180 4260 3190 4270
rect 3200 4260 3210 4270
rect 3230 4260 3240 4270
rect 4160 4260 4200 4270
rect 4290 4260 4320 4270
rect 4520 4260 4560 4270
rect 4910 4260 4960 4270
rect 5360 4260 5370 4270
rect 5450 4260 5460 4270
rect 5470 4260 5520 4270
rect 5950 4260 6380 4270
rect 6400 4260 6420 4270
rect 6530 4260 6560 4270
rect 7090 4260 7170 4270
rect 7420 4260 7440 4270
rect 8480 4260 8490 4270
rect 8590 4260 8610 4270
rect 9400 4260 9410 4270
rect 9760 4260 9780 4270
rect 9900 4260 9910 4270
rect 2810 4250 2830 4260
rect 2890 4250 2930 4260
rect 2950 4250 2970 4260
rect 3030 4250 3080 4260
rect 3130 4250 3140 4260
rect 3160 4250 3170 4260
rect 3200 4250 3210 4260
rect 3230 4250 3240 4260
rect 4160 4250 4200 4260
rect 4300 4250 4330 4260
rect 4520 4250 4550 4260
rect 4910 4250 4970 4260
rect 5370 4250 5380 4260
rect 5460 4250 5470 4260
rect 5480 4250 5520 4260
rect 5980 4250 6370 4260
rect 6520 4250 6560 4260
rect 7050 4250 7080 4260
rect 7150 4250 7160 4260
rect 7170 4250 7190 4260
rect 7370 4250 7390 4260
rect 7410 4250 7440 4260
rect 8490 4250 8500 4260
rect 8840 4250 8850 4260
rect 9750 4250 9770 4260
rect 9850 4250 9860 4260
rect 9870 4250 9880 4260
rect 2820 4240 2830 4250
rect 2870 4240 2890 4250
rect 2910 4240 2920 4250
rect 2930 4240 2960 4250
rect 3070 4240 3140 4250
rect 3170 4240 3180 4250
rect 3200 4240 3210 4250
rect 3220 4240 3230 4250
rect 3240 4240 3250 4250
rect 4160 4240 4190 4250
rect 4330 4240 4340 4250
rect 4500 4240 4530 4250
rect 4910 4240 4980 4250
rect 5470 4240 5480 4250
rect 5490 4240 5530 4250
rect 5990 4240 6300 4250
rect 6310 4240 6370 4250
rect 6520 4240 6560 4250
rect 7080 4240 7090 4250
rect 7110 4240 7150 4250
rect 7170 4240 7180 4250
rect 7290 4240 7360 4250
rect 7370 4240 7410 4250
rect 9740 4240 9760 4250
rect 9820 4240 9850 4250
rect 9870 4240 9880 4250
rect 9990 4240 9990 4250
rect 2690 4230 2700 4240
rect 2880 4230 2890 4240
rect 2900 4230 2960 4240
rect 2970 4230 2980 4240
rect 3070 4230 3090 4240
rect 3130 4230 3140 4240
rect 3240 4230 3260 4240
rect 4140 4230 4170 4240
rect 4330 4230 4350 4240
rect 4490 4230 4530 4240
rect 4910 4230 4990 4240
rect 5480 4230 5540 4240
rect 5990 4230 6070 4240
rect 6080 4230 6270 4240
rect 6330 4230 6360 4240
rect 6520 4230 6570 4240
rect 7120 4230 7150 4240
rect 7260 4230 7270 4240
rect 7330 4230 7370 4240
rect 7380 4230 7390 4240
rect 7420 4230 7450 4240
rect 8460 4230 8470 4240
rect 9730 4230 9750 4240
rect 9820 4230 9830 4240
rect 9970 4230 9990 4240
rect 2890 4220 2910 4230
rect 2920 4220 2950 4230
rect 3040 4220 3080 4230
rect 3090 4220 3100 4230
rect 3180 4220 3190 4230
rect 3210 4220 3220 4230
rect 3240 4220 3260 4230
rect 4130 4220 4170 4230
rect 4330 4220 4360 4230
rect 4490 4220 4520 4230
rect 4920 4220 4990 4230
rect 5500 4220 5550 4230
rect 6110 4220 6260 4230
rect 6510 4220 6580 4230
rect 7120 4220 7130 4230
rect 7220 4220 7240 4230
rect 7300 4220 7390 4230
rect 7450 4220 7460 4230
rect 9360 4220 9370 4230
rect 9720 4220 9740 4230
rect 9860 4220 9870 4230
rect 9940 4220 9950 4230
rect 9980 4220 9990 4230
rect 2770 4210 2800 4220
rect 3030 4210 3040 4220
rect 3100 4210 3120 4220
rect 4130 4210 4160 4220
rect 4330 4210 4360 4220
rect 4470 4210 4510 4220
rect 4950 4210 5000 4220
rect 5490 4210 5500 4220
rect 5530 4210 5550 4220
rect 6120 4210 6250 4220
rect 6320 4210 6330 4220
rect 6500 4210 6580 4220
rect 7170 4210 7180 4220
rect 7280 4210 7300 4220
rect 7340 4210 7350 4220
rect 9710 4210 9730 4220
rect 9740 4210 9750 4220
rect 9810 4210 9830 4220
rect 9880 4210 9890 4220
rect 9930 4210 9950 4220
rect 9960 4210 9970 4220
rect 2790 4200 2800 4210
rect 3030 4200 3100 4210
rect 3170 4200 3180 4210
rect 3200 4200 3210 4210
rect 3230 4200 3240 4210
rect 4120 4200 4150 4210
rect 4350 4200 4360 4210
rect 4450 4200 4480 4210
rect 4970 4200 5000 4210
rect 5490 4200 5500 4210
rect 5540 4200 5560 4210
rect 6150 4200 6160 4210
rect 6180 4200 6210 4210
rect 6240 4200 6250 4210
rect 6270 4200 6290 4210
rect 6490 4200 6580 4210
rect 9710 4200 9720 4210
rect 9750 4200 9760 4210
rect 9810 4200 9820 4210
rect 9880 4200 9900 4210
rect 3170 4190 3180 4200
rect 4120 4190 4150 4200
rect 4370 4190 4380 4200
rect 4450 4190 4480 4200
rect 4980 4190 5010 4200
rect 5390 4190 5420 4200
rect 5550 4190 5570 4200
rect 6180 4190 6190 4200
rect 6280 4190 6290 4200
rect 6480 4190 6560 4200
rect 7260 4190 7270 4200
rect 9310 4190 9320 4200
rect 9690 4190 9720 4200
rect 9780 4190 9790 4200
rect 9870 4190 9880 4200
rect 2590 4180 2600 4190
rect 2860 4180 2890 4190
rect 3020 4180 3080 4190
rect 3090 4180 3110 4190
rect 3140 4180 3150 4190
rect 3220 4180 3230 4190
rect 4110 4180 4140 4190
rect 4370 4180 4410 4190
rect 4450 4180 4460 4190
rect 4680 4180 4690 4190
rect 4990 4180 5020 4190
rect 5560 4180 5570 4190
rect 6260 4180 6280 4190
rect 6290 4180 6300 4190
rect 6480 4180 6580 4190
rect 8820 4180 8830 4190
rect 9280 4180 9290 4190
rect 9310 4180 9320 4190
rect 9690 4180 9710 4190
rect 9800 4180 9810 4190
rect 9840 4180 9850 4190
rect 9880 4180 9900 4190
rect 2590 4170 2600 4180
rect 2840 4170 2870 4180
rect 2900 4170 2940 4180
rect 3020 4170 3110 4180
rect 3130 4170 3170 4180
rect 3200 4170 3220 4180
rect 4100 4170 4120 4180
rect 4380 4170 4410 4180
rect 4440 4170 4460 4180
rect 4670 4170 4710 4180
rect 5000 4170 5020 4180
rect 5390 4170 5400 4180
rect 5570 4170 5590 4180
rect 6170 4170 6180 4180
rect 6470 4170 6580 4180
rect 7260 4170 7270 4180
rect 9310 4170 9320 4180
rect 9810 4170 9820 4180
rect 2840 4160 2850 4170
rect 2860 4160 2870 4170
rect 2890 4160 2950 4170
rect 3010 4160 3110 4170
rect 3120 4160 3130 4170
rect 3190 4160 3210 4170
rect 4100 4160 4110 4170
rect 4400 4160 4420 4170
rect 4640 4160 4710 4170
rect 5010 4160 5030 4170
rect 5410 4160 5420 4170
rect 5490 4160 5500 4170
rect 5580 4160 5600 4170
rect 6460 4160 6540 4170
rect 6560 4160 6580 4170
rect 7340 4160 7350 4170
rect 7470 4160 7480 4170
rect 9310 4160 9320 4170
rect 9820 4160 9830 4170
rect 2860 4150 2880 4160
rect 2900 4150 2920 4160
rect 2930 4150 2970 4160
rect 3010 4150 3090 4160
rect 4100 4150 4110 4160
rect 4610 4150 4720 4160
rect 5010 4150 5030 4160
rect 5430 4150 5440 4160
rect 5590 4150 5610 4160
rect 6440 4150 6540 4160
rect 6560 4150 6580 4160
rect 7470 4150 7480 4160
rect 9820 4150 9850 4160
rect 2870 4140 2880 4150
rect 2900 4140 2920 4150
rect 2930 4140 2970 4150
rect 3040 4140 3090 4150
rect 3150 4140 3190 4150
rect 3260 4140 3270 4150
rect 4090 4140 4100 4150
rect 4590 4140 4720 4150
rect 4770 4140 4900 4150
rect 5010 4140 5040 4150
rect 5440 4140 5450 4150
rect 5490 4140 5500 4150
rect 5600 4140 5620 4150
rect 6430 4140 6520 4150
rect 7380 4140 7390 4150
rect 7470 4140 7480 4150
rect 9660 4140 9670 4150
rect 9810 4140 9820 4150
rect 9860 4140 9870 4150
rect 9950 4140 9990 4150
rect 2900 4130 2910 4140
rect 2950 4130 2990 4140
rect 3020 4130 3040 4140
rect 3120 4130 3130 4140
rect 3140 4130 3170 4140
rect 3190 4130 3210 4140
rect 4080 4130 4090 4140
rect 4580 4130 4760 4140
rect 4920 4130 4950 4140
rect 4980 4130 5040 4140
rect 5440 4130 5450 4140
rect 5490 4130 5500 4140
rect 5610 4130 5630 4140
rect 6420 4130 6520 4140
rect 7240 4130 7250 4140
rect 7420 4130 7430 4140
rect 7450 4130 7460 4140
rect 9650 4130 9660 4140
rect 9860 4130 9880 4140
rect 9950 4130 9990 4140
rect 2870 4120 2880 4130
rect 2970 4120 2990 4130
rect 3020 4120 3030 4130
rect 3040 4120 3070 4130
rect 3160 4120 3200 4130
rect 3240 4120 3250 4130
rect 4080 4120 4090 4130
rect 4560 4120 4730 4130
rect 4950 4120 5030 4130
rect 5440 4120 5450 4130
rect 5620 4120 5640 4130
rect 6410 4120 6480 4130
rect 6500 4120 6520 4130
rect 7440 4120 7460 4130
rect 9820 4120 9840 4130
rect 9870 4120 9890 4130
rect 9960 4120 9970 4130
rect 2840 4110 2860 4120
rect 2870 4110 2890 4120
rect 2970 4110 3000 4120
rect 3020 4110 3080 4120
rect 3130 4110 3140 4120
rect 3170 4110 3180 4120
rect 3210 4110 3220 4120
rect 4080 4110 4090 4120
rect 4550 4110 4710 4120
rect 5030 4110 5080 4120
rect 5450 4110 5460 4120
rect 5630 4110 5650 4120
rect 6400 4110 6470 4120
rect 6500 4110 6520 4120
rect 7450 4110 7470 4120
rect 9820 4110 9910 4120
rect 9970 4110 9980 4120
rect 2830 4100 2840 4110
rect 2860 4100 2870 4110
rect 2960 4100 3010 4110
rect 3090 4100 3170 4110
rect 4070 4100 4080 4110
rect 4550 4100 4670 4110
rect 5010 4100 5030 4110
rect 5050 4100 5080 4110
rect 5450 4100 5460 4110
rect 5640 4100 5660 4110
rect 6390 4100 6460 4110
rect 6500 4100 6510 4110
rect 7230 4100 7240 4110
rect 7470 4100 7480 4110
rect 9790 4100 9920 4110
rect 2820 4090 2840 4100
rect 2950 4090 2960 4100
rect 2970 4090 3010 4100
rect 3270 4090 3280 4100
rect 4070 4090 4080 4100
rect 4540 4090 4670 4100
rect 4900 4090 4920 4100
rect 5060 4090 5090 4100
rect 5430 4090 5460 4100
rect 5660 4090 5680 4100
rect 6370 4090 6440 4100
rect 6500 4090 6510 4100
rect 7480 4090 7490 4100
rect 7500 4090 7510 4100
rect 9620 4090 9630 4100
rect 9870 4090 9900 4100
rect 9920 4090 9940 4100
rect 2830 4080 2850 4090
rect 2970 4080 2990 4090
rect 3070 4080 3080 4090
rect 3130 4080 3170 4090
rect 3270 4080 3280 4090
rect 4060 4080 4070 4090
rect 4540 4080 4650 4090
rect 4850 4080 4880 4090
rect 5070 4080 5100 4090
rect 5430 4080 5440 4090
rect 5670 4080 5690 4090
rect 6360 4080 6430 4090
rect 6500 4080 6510 4090
rect 7220 4080 7230 4090
rect 7500 4080 7520 4090
rect 7550 4080 7570 4090
rect 8780 4080 8790 4090
rect 9200 4080 9210 4090
rect 9610 4080 9650 4090
rect 9690 4080 9730 4090
rect 9940 4080 9950 4090
rect 2830 4070 2880 4080
rect 3020 4070 3050 4080
rect 3090 4070 3110 4080
rect 3240 4070 3250 4080
rect 4550 4070 4640 4080
rect 5080 4070 5110 4080
rect 5420 4070 5440 4080
rect 5670 4070 5710 4080
rect 6340 4070 6420 4080
rect 6500 4070 6510 4080
rect 7600 4070 7610 4080
rect 8790 4070 8800 4080
rect 9210 4070 9220 4080
rect 9940 4070 9970 4080
rect 2840 4060 2850 4070
rect 2870 4060 2880 4070
rect 2930 4060 2950 4070
rect 3010 4060 3020 4070
rect 3030 4060 3080 4070
rect 3130 4060 3140 4070
rect 3240 4060 3250 4070
rect 3260 4060 3270 4070
rect 4050 4060 4060 4070
rect 4550 4060 4640 4070
rect 5080 4060 5110 4070
rect 5420 4060 5430 4070
rect 5680 4060 5720 4070
rect 6320 4060 6410 4070
rect 6500 4060 6510 4070
rect 7210 4060 7220 4070
rect 7590 4060 7600 4070
rect 8790 4060 8800 4070
rect 2850 4050 2870 4060
rect 2940 4050 2950 4060
rect 2970 4050 2990 4060
rect 3010 4050 3060 4060
rect 3110 4050 3120 4060
rect 3150 4050 3160 4060
rect 3240 4050 3250 4060
rect 4050 4050 4060 4060
rect 4540 4050 4630 4060
rect 5080 4050 5110 4060
rect 5420 4050 5430 4060
rect 5700 4050 5730 4060
rect 6310 4050 6400 4060
rect 6500 4050 6510 4060
rect 7620 4050 7630 4060
rect 7660 4050 7670 4060
rect 8650 4050 8660 4060
rect 2870 4040 2880 4050
rect 2960 4040 2970 4050
rect 2980 4040 2990 4050
rect 3030 4040 3070 4050
rect 3140 4040 3150 4050
rect 4040 4040 4050 4050
rect 4540 4040 4630 4050
rect 5080 4040 5110 4050
rect 5420 4040 5430 4050
rect 5710 4040 5750 4050
rect 6300 4040 6390 4050
rect 6500 4040 6510 4050
rect 7200 4040 7210 4050
rect 7650 4040 7670 4050
rect 8770 4040 8790 4050
rect 2770 4030 2820 4040
rect 2870 4030 2880 4040
rect 2950 4030 2980 4040
rect 3050 4030 3100 4040
rect 3150 4030 3160 4040
rect 3170 4030 3180 4040
rect 4040 4030 4050 4040
rect 4540 4030 4620 4040
rect 4770 4030 4780 4040
rect 5090 4030 5110 4040
rect 5410 4030 5420 4040
rect 5720 4030 5760 4040
rect 6290 4030 6390 4040
rect 6500 4030 6510 4040
rect 7690 4030 7700 4040
rect 7710 4030 7720 4040
rect 8530 4030 8550 4040
rect 8610 4030 8620 4040
rect 8640 4030 8650 4040
rect 8660 4030 8670 4040
rect 2770 4020 2790 4030
rect 2810 4020 2820 4030
rect 2870 4020 2880 4030
rect 2950 4020 2980 4030
rect 3060 4020 3120 4030
rect 3160 4020 3180 4030
rect 4030 4020 4040 4030
rect 4550 4020 4620 4030
rect 4750 4020 4760 4030
rect 5100 4020 5120 4030
rect 5410 4020 5420 4030
rect 5730 4020 5820 4030
rect 6250 4020 6400 4030
rect 6500 4020 6520 4030
rect 6590 4020 6600 4030
rect 7710 4020 7720 4030
rect 7730 4020 7740 4030
rect 8530 4020 8540 4030
rect 8620 4020 8650 4030
rect 8670 4020 8680 4030
rect 2780 4010 2790 4020
rect 2950 4010 2980 4020
rect 3070 4010 3120 4020
rect 3180 4010 3190 4020
rect 4030 4010 4040 4020
rect 4550 4010 4620 4020
rect 4860 4010 4880 4020
rect 5100 4010 5130 4020
rect 5740 4010 5910 4020
rect 5920 4010 5940 4020
rect 6010 4010 6020 4020
rect 6240 4010 6410 4020
rect 6510 4010 6580 4020
rect 7190 4010 7200 4020
rect 7760 4010 7770 4020
rect 8440 4010 8450 4020
rect 8460 4010 8480 4020
rect 8500 4010 8510 4020
rect 8640 4010 8650 4020
rect 8680 4010 8690 4020
rect 2770 4000 2790 4010
rect 2840 4000 2850 4010
rect 2950 4000 2980 4010
rect 3080 4000 3130 4010
rect 3170 4000 3190 4010
rect 3220 4000 3230 4010
rect 4550 4000 4630 4010
rect 4710 4000 4720 4010
rect 4840 4000 4880 4010
rect 5100 4000 5140 4010
rect 5760 4000 5960 4010
rect 5970 4000 6010 4010
rect 6080 4000 6100 4010
rect 6220 4000 6400 4010
rect 7180 4000 7190 4010
rect 7750 4000 7760 4010
rect 7780 4000 7790 4010
rect 8380 4000 8390 4010
rect 8490 4000 8520 4010
rect 8530 4000 8540 4010
rect 8650 4000 8660 4010
rect 8700 4000 8710 4010
rect 8760 4000 8770 4010
rect 2770 3990 2800 4000
rect 2840 3990 2850 4000
rect 2950 3990 2970 4000
rect 3090 3990 3120 4000
rect 3130 3990 3150 4000
rect 3170 3990 3180 4000
rect 3220 3990 3230 4000
rect 3240 3990 3260 4000
rect 4010 3990 4030 4000
rect 4560 3990 4630 4000
rect 4690 3990 4700 4000
rect 4810 3990 4860 4000
rect 5110 3990 5150 4000
rect 5490 3990 5500 4000
rect 5780 3990 6110 4000
rect 6130 3990 6190 4000
rect 6200 3990 6300 4000
rect 6310 3990 6400 4000
rect 7170 3990 7180 4000
rect 7780 3990 7790 4000
rect 7810 3990 7820 4000
rect 8510 3990 8520 4000
rect 8530 3990 8540 4000
rect 8560 3990 8570 4000
rect 8660 3990 8670 4000
rect 8710 3990 8720 4000
rect 8730 3990 8740 4000
rect 8760 3990 8770 4000
rect 2770 3980 2800 3990
rect 2950 3980 2970 3990
rect 3100 3980 3130 3990
rect 3140 3980 3150 3990
rect 3170 3980 3190 3990
rect 3220 3980 3230 3990
rect 3250 3980 3260 3990
rect 4010 3980 4020 3990
rect 4220 3980 4250 3990
rect 4560 3980 4610 3990
rect 4620 3980 4630 3990
rect 4660 3980 4670 3990
rect 4790 3980 4820 3990
rect 4840 3980 4850 3990
rect 5120 3980 5150 3990
rect 5490 3980 5500 3990
rect 5800 3980 6280 3990
rect 6310 3980 6400 3990
rect 7160 3980 7180 3990
rect 8400 3980 8410 3990
rect 8430 3980 8450 3990
rect 8520 3980 8550 3990
rect 8700 3980 8710 3990
rect 8720 3980 8730 3990
rect 2890 3970 2900 3980
rect 2950 3970 2970 3980
rect 3130 3970 3140 3980
rect 3170 3970 3180 3980
rect 3190 3970 3200 3980
rect 3250 3970 3270 3980
rect 4000 3970 4010 3980
rect 4200 3970 4280 3980
rect 4560 3970 4580 3980
rect 4760 3970 4790 3980
rect 4830 3970 4840 3980
rect 5120 3970 5150 3980
rect 5830 3970 5860 3980
rect 5870 3970 5890 3980
rect 5900 3970 5930 3980
rect 5950 3970 6260 3980
rect 6310 3970 6400 3980
rect 7160 3970 7170 3980
rect 7830 3970 7840 3980
rect 8310 3970 8330 3980
rect 8420 3970 8450 3980
rect 8510 3970 8520 3980
rect 8550 3970 8570 3980
rect 8710 3970 8720 3980
rect 2890 3960 2900 3970
rect 2950 3960 2970 3970
rect 3130 3960 3140 3970
rect 3170 3960 3200 3970
rect 3990 3960 4010 3970
rect 4160 3960 4290 3970
rect 4720 3960 4770 3970
rect 4790 3960 4810 3970
rect 5130 3960 5160 3970
rect 5480 3960 5490 3970
rect 6000 3960 6230 3970
rect 6240 3960 6250 3970
rect 6310 3960 6400 3970
rect 7160 3960 7170 3970
rect 7890 3960 7900 3970
rect 8220 3960 8230 3970
rect 8320 3960 8330 3970
rect 8430 3960 8440 3970
rect 8730 3960 8750 3970
rect 2820 3950 2830 3960
rect 2940 3950 2970 3960
rect 3120 3950 3130 3960
rect 3160 3950 3190 3960
rect 3250 3950 3260 3960
rect 3980 3950 3990 3960
rect 4150 3950 4300 3960
rect 4700 3950 4750 3960
rect 4760 3950 4790 3960
rect 5140 3950 5170 3960
rect 5410 3950 5420 3960
rect 5430 3950 5450 3960
rect 5470 3950 5490 3960
rect 6040 3950 6060 3960
rect 6140 3950 6150 3960
rect 6320 3950 6400 3960
rect 7160 3950 7170 3960
rect 7880 3950 7890 3960
rect 8170 3950 8230 3960
rect 8300 3950 8320 3960
rect 8440 3950 8450 3960
rect 8570 3950 8580 3960
rect 9670 3950 9710 3960
rect 2950 3940 2970 3950
rect 3110 3940 3130 3950
rect 3150 3940 3190 3950
rect 3200 3940 3230 3950
rect 3250 3940 3260 3950
rect 3950 3940 3980 3950
rect 4140 3940 4300 3950
rect 4700 3940 4770 3950
rect 5150 3940 5180 3950
rect 5420 3940 5490 3950
rect 6320 3940 6400 3950
rect 7930 3940 7940 3950
rect 8130 3940 8140 3950
rect 8330 3940 8340 3950
rect 8410 3940 8420 3950
rect 8450 3940 8460 3950
rect 8500 3940 8510 3950
rect 8530 3940 8540 3950
rect 8650 3940 8660 3950
rect 8690 3940 8710 3950
rect 9670 3940 9680 3950
rect 2930 3930 2970 3940
rect 3050 3930 3060 3940
rect 3120 3930 3140 3940
rect 3160 3930 3170 3940
rect 3180 3930 3230 3940
rect 3250 3930 3270 3940
rect 3940 3930 3960 3940
rect 4120 3930 4200 3940
rect 4250 3930 4260 3940
rect 4270 3930 4310 3940
rect 5160 3930 5190 3940
rect 6320 3930 6400 3940
rect 7150 3930 7160 3940
rect 7920 3930 7930 3940
rect 7950 3930 7960 3940
rect 8110 3930 8120 3940
rect 8200 3930 8210 3940
rect 8260 3930 8280 3940
rect 8540 3930 8560 3940
rect 8580 3930 8590 3940
rect 8660 3930 8680 3940
rect 9640 3930 9650 3940
rect 9730 3930 9740 3940
rect 2930 3920 2960 3930
rect 3020 3920 3060 3930
rect 3100 3920 3160 3930
rect 3200 3920 3210 3930
rect 3220 3920 3230 3930
rect 3920 3920 3950 3930
rect 4110 3920 4160 3930
rect 4170 3920 4190 3930
rect 4260 3920 4320 3930
rect 5170 3920 5200 3930
rect 6320 3920 6330 3930
rect 6340 3920 6400 3930
rect 7950 3920 7960 3930
rect 8020 3920 8040 3930
rect 8050 3920 8060 3930
rect 8120 3920 8130 3930
rect 8140 3920 8160 3930
rect 8170 3920 8180 3930
rect 8190 3920 8200 3930
rect 8260 3920 8300 3930
rect 8440 3920 8450 3930
rect 8510 3920 8520 3930
rect 8550 3920 8560 3930
rect 8570 3920 8580 3930
rect 9630 3920 9640 3930
rect 9660 3920 9680 3930
rect 2860 3910 2880 3920
rect 2940 3910 2960 3920
rect 3030 3910 3150 3920
rect 3170 3910 3180 3920
rect 3190 3910 3200 3920
rect 3910 3910 3940 3920
rect 4090 3910 4190 3920
rect 4270 3910 4320 3920
rect 5180 3910 5200 3920
rect 6330 3910 6410 3920
rect 7960 3910 7970 3920
rect 8140 3910 8180 3920
rect 8190 3910 8200 3920
rect 8270 3910 8280 3920
rect 8520 3910 8530 3920
rect 8550 3910 8560 3920
rect 8640 3910 8650 3920
rect 8700 3910 8710 3920
rect 9610 3910 9630 3920
rect 9750 3910 9760 3920
rect 2860 3900 2920 3910
rect 2940 3900 2960 3910
rect 3030 3900 3140 3910
rect 3170 3900 3180 3910
rect 3190 3900 3200 3910
rect 3910 3900 3930 3910
rect 4090 3900 4140 3910
rect 4290 3900 4330 3910
rect 5180 3900 5220 3910
rect 6330 3900 6410 3910
rect 7980 3900 7990 3910
rect 8060 3900 8070 3910
rect 8190 3900 8200 3910
rect 8270 3900 8280 3910
rect 8510 3900 8550 3910
rect 9600 3900 9620 3910
rect 9780 3900 9790 3910
rect 2810 3890 2820 3900
rect 2860 3890 2920 3900
rect 2940 3890 2960 3900
rect 3000 3890 3120 3900
rect 3150 3890 3220 3900
rect 3900 3890 3920 3900
rect 4080 3890 4110 3900
rect 4300 3890 4330 3900
rect 5190 3890 5220 3900
rect 6330 3890 6410 3900
rect 8000 3890 8010 3900
rect 8190 3890 8200 3900
rect 8270 3890 8280 3900
rect 8340 3890 8350 3900
rect 8420 3890 8440 3900
rect 8530 3890 8540 3900
rect 8610 3890 8620 3900
rect 8650 3890 8660 3900
rect 8690 3890 8710 3900
rect 9560 3890 9590 3900
rect 9740 3890 9750 3900
rect 9760 3890 9770 3900
rect 2860 3880 2920 3890
rect 2930 3880 2980 3890
rect 3010 3880 3090 3890
rect 3130 3880 3140 3890
rect 3890 3880 3910 3890
rect 4050 3880 4110 3890
rect 4300 3880 4330 3890
rect 5190 3880 5220 3890
rect 6340 3880 6420 3890
rect 8010 3880 8020 3890
rect 8060 3880 8070 3890
rect 8200 3880 8210 3890
rect 8280 3880 8290 3890
rect 8340 3880 8350 3890
rect 8420 3880 8440 3890
rect 8460 3880 8470 3890
rect 8560 3880 8570 3890
rect 8640 3880 8650 3890
rect 8670 3880 8680 3890
rect 9460 3880 9470 3890
rect 9490 3880 9550 3890
rect 9720 3880 9730 3890
rect 9800 3880 9810 3890
rect 2870 3870 2980 3880
rect 2990 3870 3070 3880
rect 3890 3870 3900 3880
rect 4040 3870 4110 3880
rect 4310 3870 4330 3880
rect 5200 3870 5230 3880
rect 6340 3870 6430 3880
rect 7120 3870 7130 3880
rect 8040 3870 8050 3880
rect 8290 3870 8300 3880
rect 8320 3870 8340 3880
rect 8440 3870 8460 3880
rect 8470 3870 8480 3880
rect 8550 3870 8560 3880
rect 9460 3870 9480 3880
rect 9520 3870 9550 3880
rect 9720 3870 9730 3880
rect 9810 3870 9820 3880
rect 2800 3860 2820 3870
rect 2880 3860 2940 3870
rect 2950 3860 3070 3870
rect 3100 3860 3120 3870
rect 3160 3860 3180 3870
rect 3880 3860 3900 3870
rect 4050 3860 4110 3870
rect 4300 3860 4340 3870
rect 5200 3860 5230 3870
rect 6310 3860 6320 3870
rect 6340 3860 6440 3870
rect 8040 3860 8060 3870
rect 8220 3860 8230 3870
rect 8440 3860 8460 3870
rect 8620 3860 8640 3870
rect 8670 3860 8700 3870
rect 9430 3860 9440 3870
rect 9450 3860 9490 3870
rect 9530 3860 9550 3870
rect 9780 3860 9790 3870
rect 2880 3850 3050 3860
rect 3070 3850 3090 3860
rect 3140 3850 3170 3860
rect 4060 3850 4120 3860
rect 4280 3850 4340 3860
rect 5200 3850 5240 3860
rect 6340 3850 6500 3860
rect 8230 3850 8240 3860
rect 8440 3850 8470 3860
rect 8570 3850 8590 3860
rect 8620 3850 8650 3860
rect 9460 3850 9470 3860
rect 9560 3850 9570 3860
rect 2890 3840 3030 3850
rect 3060 3840 3080 3850
rect 3100 3840 3140 3850
rect 3150 3840 3160 3850
rect 3270 3840 3280 3850
rect 3870 3840 3880 3850
rect 4060 3840 4120 3850
rect 4280 3840 4340 3850
rect 5200 3840 5240 3850
rect 6340 3840 6510 3850
rect 8230 3840 8250 3850
rect 8460 3840 8480 3850
rect 8640 3840 8650 3850
rect 9730 3840 9740 3850
rect 9860 3840 9880 3850
rect 2690 3830 2700 3840
rect 2900 3830 2940 3840
rect 2950 3830 2980 3840
rect 3040 3830 3060 3840
rect 3070 3830 3100 3840
rect 3120 3830 3140 3840
rect 3150 3830 3160 3840
rect 3260 3830 3280 3840
rect 3870 3830 3880 3840
rect 4070 3830 4100 3840
rect 4290 3830 4340 3840
rect 5210 3830 5250 3840
rect 6340 3830 6510 3840
rect 8220 3830 8250 3840
rect 8610 3830 8620 3840
rect 8650 3830 8670 3840
rect 9730 3830 9740 3840
rect 9850 3830 9860 3840
rect 2690 3820 2700 3830
rect 2890 3820 2940 3830
rect 3000 3820 3070 3830
rect 3120 3820 3140 3830
rect 3260 3820 3270 3830
rect 3870 3820 3880 3830
rect 4060 3820 4090 3830
rect 4290 3820 4300 3830
rect 4320 3820 4330 3830
rect 5220 3820 5260 3830
rect 6310 3820 6520 3830
rect 7090 3820 7100 3830
rect 8090 3820 8100 3830
rect 8220 3820 8240 3830
rect 8480 3820 8490 3830
rect 8500 3820 8510 3830
rect 8600 3820 8610 3830
rect 8630 3820 8640 3830
rect 8670 3820 8680 3830
rect 9600 3820 9610 3830
rect 9790 3820 9800 3830
rect 2700 3810 2710 3820
rect 2980 3810 3010 3820
rect 3040 3810 3120 3820
rect 3180 3810 3200 3820
rect 3260 3810 3280 3820
rect 3870 3810 3880 3820
rect 4060 3810 4080 3820
rect 5220 3810 5260 3820
rect 6300 3810 6530 3820
rect 8180 3810 8190 3820
rect 8220 3810 8240 3820
rect 8440 3810 8460 3820
rect 8490 3810 8500 3820
rect 8610 3810 8620 3820
rect 9760 3810 9770 3820
rect 2700 3800 2720 3810
rect 2900 3800 2920 3810
rect 2960 3800 2990 3810
rect 3070 3800 3120 3810
rect 3150 3800 3160 3810
rect 3870 3800 3880 3810
rect 4040 3800 4060 3810
rect 4300 3800 4310 3810
rect 5230 3800 5270 3810
rect 6300 3800 6530 3810
rect 8130 3800 8140 3810
rect 8180 3800 8230 3810
rect 8240 3800 8270 3810
rect 8280 3800 8290 3810
rect 8300 3800 8310 3810
rect 8440 3800 8450 3810
rect 8470 3800 8480 3810
rect 8630 3800 8670 3810
rect 9820 3800 9830 3810
rect 2700 3790 2720 3800
rect 2730 3790 2740 3800
rect 2810 3790 2820 3800
rect 2900 3790 2920 3800
rect 2940 3790 2990 3800
rect 3070 3790 3100 3800
rect 3130 3790 3160 3800
rect 3260 3790 3270 3800
rect 3880 3790 3890 3800
rect 4030 3790 4050 3800
rect 4270 3790 4280 3800
rect 5220 3790 5270 3800
rect 6300 3790 6530 3800
rect 7070 3790 7080 3800
rect 8140 3790 8150 3800
rect 8190 3790 8200 3800
rect 8270 3790 8300 3800
rect 8450 3790 8460 3800
rect 8650 3790 8670 3800
rect 9610 3790 9620 3800
rect 9820 3790 9830 3800
rect 3090 3780 3110 3790
rect 3130 3780 3150 3790
rect 3890 3780 3910 3790
rect 4020 3780 4030 3790
rect 4250 3780 4260 3790
rect 5220 3780 5270 3790
rect 6300 3780 6530 3790
rect 8230 3780 8250 3790
rect 8320 3780 8350 3790
rect 8500 3780 8510 3790
rect 9810 3780 9820 3790
rect 2930 3770 2940 3780
rect 3050 3770 3110 3780
rect 3190 3770 3200 3780
rect 3890 3770 3920 3780
rect 4000 3770 4020 3780
rect 5230 3770 5280 3780
rect 6310 3770 6540 3780
rect 8190 3770 8220 3780
rect 8260 3770 8330 3780
rect 8360 3770 8370 3780
rect 8480 3770 8490 3780
rect 8510 3770 8520 3780
rect 9820 3770 9840 3780
rect 9850 3770 9860 3780
rect 2930 3760 2940 3770
rect 3030 3760 3050 3770
rect 3080 3760 3100 3770
rect 3120 3760 3130 3770
rect 3190 3760 3200 3770
rect 3270 3760 3280 3770
rect 3290 3760 3300 3770
rect 3900 3760 3940 3770
rect 3990 3760 4010 3770
rect 4190 3760 4200 3770
rect 5230 3760 5280 3770
rect 6320 3760 6530 3770
rect 7050 3760 7060 3770
rect 8220 3760 8320 3770
rect 8370 3760 8380 3770
rect 8500 3760 8510 3770
rect 9720 3760 9730 3770
rect 9750 3760 9770 3770
rect 9810 3760 9820 3770
rect 2770 3750 2780 3760
rect 2850 3750 2870 3760
rect 2900 3750 2940 3760
rect 3020 3750 3040 3760
rect 3060 3750 3120 3760
rect 3210 3750 3220 3760
rect 3270 3750 3280 3760
rect 3290 3750 3300 3760
rect 3890 3750 3930 3760
rect 3980 3750 4000 3760
rect 4150 3750 4160 3760
rect 5240 3750 5290 3760
rect 6330 3750 6350 3760
rect 6360 3750 6370 3760
rect 6440 3750 6530 3760
rect 8150 3750 8160 3760
rect 8170 3750 8320 3760
rect 8380 3750 8390 3760
rect 8520 3750 8530 3760
rect 8540 3750 8550 3760
rect 9660 3750 9670 3760
rect 9820 3750 9830 3760
rect 9860 3750 9870 3760
rect 2850 3740 2860 3750
rect 2890 3740 2950 3750
rect 3020 3740 3030 3750
rect 3060 3740 3110 3750
rect 3200 3740 3210 3750
rect 3270 3740 3280 3750
rect 3290 3740 3300 3750
rect 3890 3740 3930 3750
rect 3970 3740 3990 3750
rect 5240 3740 5290 3750
rect 6350 3740 6360 3750
rect 6440 3740 6530 3750
rect 8160 3740 8170 3750
rect 8210 3740 8310 3750
rect 8390 3740 8400 3750
rect 8530 3740 8560 3750
rect 9820 3740 9830 3750
rect 2890 3730 2960 3740
rect 3070 3730 3100 3740
rect 3120 3730 3150 3740
rect 3290 3730 3300 3740
rect 3890 3730 3920 3740
rect 3950 3730 3980 3740
rect 4220 3730 4250 3740
rect 5250 3730 5290 3740
rect 6440 3730 6540 3740
rect 7030 3730 7040 3740
rect 8170 3730 8180 3740
rect 8190 3730 8310 3740
rect 8390 3730 8410 3740
rect 8530 3730 8540 3740
rect 8570 3730 8580 3740
rect 9830 3730 9850 3740
rect 9880 3730 9900 3740
rect 9960 3730 9980 3740
rect 2880 3720 2960 3730
rect 3050 3720 3110 3730
rect 3120 3720 3170 3730
rect 3290 3720 3300 3730
rect 3890 3720 3910 3730
rect 3940 3720 3970 3730
rect 4050 3720 4060 3730
rect 4200 3720 4250 3730
rect 4850 3720 4870 3730
rect 5270 3720 5300 3730
rect 6450 3720 6530 3730
rect 8200 3720 8330 3730
rect 8360 3720 8370 3730
rect 8410 3720 8430 3730
rect 9690 3720 9700 3730
rect 9760 3720 9790 3730
rect 9960 3720 9990 3730
rect 2880 3710 2910 3720
rect 2920 3710 2970 3720
rect 2990 3710 3000 3720
rect 3080 3710 3100 3720
rect 3110 3710 3120 3720
rect 3130 3710 3180 3720
rect 3290 3710 3310 3720
rect 3880 3710 3890 3720
rect 3950 3710 3960 3720
rect 4030 3710 4040 3720
rect 4180 3710 4250 3720
rect 4830 3710 4910 3720
rect 5270 3710 5300 3720
rect 6450 3710 6540 3720
rect 8210 3710 8350 3720
rect 8380 3710 8390 3720
rect 8410 3710 8440 3720
rect 8540 3710 8550 3720
rect 8600 3710 8610 3720
rect 9690 3710 9700 3720
rect 9870 3710 9880 3720
rect 2900 3700 2950 3710
rect 3000 3700 3010 3710
rect 3020 3700 3030 3710
rect 3160 3700 3170 3710
rect 3280 3700 3300 3710
rect 3940 3700 3960 3710
rect 4020 3700 4030 3710
rect 4150 3700 4230 3710
rect 4840 3700 4940 3710
rect 5270 3700 5300 3710
rect 6450 3700 6540 3710
rect 8190 3700 8200 3710
rect 8220 3700 8250 3710
rect 8440 3700 8460 3710
rect 8610 3700 8620 3710
rect 9870 3700 9880 3710
rect 9950 3700 9960 3710
rect 2900 3690 2940 3700
rect 3040 3690 3060 3700
rect 3220 3690 3250 3700
rect 3290 3690 3300 3700
rect 3880 3690 3890 3700
rect 3930 3690 3960 3700
rect 4000 3690 4020 3700
rect 4120 3690 4190 3700
rect 4200 3690 4220 3700
rect 4850 3690 4870 3700
rect 4900 3690 4960 3700
rect 5280 3690 5310 3700
rect 6470 3690 6550 3700
rect 8470 3690 8480 3700
rect 8550 3690 8560 3700
rect 9870 3690 9880 3700
rect 3060 3680 3080 3690
rect 3090 3680 3110 3690
rect 3220 3680 3260 3690
rect 3290 3680 3300 3690
rect 3310 3680 3320 3690
rect 3880 3680 3890 3690
rect 3920 3680 3940 3690
rect 3990 3680 4000 3690
rect 4090 3680 4160 3690
rect 4180 3680 4200 3690
rect 4870 3680 4880 3690
rect 4940 3680 5000 3690
rect 5280 3680 5310 3690
rect 6470 3680 6550 3690
rect 8200 3680 8210 3690
rect 8390 3680 8400 3690
rect 8490 3680 8500 3690
rect 8610 3680 8620 3690
rect 9840 3680 9850 3690
rect 9920 3680 9930 3690
rect 3070 3670 3090 3680
rect 3210 3670 3240 3680
rect 3880 3670 3930 3680
rect 3980 3670 3990 3680
rect 4080 3670 4090 3680
rect 4130 3670 4180 3680
rect 4880 3670 4910 3680
rect 4960 3670 5030 3680
rect 5280 3670 5310 3680
rect 6470 3670 6550 3680
rect 8200 3670 8210 3680
rect 8500 3670 8510 3680
rect 8560 3670 8570 3680
rect 8600 3670 8610 3680
rect 3090 3660 3110 3670
rect 3210 3660 3230 3670
rect 3320 3660 3330 3670
rect 3970 3660 3980 3670
rect 4070 3660 4110 3670
rect 4910 3660 4930 3670
rect 4990 3660 5100 3670
rect 5290 3660 5320 3670
rect 6480 3660 6550 3670
rect 8400 3660 8410 3670
rect 8520 3660 8530 3670
rect 8570 3660 8580 3670
rect 9580 3660 9620 3670
rect 3130 3650 3140 3660
rect 3170 3650 3180 3660
rect 3200 3650 3230 3660
rect 3290 3650 3300 3660
rect 3320 3650 3340 3660
rect 3960 3650 3970 3660
rect 4920 3650 4960 3660
rect 5010 3650 5130 3660
rect 5290 3650 5320 3660
rect 6480 3650 6540 3660
rect 8210 3650 8220 3660
rect 8400 3650 8410 3660
rect 8540 3650 8550 3660
rect 9570 3650 9640 3660
rect 9870 3650 9890 3660
rect 3140 3640 3150 3650
rect 3180 3640 3240 3650
rect 3260 3640 3300 3650
rect 3320 3640 3340 3650
rect 4940 3640 4970 3650
rect 5030 3640 5130 3650
rect 5300 3640 5320 3650
rect 6460 3640 6540 3650
rect 6960 3640 6970 3650
rect 8220 3640 8230 3650
rect 8340 3640 8360 3650
rect 8390 3640 8400 3650
rect 9550 3640 9650 3650
rect 9870 3640 9880 3650
rect 3160 3630 3190 3640
rect 3200 3630 3230 3640
rect 3250 3630 3270 3640
rect 3290 3630 3300 3640
rect 3320 3630 3330 3640
rect 3340 3630 3350 3640
rect 3950 3630 3960 3640
rect 4950 3630 4990 3640
rect 5020 3630 5130 3640
rect 5290 3630 5320 3640
rect 6460 3630 6540 3640
rect 8240 3630 8250 3640
rect 8350 3630 8360 3640
rect 8370 3630 8380 3640
rect 8510 3630 8520 3640
rect 8530 3630 8550 3640
rect 9540 3630 9560 3640
rect 9570 3630 9590 3640
rect 9600 3630 9660 3640
rect 9890 3630 9910 3640
rect 3180 3620 3190 3630
rect 3210 3620 3240 3630
rect 3250 3620 3260 3630
rect 3290 3620 3300 3630
rect 3330 3620 3350 3630
rect 3940 3620 3950 3630
rect 4960 3620 5000 3630
rect 5030 3620 5130 3630
rect 5300 3620 5330 3630
rect 6460 3620 6540 3630
rect 8530 3620 8550 3630
rect 9530 3620 9550 3630
rect 9570 3620 9580 3630
rect 9620 3620 9660 3630
rect 9820 3620 9850 3630
rect 9930 3620 9940 3630
rect 3190 3610 3210 3620
rect 3240 3610 3260 3620
rect 3280 3610 3300 3620
rect 3350 3610 3360 3620
rect 3930 3610 3940 3620
rect 4970 3610 5130 3620
rect 5300 3610 5330 3620
rect 6450 3610 6530 3620
rect 6940 3610 6950 3620
rect 8260 3610 8270 3620
rect 8360 3610 8380 3620
rect 8520 3610 8530 3620
rect 9520 3610 9540 3620
rect 9560 3610 9570 3620
rect 9650 3610 9660 3620
rect 3220 3600 3230 3610
rect 3250 3600 3310 3610
rect 3920 3600 3930 3610
rect 4990 3600 5130 3610
rect 5300 3600 5330 3610
rect 6440 3600 6520 3610
rect 6930 3600 6940 3610
rect 8360 3600 8380 3610
rect 8510 3600 8520 3610
rect 9500 3600 9530 3610
rect 9550 3600 9560 3610
rect 9680 3600 9690 3610
rect 9910 3600 9920 3610
rect 3250 3590 3270 3600
rect 3310 3590 3320 3600
rect 3920 3590 3930 3600
rect 4790 3590 4820 3600
rect 5040 3590 5130 3600
rect 5300 3590 5330 3600
rect 6450 3590 6510 3600
rect 8280 3590 8290 3600
rect 8390 3590 8410 3600
rect 9470 3590 9500 3600
rect 9540 3590 9550 3600
rect 9670 3590 9680 3600
rect 9920 3590 9940 3600
rect 3250 3580 3280 3590
rect 3300 3580 3310 3590
rect 3340 3580 3360 3590
rect 3910 3580 3930 3590
rect 4770 3580 4780 3590
rect 4790 3580 4820 3590
rect 5060 3580 5130 3590
rect 5300 3580 5330 3590
rect 6430 3580 6510 3590
rect 8420 3580 8450 3590
rect 8500 3580 8510 3590
rect 9450 3580 9490 3590
rect 9530 3580 9540 3590
rect 9660 3580 9680 3590
rect 9740 3580 9750 3590
rect 3250 3570 3260 3580
rect 3270 3570 3280 3580
rect 3320 3570 3330 3580
rect 3340 3570 3360 3580
rect 3920 3570 3940 3580
rect 4750 3570 4770 3580
rect 4800 3570 4810 3580
rect 5070 3570 5140 3580
rect 5300 3570 5330 3580
rect 6400 3570 6420 3580
rect 6430 3570 6510 3580
rect 6910 3570 6920 3580
rect 8400 3570 8410 3580
rect 8490 3570 8500 3580
rect 9430 3570 9470 3580
rect 9530 3570 9540 3580
rect 9660 3570 9670 3580
rect 9720 3570 9740 3580
rect 3250 3560 3260 3570
rect 3320 3560 3330 3570
rect 3340 3560 3350 3570
rect 3370 3560 3380 3570
rect 3920 3560 3980 3570
rect 4710 3560 4720 3570
rect 4730 3560 4750 3570
rect 4790 3560 4810 3570
rect 5080 3560 5130 3570
rect 5300 3560 5330 3570
rect 6390 3560 6510 3570
rect 6900 3560 6910 3570
rect 8380 3560 8390 3570
rect 8440 3560 8450 3570
rect 8490 3560 8500 3570
rect 9410 3560 9440 3570
rect 9510 3560 9530 3570
rect 3260 3550 3270 3560
rect 3330 3550 3340 3560
rect 3350 3550 3360 3560
rect 3930 3550 3980 3560
rect 4690 3550 4740 3560
rect 4770 3550 4810 3560
rect 5100 3550 5140 3560
rect 5300 3550 5330 3560
rect 6370 3550 6510 3560
rect 6890 3550 6900 3560
rect 8380 3550 8390 3560
rect 8490 3550 8500 3560
rect 9300 3550 9320 3560
rect 9370 3550 9430 3560
rect 9500 3550 9510 3560
rect 9660 3550 9670 3560
rect 3340 3540 3360 3550
rect 3930 3540 3980 3550
rect 4690 3540 4730 3550
rect 4760 3540 4790 3550
rect 5050 3540 5070 3550
rect 5110 3540 5140 3550
rect 5300 3540 5340 3550
rect 6370 3540 6500 3550
rect 6880 3540 6890 3550
rect 8420 3540 8430 3550
rect 9280 3540 9420 3550
rect 9480 3540 9500 3550
rect 9650 3540 9660 3550
rect 3350 3530 3370 3540
rect 3930 3530 3990 3540
rect 4680 3530 4720 3540
rect 4750 3530 4780 3540
rect 5040 3530 5080 3540
rect 5110 3530 5140 3540
rect 5300 3530 5340 3540
rect 6350 3530 6480 3540
rect 8390 3530 8400 3540
rect 8410 3530 8420 3540
rect 9270 3530 9400 3540
rect 9470 3530 9480 3540
rect 3310 3520 3320 3530
rect 3350 3520 3360 3530
rect 3930 3520 3990 3530
rect 4340 3520 4360 3530
rect 4670 3520 4710 3530
rect 4740 3520 4780 3530
rect 5020 3520 5070 3530
rect 5110 3520 5130 3530
rect 5310 3520 5330 3530
rect 6350 3520 6360 3530
rect 6370 3520 6470 3530
rect 8350 3520 8360 3530
rect 8400 3520 8430 3530
rect 8440 3520 8450 3530
rect 8490 3520 8500 3530
rect 9260 3520 9390 3530
rect 9450 3520 9460 3530
rect 9630 3520 9660 3530
rect 3300 3510 3310 3520
rect 3330 3510 3340 3520
rect 3930 3510 3990 3520
rect 4330 3510 4370 3520
rect 4670 3510 4710 3520
rect 4730 3510 4780 3520
rect 5010 3510 5070 3520
rect 5310 3510 5340 3520
rect 6370 3510 6470 3520
rect 6860 3510 6870 3520
rect 8360 3510 8370 3520
rect 9230 3510 9240 3520
rect 9250 3510 9360 3520
rect 9430 3510 9440 3520
rect 9620 3510 9640 3520
rect 2540 3500 2550 3510
rect 3300 3500 3310 3510
rect 3400 3500 3410 3510
rect 3940 3500 3990 3510
rect 4320 3500 4370 3510
rect 4640 3500 4770 3510
rect 4990 3500 5010 3510
rect 5050 3500 5060 3510
rect 5310 3500 5340 3510
rect 6350 3500 6480 3510
rect 6850 3500 6860 3510
rect 8430 3500 8440 3510
rect 8500 3500 8510 3510
rect 9210 3500 9290 3510
rect 9410 3500 9420 3510
rect 9600 3500 9630 3510
rect 2480 3490 2490 3500
rect 2590 3490 2610 3500
rect 2630 3490 2680 3500
rect 3940 3490 3980 3500
rect 4300 3490 4370 3500
rect 4500 3490 4570 3500
rect 4600 3490 4760 3500
rect 4980 3490 4990 3500
rect 5050 3490 5060 3500
rect 5310 3490 5340 3500
rect 6340 3490 6480 3500
rect 8390 3490 8400 3500
rect 8510 3490 8520 3500
rect 9200 3490 9270 3500
rect 9380 3490 9390 3500
rect 9580 3490 9630 3500
rect 2420 3480 2450 3490
rect 2680 3480 2690 3490
rect 2750 3480 2760 3490
rect 3410 3480 3420 3490
rect 3940 3480 3980 3490
rect 4300 3480 4320 3490
rect 4350 3480 4380 3490
rect 4490 3480 4670 3490
rect 4680 3480 4750 3490
rect 4960 3480 4970 3490
rect 5040 3480 5050 3490
rect 5310 3480 5340 3490
rect 6330 3480 6470 3490
rect 8450 3480 8470 3490
rect 8520 3480 8530 3490
rect 9190 3480 9260 3490
rect 9360 3480 9380 3490
rect 9570 3480 9600 3490
rect 9620 3480 9630 3490
rect 2390 3470 2400 3480
rect 2700 3470 2720 3480
rect 2740 3470 2760 3480
rect 3320 3470 3330 3480
rect 3340 3470 3350 3480
rect 3950 3470 3990 3480
rect 4280 3470 4320 3480
rect 4350 3470 4390 3480
rect 4480 3470 4520 3480
rect 4620 3470 4630 3480
rect 4690 3470 4740 3480
rect 4940 3470 4960 3480
rect 5040 3470 5050 3480
rect 5310 3470 5340 3480
rect 6320 3470 6460 3480
rect 8470 3470 8480 3480
rect 9170 3470 9240 3480
rect 9320 3470 9340 3480
rect 9560 3470 9590 3480
rect 9610 3470 9620 3480
rect 2370 3460 2380 3470
rect 2750 3460 2770 3470
rect 2780 3460 2810 3470
rect 3340 3460 3360 3470
rect 3400 3460 3410 3470
rect 3950 3460 4000 3470
rect 4270 3460 4300 3470
rect 4350 3460 4410 3470
rect 4460 3460 4510 3470
rect 4690 3460 4740 3470
rect 4930 3460 4940 3470
rect 5030 3460 5040 3470
rect 5310 3460 5340 3470
rect 6320 3460 6450 3470
rect 8430 3460 8450 3470
rect 9160 3460 9220 3470
rect 9300 3460 9310 3470
rect 9540 3460 9570 3470
rect 9600 3460 9610 3470
rect 2340 3450 2360 3460
rect 2730 3450 2740 3460
rect 2810 3450 2850 3460
rect 3380 3450 3390 3460
rect 3420 3450 3430 3460
rect 3950 3450 4000 3460
rect 4270 3450 4310 3460
rect 4350 3450 4420 3460
rect 4440 3450 4480 3460
rect 4690 3450 4750 3460
rect 4910 3450 4920 3460
rect 5310 3450 5340 3460
rect 6320 3450 6440 3460
rect 8480 3450 8490 3460
rect 8530 3450 8540 3460
rect 9160 3450 9210 3460
rect 9280 3450 9290 3460
rect 9530 3450 9550 3460
rect 2290 3440 2320 3450
rect 2870 3440 2880 3450
rect 3440 3440 3450 3450
rect 3960 3440 4000 3450
rect 4270 3440 4300 3450
rect 4340 3440 4460 3450
rect 4680 3440 4750 3450
rect 4880 3440 4900 3450
rect 5300 3440 5330 3450
rect 6280 3440 6300 3450
rect 6320 3440 6380 3450
rect 6390 3440 6430 3450
rect 8530 3440 8540 3450
rect 9160 3440 9200 3450
rect 9260 3440 9270 3450
rect 9520 3440 9540 3450
rect 9580 3440 9600 3450
rect 2270 3430 2290 3440
rect 3440 3430 3450 3440
rect 3960 3430 4000 3440
rect 4270 3430 4300 3440
rect 4340 3430 4360 3440
rect 4380 3430 4410 3440
rect 4670 3430 4750 3440
rect 4860 3430 4900 3440
rect 5020 3430 5030 3440
rect 5300 3430 5330 3440
rect 6270 3430 6380 3440
rect 6390 3430 6430 3440
rect 8480 3430 8490 3440
rect 9150 3430 9190 3440
rect 9240 3430 9250 3440
rect 9450 3430 9460 3440
rect 9510 3430 9530 3440
rect 2250 3420 2260 3430
rect 2900 3420 2920 3430
rect 3970 3420 4000 3430
rect 4270 3420 4300 3430
rect 4330 3420 4350 3430
rect 4390 3420 4420 3430
rect 4660 3420 4750 3430
rect 4840 3420 4880 3430
rect 5020 3420 5030 3430
rect 5300 3420 5330 3430
rect 6240 3420 6370 3430
rect 6380 3420 6410 3430
rect 8490 3420 8510 3430
rect 9150 3420 9170 3430
rect 9440 3420 9470 3430
rect 9510 3420 9530 3430
rect 9570 3420 9580 3430
rect 2240 3410 2250 3420
rect 2900 3410 2960 3420
rect 3970 3410 4010 3420
rect 4260 3410 4290 3420
rect 4330 3410 4350 3420
rect 4390 3410 4430 3420
rect 4640 3410 4700 3420
rect 4710 3410 4740 3420
rect 4780 3410 4870 3420
rect 4950 3410 5000 3420
rect 5020 3410 5030 3420
rect 5310 3410 5330 3420
rect 6230 3410 6400 3420
rect 8500 3410 8510 3420
rect 9070 3410 9090 3420
rect 9120 3410 9160 3420
rect 9440 3410 9480 3420
rect 9510 3410 9530 3420
rect 9560 3410 9570 3420
rect 2230 3400 2240 3410
rect 2970 3400 2980 3410
rect 3980 3400 4010 3410
rect 4260 3400 4280 3410
rect 4330 3400 4350 3410
rect 4420 3400 4450 3410
rect 4610 3400 4620 3410
rect 4700 3400 4720 3410
rect 4740 3400 4850 3410
rect 4930 3400 4940 3410
rect 4980 3400 5000 3410
rect 5300 3400 5330 3410
rect 6210 3400 6400 3410
rect 8520 3400 8530 3410
rect 9060 3400 9090 3410
rect 9200 3400 9210 3410
rect 9430 3400 9520 3410
rect 9550 3400 9560 3410
rect 2220 3390 2230 3400
rect 3980 3390 4010 3400
rect 4260 3390 4280 3400
rect 4330 3390 4350 3400
rect 4420 3390 4460 3400
rect 4550 3390 4620 3400
rect 4630 3390 4640 3400
rect 4690 3390 4700 3400
rect 4740 3390 4750 3400
rect 4770 3390 4830 3400
rect 4920 3390 4930 3400
rect 4990 3390 5010 3400
rect 5300 3390 5330 3400
rect 6200 3390 6380 3400
rect 8530 3390 8540 3400
rect 9070 3390 9100 3400
rect 9420 3390 9520 3400
rect 9540 3390 9550 3400
rect 2200 3380 2220 3390
rect 3000 3380 3020 3390
rect 3490 3380 3510 3390
rect 3980 3380 4020 3390
rect 4260 3380 4270 3390
rect 4320 3380 4360 3390
rect 4430 3380 4440 3390
rect 4460 3380 4470 3390
rect 4480 3380 4620 3390
rect 4630 3380 4680 3390
rect 4720 3380 4750 3390
rect 4780 3380 4810 3390
rect 4990 3380 5010 3390
rect 5300 3380 5330 3390
rect 6200 3380 6380 3390
rect 6730 3380 6740 3390
rect 9090 3380 9110 3390
rect 9430 3380 9510 3390
rect 9530 3380 9540 3390
rect 9760 3380 9770 3390
rect 2190 3370 2210 3380
rect 3020 3370 3030 3380
rect 3490 3370 3510 3380
rect 3530 3370 3540 3380
rect 3990 3370 4020 3380
rect 4250 3370 4270 3380
rect 4330 3370 4360 3380
rect 4500 3370 4650 3380
rect 4710 3370 4740 3380
rect 4760 3370 4770 3380
rect 4890 3370 4910 3380
rect 4990 3370 5010 3380
rect 5300 3370 5330 3380
rect 6170 3370 6370 3380
rect 8520 3370 8530 3380
rect 9100 3370 9110 3380
rect 9420 3370 9500 3380
rect 9520 3370 9530 3380
rect 9740 3370 9750 3380
rect 9810 3370 9820 3380
rect 2180 3360 2190 3370
rect 3500 3360 3510 3370
rect 3990 3360 4040 3370
rect 4240 3360 4270 3370
rect 4320 3360 4360 3370
rect 4520 3360 4610 3370
rect 4700 3360 4710 3370
rect 4880 3360 4900 3370
rect 5000 3360 5020 3370
rect 5300 3360 5320 3370
rect 6160 3360 6360 3370
rect 8520 3360 8530 3370
rect 9080 3360 9110 3370
rect 9430 3360 9490 3370
rect 9810 3360 9820 3370
rect 2170 3350 2190 3360
rect 3510 3350 3520 3360
rect 4010 3350 4060 3360
rect 4070 3350 4080 3360
rect 4230 3350 4260 3360
rect 4320 3350 4360 3360
rect 4680 3350 4690 3360
rect 4870 3350 4880 3360
rect 4980 3350 4990 3360
rect 5000 3350 5020 3360
rect 5290 3350 5320 3360
rect 6160 3350 6340 3360
rect 6690 3350 6700 3360
rect 9080 3350 9100 3360
rect 9440 3350 9490 3360
rect 2150 3340 2180 3350
rect 3490 3340 3500 3350
rect 4010 3340 4150 3350
rect 4230 3340 4260 3350
rect 4320 3340 4350 3350
rect 4630 3340 4660 3350
rect 4860 3340 4870 3350
rect 5000 3340 5020 3350
rect 5290 3340 5320 3350
rect 6160 3340 6340 3350
rect 6680 3340 6690 3350
rect 8500 3340 8520 3350
rect 9060 3340 9080 3350
rect 9140 3340 9150 3350
rect 9430 3340 9480 3350
rect 9720 3340 9730 3350
rect 2140 3330 2170 3340
rect 3080 3330 3090 3340
rect 3520 3330 3530 3340
rect 4010 3330 4170 3340
rect 4210 3330 4250 3340
rect 4320 3330 4350 3340
rect 4580 3330 4630 3340
rect 4850 3330 4860 3340
rect 4990 3330 5000 3340
rect 5010 3330 5020 3340
rect 5290 3330 5320 3340
rect 6160 3330 6340 3340
rect 8490 3330 8510 3340
rect 9010 3330 9040 3340
rect 9430 3330 9460 3340
rect 9490 3330 9500 3340
rect 9690 3330 9700 3340
rect 2130 3320 2160 3330
rect 3500 3320 3510 3330
rect 4020 3320 4170 3330
rect 4190 3320 4200 3330
rect 4210 3320 4240 3330
rect 4320 3320 4350 3330
rect 4550 3320 4610 3330
rect 4840 3320 4850 3330
rect 4990 3320 5000 3330
rect 5010 3320 5020 3330
rect 5290 3320 5320 3330
rect 6170 3320 6310 3330
rect 8980 3320 9010 3330
rect 9020 3320 9060 3330
rect 9420 3320 9450 3330
rect 9480 3320 9490 3330
rect 9660 3320 9710 3330
rect 2120 3310 2160 3320
rect 3510 3310 3520 3320
rect 4030 3310 4180 3320
rect 4190 3310 4240 3320
rect 4320 3310 4350 3320
rect 4540 3310 4600 3320
rect 4780 3310 4830 3320
rect 4980 3310 5000 3320
rect 5290 3310 5310 3320
rect 6170 3310 6300 3320
rect 6650 3310 6670 3320
rect 8490 3310 8510 3320
rect 9050 3310 9070 3320
rect 9120 3310 9130 3320
rect 9340 3310 9370 3320
rect 9410 3310 9440 3320
rect 9470 3310 9480 3320
rect 9650 3310 9700 3320
rect 2110 3300 2140 3310
rect 3110 3300 3120 3310
rect 3510 3300 3520 3310
rect 3530 3300 3540 3310
rect 3580 3300 3590 3310
rect 4040 3300 4240 3310
rect 4320 3300 4340 3310
rect 4520 3300 4590 3310
rect 4760 3300 4780 3310
rect 4810 3300 4820 3310
rect 5290 3300 5310 3310
rect 6180 3300 6240 3310
rect 6270 3300 6290 3310
rect 6650 3300 6660 3310
rect 9060 3300 9070 3310
rect 9330 3300 9430 3310
rect 9460 3300 9470 3310
rect 9630 3300 9670 3310
rect 2110 3290 2140 3300
rect 3530 3290 3540 3300
rect 3550 3290 3570 3300
rect 4060 3290 4230 3300
rect 4310 3290 4340 3300
rect 4500 3290 4580 3300
rect 4740 3290 4760 3300
rect 4810 3290 4820 3300
rect 4970 3290 4980 3300
rect 5000 3290 5010 3300
rect 5290 3290 5310 3300
rect 6170 3290 6250 3300
rect 6640 3290 6670 3300
rect 9040 3290 9060 3300
rect 9100 3290 9120 3300
rect 9330 3290 9420 3300
rect 9450 3290 9460 3300
rect 9620 3290 9650 3300
rect 2100 3280 2130 3290
rect 3120 3280 3130 3290
rect 3530 3280 3540 3290
rect 4070 3280 4230 3290
rect 4310 3280 4340 3290
rect 4480 3280 4510 3290
rect 4520 3280 4550 3290
rect 4730 3280 4760 3290
rect 4800 3280 4810 3290
rect 4950 3280 4960 3290
rect 5290 3280 5310 3290
rect 6180 3280 6240 3290
rect 6590 3280 6620 3290
rect 6640 3280 6660 3290
rect 8470 3280 8480 3290
rect 8950 3280 8960 3290
rect 8970 3280 9010 3290
rect 9030 3280 9050 3290
rect 9080 3280 9120 3290
rect 9330 3280 9400 3290
rect 9440 3280 9450 3290
rect 9610 3280 9640 3290
rect 9720 3280 9740 3290
rect 2100 3270 2120 3280
rect 3120 3270 3130 3280
rect 4090 3270 4230 3280
rect 4310 3270 4350 3280
rect 4460 3270 4490 3280
rect 4700 3270 4750 3280
rect 4950 3270 4970 3280
rect 4990 3270 5000 3280
rect 5280 3270 5300 3280
rect 6190 3270 6240 3280
rect 6600 3270 6620 3280
rect 6640 3270 6660 3280
rect 8930 3270 8970 3280
rect 9030 3270 9050 3280
rect 9060 3270 9070 3280
rect 9100 3270 9120 3280
rect 9330 3270 9390 3280
rect 9430 3270 9440 3280
rect 9600 3270 9630 3280
rect 9680 3270 9730 3280
rect 2100 3260 2120 3270
rect 4110 3260 4230 3270
rect 4320 3260 4370 3270
rect 4430 3260 4450 3270
rect 4700 3260 4730 3270
rect 4750 3260 4760 3270
rect 4780 3260 4790 3270
rect 4940 3260 4960 3270
rect 4990 3260 5000 3270
rect 5280 3260 5300 3270
rect 6190 3260 6250 3270
rect 6590 3260 6610 3270
rect 6630 3260 6650 3270
rect 8460 3260 8470 3270
rect 9030 3260 9050 3270
rect 9100 3260 9120 3270
rect 9330 3260 9380 3270
rect 9420 3260 9440 3270
rect 9580 3260 9620 3270
rect 9690 3260 9720 3270
rect 2090 3250 2120 3260
rect 3130 3250 3140 3260
rect 3580 3250 3590 3260
rect 4110 3250 4230 3260
rect 4310 3250 4430 3260
rect 4660 3250 4670 3260
rect 4720 3250 4740 3260
rect 4750 3250 4780 3260
rect 4940 3250 4950 3260
rect 4990 3250 5000 3260
rect 5280 3250 5300 3260
rect 6200 3250 6250 3260
rect 6590 3250 6610 3260
rect 6630 3250 6650 3260
rect 9010 3250 9040 3260
rect 9090 3250 9110 3260
rect 9320 3250 9330 3260
rect 9340 3250 9370 3260
rect 9420 3250 9430 3260
rect 9570 3250 9600 3260
rect 9700 3250 9710 3260
rect 2080 3240 2110 3250
rect 3570 3240 3580 3250
rect 4120 3240 4230 3250
rect 4260 3240 4280 3250
rect 4340 3240 4400 3250
rect 4730 3240 4740 3250
rect 4750 3240 4760 3250
rect 4940 3240 4950 3250
rect 5280 3240 5300 3250
rect 6200 3240 6250 3250
rect 6510 3240 6520 3250
rect 6590 3240 6610 3250
rect 6620 3240 6650 3250
rect 9000 3240 9020 3250
rect 9090 3240 9100 3250
rect 9120 3240 9130 3250
rect 9310 3240 9330 3250
rect 9350 3240 9370 3250
rect 9410 3240 9420 3250
rect 9520 3240 9590 3250
rect 9700 3240 9710 3250
rect 2070 3230 2100 3240
rect 3140 3230 3150 3240
rect 3610 3230 3620 3240
rect 4120 3230 4240 3240
rect 4260 3230 4280 3240
rect 4650 3230 4660 3240
rect 4920 3230 4950 3240
rect 4980 3230 4990 3240
rect 5270 3230 5290 3240
rect 6200 3230 6260 3240
rect 6490 3230 6500 3240
rect 6590 3230 6610 3240
rect 6620 3230 6640 3240
rect 8980 3230 9000 3240
rect 9300 3230 9320 3240
rect 9350 3230 9360 3240
rect 9400 3230 9420 3240
rect 9490 3230 9570 3240
rect 9610 3230 9620 3240
rect 9630 3230 9640 3240
rect 9660 3230 9670 3240
rect 9940 3230 9950 3240
rect 2070 3220 2100 3230
rect 3600 3220 3610 3230
rect 4140 3220 4280 3230
rect 4650 3220 4660 3230
rect 4680 3220 4700 3230
rect 4920 3220 4940 3230
rect 5270 3220 5290 3230
rect 6210 3220 6270 3230
rect 6590 3220 6610 3230
rect 6620 3220 6650 3230
rect 8440 3220 8450 3230
rect 8960 3220 8980 3230
rect 9140 3220 9160 3230
rect 9290 3220 9300 3230
rect 9340 3220 9350 3230
rect 9390 3220 9410 3230
rect 9480 3220 9560 3230
rect 9600 3220 9610 3230
rect 9940 3220 9950 3230
rect 9970 3220 9980 3230
rect 2070 3210 2090 3220
rect 3150 3210 3160 3220
rect 3600 3210 3620 3220
rect 4150 3210 4280 3220
rect 4600 3210 4650 3220
rect 4910 3210 4930 3220
rect 5260 3210 5290 3220
rect 6210 3210 6270 3220
rect 6590 3210 6640 3220
rect 8940 3210 8960 3220
rect 9070 3210 9080 3220
rect 9150 3210 9170 3220
rect 9240 3210 9250 3220
rect 9280 3210 9300 3220
rect 9330 3210 9340 3220
rect 9380 3210 9400 3220
rect 9470 3210 9520 3220
rect 9940 3210 9950 3220
rect 2070 3200 2090 3210
rect 3600 3200 3610 3210
rect 4150 3200 4280 3210
rect 4540 3200 4620 3210
rect 4900 3200 4920 3210
rect 5270 3200 5280 3210
rect 6210 3200 6290 3210
rect 6430 3200 6440 3210
rect 6590 3200 6630 3210
rect 8430 3200 8440 3210
rect 8900 3200 8930 3210
rect 9060 3200 9070 3210
rect 9160 3200 9190 3210
rect 9200 3200 9280 3210
rect 9330 3200 9340 3210
rect 9370 3200 9400 3210
rect 9470 3200 9500 3210
rect 9590 3200 9600 3210
rect 9990 3200 9990 3210
rect 2070 3190 2090 3200
rect 3160 3190 3170 3200
rect 4160 3190 4290 3200
rect 4510 3190 4600 3200
rect 4890 3190 4920 3200
rect 4960 3190 4970 3200
rect 5270 3190 5280 3200
rect 6210 3190 6290 3200
rect 6400 3190 6410 3200
rect 6580 3190 6630 3200
rect 8820 3190 8890 3200
rect 9040 3190 9060 3200
rect 9200 3190 9210 3200
rect 9220 3190 9250 3200
rect 9260 3190 9280 3200
rect 9370 3190 9390 3200
rect 9460 3190 9510 3200
rect 2070 3180 2080 3190
rect 4170 3180 4300 3190
rect 4490 3180 4550 3190
rect 4580 3180 4590 3190
rect 4880 3180 4900 3190
rect 4950 3180 4960 3190
rect 5260 3180 5280 3190
rect 6220 3180 6290 3190
rect 6360 3180 6380 3190
rect 6580 3180 6630 3190
rect 9020 3180 9040 3190
rect 9260 3180 9280 3190
rect 9290 3180 9310 3190
rect 9370 3180 9380 3190
rect 9460 3180 9490 3190
rect 9590 3180 9600 3190
rect 2060 3170 2080 3180
rect 3170 3170 3180 3180
rect 4170 3170 4240 3180
rect 4250 3170 4260 3180
rect 4290 3170 4300 3180
rect 4490 3170 4570 3180
rect 4580 3170 4590 3180
rect 4880 3170 4900 3180
rect 4940 3170 4960 3180
rect 5260 3170 5280 3180
rect 6230 3170 6310 3180
rect 6340 3170 6360 3180
rect 6580 3170 6630 3180
rect 8980 3170 9030 3180
rect 9370 3170 9390 3180
rect 9460 3170 9490 3180
rect 9540 3170 9550 3180
rect 9560 3170 9590 3180
rect 9950 3170 9960 3180
rect 2060 3160 2080 3170
rect 3170 3160 3180 3170
rect 4170 3160 4230 3170
rect 4300 3160 4370 3170
rect 4380 3160 4400 3170
rect 4480 3160 4560 3170
rect 4570 3160 4590 3170
rect 4620 3160 4630 3170
rect 4870 3160 4890 3170
rect 4940 3160 4950 3170
rect 5260 3160 5270 3170
rect 5890 3160 5900 3170
rect 6240 3160 6310 3170
rect 6580 3160 6630 3170
rect 8950 3160 9020 3170
rect 9060 3160 9090 3170
rect 9320 3160 9350 3170
rect 9370 3160 9380 3170
rect 9440 3160 9480 3170
rect 9530 3160 9550 3170
rect 9630 3160 9640 3170
rect 9890 3160 9900 3170
rect 2060 3150 2080 3160
rect 3170 3150 3180 3160
rect 4180 3150 4230 3160
rect 4310 3150 4350 3160
rect 4400 3150 4410 3160
rect 4480 3150 4560 3160
rect 4580 3150 4600 3160
rect 4620 3150 4630 3160
rect 4860 3150 4870 3160
rect 4930 3150 4950 3160
rect 5260 3150 5270 3160
rect 6250 3150 6280 3160
rect 6580 3150 6630 3160
rect 8910 3150 8950 3160
rect 8980 3150 9000 3160
rect 9040 3150 9090 3160
rect 9300 3150 9350 3160
rect 9370 3150 9400 3160
rect 9420 3150 9470 3160
rect 9530 3150 9550 3160
rect 9590 3150 9600 3160
rect 9890 3150 9900 3160
rect 9970 3150 9980 3160
rect 2050 3140 2080 3150
rect 4190 3140 4230 3150
rect 4320 3140 4350 3150
rect 4420 3140 4430 3150
rect 4480 3140 4570 3150
rect 4590 3140 4640 3150
rect 4850 3140 4870 3150
rect 4920 3140 4940 3150
rect 5250 3140 5270 3150
rect 6580 3140 6620 3150
rect 8870 3140 8930 3150
rect 8970 3140 8990 3150
rect 9020 3140 9030 3150
rect 9080 3140 9090 3150
rect 9290 3140 9350 3150
rect 9360 3140 9460 3150
rect 9530 3140 9560 3150
rect 9600 3140 9610 3150
rect 9890 3140 9900 3150
rect 9910 3140 9920 3150
rect 2040 3130 2080 3140
rect 3170 3130 3180 3140
rect 4200 3130 4230 3140
rect 4330 3130 4340 3140
rect 4440 3130 4450 3140
rect 4490 3130 4580 3140
rect 4590 3130 4650 3140
rect 4830 3130 4850 3140
rect 4910 3130 4940 3140
rect 5250 3130 5260 3140
rect 6580 3130 6620 3140
rect 8840 3130 8890 3140
rect 8950 3130 8970 3140
rect 8990 3130 9010 3140
rect 9070 3130 9090 3140
rect 9270 3130 9350 3140
rect 9360 3130 9450 3140
rect 9540 3130 9560 3140
rect 9850 3130 9860 3140
rect 9920 3130 9930 3140
rect 2040 3120 2070 3130
rect 3170 3120 3180 3130
rect 4200 3120 4230 3130
rect 4520 3120 4580 3130
rect 4620 3120 4650 3130
rect 4820 3120 4840 3130
rect 4910 3120 4930 3130
rect 5250 3120 5260 3130
rect 6580 3120 6610 3130
rect 8820 3120 8840 3130
rect 8930 3120 8950 3130
rect 8970 3120 8990 3130
rect 9060 3120 9080 3130
rect 9220 3120 9440 3130
rect 9550 3120 9560 3130
rect 2040 3110 2070 3120
rect 3170 3110 3180 3120
rect 3870 3110 3880 3120
rect 4120 3110 4140 3120
rect 4210 3110 4240 3120
rect 4540 3110 4590 3120
rect 4810 3110 4830 3120
rect 4910 3110 4930 3120
rect 5240 3110 5250 3120
rect 6580 3110 6610 3120
rect 8920 3110 8940 3120
rect 8950 3110 8970 3120
rect 9050 3110 9070 3120
rect 9220 3110 9230 3120
rect 9280 3110 9340 3120
rect 9350 3110 9420 3120
rect 9540 3110 9550 3120
rect 9830 3110 9840 3120
rect 9880 3110 9890 3120
rect 9930 3110 9940 3120
rect 2040 3100 2070 3110
rect 3170 3100 3180 3110
rect 3870 3100 3880 3110
rect 4130 3100 4150 3110
rect 4220 3100 4240 3110
rect 4560 3100 4600 3110
rect 4780 3100 4810 3110
rect 4900 3100 4930 3110
rect 5240 3100 5250 3110
rect 6580 3100 6620 3110
rect 8900 3100 8920 3110
rect 8930 3100 8950 3110
rect 9040 3100 9060 3110
rect 9220 3100 9230 3110
rect 9270 3100 9280 3110
rect 9290 3100 9330 3110
rect 9340 3100 9400 3110
rect 9530 3100 9540 3110
rect 9880 3100 9890 3110
rect 2040 3090 2070 3100
rect 3170 3090 3180 3100
rect 3860 3090 3880 3100
rect 3890 3090 3900 3100
rect 4130 3090 4160 3100
rect 4230 3090 4250 3100
rect 4490 3090 4500 3100
rect 4590 3090 4620 3100
rect 4760 3090 4790 3100
rect 4890 3090 4920 3100
rect 6570 3090 6610 3100
rect 8420 3090 8430 3100
rect 8440 3090 8450 3100
rect 8880 3090 8930 3100
rect 9030 3090 9060 3100
rect 9230 3090 9390 3100
rect 9520 3090 9530 3100
rect 2030 3080 2070 3090
rect 3160 3080 3180 3090
rect 3870 3080 3900 3090
rect 4140 3080 4170 3090
rect 4240 3080 4270 3090
rect 4500 3080 4510 3090
rect 4620 3080 4750 3090
rect 4880 3080 4920 3090
rect 5230 3080 5240 3090
rect 6570 3080 6610 3090
rect 8430 3080 8440 3090
rect 8870 3080 8910 3090
rect 9020 3080 9060 3090
rect 9240 3080 9370 3090
rect 9510 3080 9520 3090
rect 2030 3070 2060 3080
rect 3170 3070 3180 3080
rect 3880 3070 3900 3080
rect 4150 3070 4180 3080
rect 4250 3070 4270 3080
rect 4510 3070 4520 3080
rect 4880 3070 4910 3080
rect 5210 3070 5240 3080
rect 6570 3070 6610 3080
rect 8370 3070 8380 3080
rect 8430 3070 8440 3080
rect 8880 3070 8890 3080
rect 9000 3070 9050 3080
rect 9260 3070 9360 3080
rect 9500 3070 9510 3080
rect 2020 3060 2060 3070
rect 3160 3060 3170 3070
rect 3770 3060 3800 3070
rect 3810 3060 3830 3070
rect 3880 3060 3910 3070
rect 4150 3060 4190 3070
rect 4260 3060 4290 3070
rect 4520 3060 4540 3070
rect 4870 3060 4900 3070
rect 5210 3060 5230 3070
rect 6570 3060 6610 3070
rect 8430 3060 8440 3070
rect 8970 3060 9050 3070
rect 9290 3060 9330 3070
rect 9500 3060 9510 3070
rect 9890 3060 9900 3070
rect 2020 3050 2060 3060
rect 3150 3050 3170 3060
rect 3760 3050 3770 3060
rect 3780 3050 3830 3060
rect 3870 3050 3910 3060
rect 4160 3050 4200 3060
rect 4280 3050 4300 3060
rect 4530 3050 4550 3060
rect 4860 3050 4900 3060
rect 5210 3050 5230 3060
rect 6570 3050 6600 3060
rect 8430 3050 8440 3060
rect 8950 3050 9040 3060
rect 9500 3050 9510 3060
rect 2020 3040 2050 3050
rect 3150 3040 3170 3050
rect 3790 3040 3830 3050
rect 3850 3040 3890 3050
rect 4160 3040 4210 3050
rect 4290 3040 4310 3050
rect 4530 3040 4570 3050
rect 4850 3040 4890 3050
rect 5210 3040 5220 3050
rect 6570 3040 6600 3050
rect 8930 3040 9040 3050
rect 2020 3030 2050 3040
rect 3150 3030 3170 3040
rect 3750 3030 3770 3040
rect 3780 3030 3880 3040
rect 4030 3030 4040 3040
rect 4180 3030 4220 3040
rect 4300 3030 4320 3040
rect 4530 3030 4590 3040
rect 4820 3030 4890 3040
rect 5210 3030 5220 3040
rect 6570 3030 6590 3040
rect 8350 3030 8360 3040
rect 8910 3030 9040 3040
rect 9490 3030 9500 3040
rect 9760 3030 9770 3040
rect 9900 3030 9910 3040
rect 2020 3020 2040 3030
rect 3150 3020 3170 3030
rect 3750 3020 3760 3030
rect 3770 3020 3800 3030
rect 3830 3020 3840 3030
rect 3860 3020 3890 3030
rect 4190 3020 4230 3030
rect 4310 3020 4340 3030
rect 4470 3020 4600 3030
rect 4800 3020 4890 3030
rect 5200 3020 5210 3030
rect 6570 3020 6590 3030
rect 8420 3020 8440 3030
rect 8900 3020 9040 3030
rect 9430 3020 9460 3030
rect 9480 3020 9490 3030
rect 9750 3020 9760 3030
rect 2020 3010 2040 3020
rect 3150 3010 3160 3020
rect 3780 3010 3790 3020
rect 3830 3010 3840 3020
rect 3870 3010 3890 3020
rect 3910 3010 3920 3020
rect 4040 3010 4050 3020
rect 4200 3010 4240 3020
rect 4320 3010 4350 3020
rect 4460 3010 4620 3020
rect 4780 3010 4890 3020
rect 5200 3010 5210 3020
rect 6560 3010 6590 3020
rect 8880 3010 8920 3020
rect 8930 3010 8940 3020
rect 8950 3010 9040 3020
rect 9420 3010 9490 3020
rect 9750 3010 9760 3020
rect 9800 3010 9820 3020
rect 9910 3010 9930 3020
rect 2010 3000 2040 3010
rect 3150 3000 3160 3010
rect 3850 3000 3870 3010
rect 3880 3000 3890 3010
rect 4030 3000 4050 3010
rect 4220 3000 4240 3010
rect 4330 3000 4360 3010
rect 4460 3000 4660 3010
rect 4770 3000 4890 3010
rect 5190 3000 5200 3010
rect 6560 3000 6590 3010
rect 8440 3000 8450 3010
rect 8740 3000 8770 3010
rect 8900 3000 9030 3010
rect 9420 3000 9480 3010
rect 9770 3000 9840 3010
rect 9860 3000 9890 3010
rect 9900 3000 9940 3010
rect 2020 2990 2040 3000
rect 3150 2990 3160 3000
rect 3880 2990 3900 3000
rect 4050 2990 4070 3000
rect 4330 2990 4370 3000
rect 4460 2990 4510 3000
rect 4520 2990 4620 3000
rect 4630 2990 4660 3000
rect 4760 2990 4880 3000
rect 5190 2990 5200 3000
rect 6560 2990 6590 3000
rect 8400 2990 8410 3000
rect 8710 2990 8850 3000
rect 8910 2990 9020 3000
rect 9380 2990 9400 3000
rect 9410 2990 9460 3000
rect 9780 2990 9880 3000
rect 2010 2980 2040 2990
rect 3150 2980 3160 2990
rect 3880 2980 3900 2990
rect 4050 2980 4070 2990
rect 4080 2980 4090 2990
rect 4350 2980 4370 2990
rect 4470 2980 4510 2990
rect 4520 2980 4660 2990
rect 4670 2980 4900 2990
rect 6560 2980 6580 2990
rect 8710 2980 8860 2990
rect 8920 2980 8940 2990
rect 8950 2980 9000 2990
rect 9360 2980 9460 2990
rect 9800 2980 9870 2990
rect 9950 2980 9960 2990
rect 2020 2970 2040 2980
rect 3140 2970 3160 2980
rect 3880 2970 3890 2980
rect 4050 2970 4060 2980
rect 4070 2970 4080 2980
rect 4350 2970 4390 2980
rect 4480 2970 4510 2980
rect 4520 2970 4900 2980
rect 5180 2970 5190 2980
rect 6560 2970 6580 2980
rect 8400 2970 8410 2980
rect 8710 2970 8850 2980
rect 8920 2970 8930 2980
rect 8950 2970 8990 2980
rect 9150 2970 9190 2980
rect 9330 2970 9460 2980
rect 9810 2970 9830 2980
rect 9910 2970 9940 2980
rect 2020 2960 2040 2970
rect 3140 2960 3160 2970
rect 4360 2960 4390 2970
rect 4490 2960 4510 2970
rect 4520 2960 4530 2970
rect 4540 2960 4910 2970
rect 6560 2960 6580 2970
rect 8310 2960 8320 2970
rect 8730 2960 8750 2970
rect 8760 2960 8830 2970
rect 8930 2960 8970 2970
rect 9130 2960 9190 2970
rect 9290 2960 9300 2970
rect 9320 2960 9460 2970
rect 9910 2960 9940 2970
rect 2010 2950 2040 2960
rect 3130 2950 3160 2960
rect 4370 2950 4420 2960
rect 4500 2950 4530 2960
rect 4560 2950 4900 2960
rect 5170 2950 5180 2960
rect 6560 2950 6580 2960
rect 8440 2950 8450 2960
rect 8900 2950 8910 2960
rect 8930 2950 8960 2960
rect 9130 2950 9190 2960
rect 9280 2950 9300 2960
rect 9310 2950 9450 2960
rect 9930 2950 9940 2960
rect 2010 2940 2040 2950
rect 3130 2940 3160 2950
rect 3830 2940 3840 2950
rect 3850 2940 3860 2950
rect 4000 2940 4020 2950
rect 4050 2940 4060 2950
rect 4380 2940 4430 2950
rect 4510 2940 4540 2950
rect 4560 2940 4950 2950
rect 5160 2940 5170 2950
rect 6570 2940 6580 2950
rect 8820 2940 8890 2950
rect 8910 2940 8940 2950
rect 9120 2940 9200 2950
rect 9270 2940 9440 2950
rect 9700 2940 9710 2950
rect 9930 2940 9950 2950
rect 2010 2930 2040 2940
rect 3140 2930 3160 2940
rect 3810 2930 3830 2940
rect 4400 2930 4440 2940
rect 4520 2930 4550 2940
rect 4560 2930 4930 2940
rect 5160 2930 5170 2940
rect 6560 2930 6580 2940
rect 8750 2930 8930 2940
rect 9110 2930 9210 2940
rect 9270 2930 9380 2940
rect 9420 2930 9430 2940
rect 9930 2930 9950 2940
rect 2010 2920 2040 2930
rect 3130 2920 3160 2930
rect 3830 2920 3850 2930
rect 3990 2920 4010 2930
rect 4030 2920 4040 2930
rect 4410 2920 4440 2930
rect 4530 2920 4930 2930
rect 4940 2920 4960 2930
rect 5150 2920 5160 2930
rect 6550 2920 6580 2930
rect 8690 2920 8980 2930
rect 9110 2920 9210 2930
rect 9250 2920 9370 2930
rect 9410 2920 9420 2930
rect 9700 2920 9710 2930
rect 9730 2920 9740 2930
rect 2010 2910 2030 2920
rect 3130 2910 3150 2920
rect 3990 2910 4000 2920
rect 4420 2910 4470 2920
rect 4540 2910 4930 2920
rect 5150 2910 5160 2920
rect 6550 2910 6570 2920
rect 8670 2910 8770 2920
rect 8780 2910 8960 2920
rect 9100 2910 9150 2920
rect 9170 2910 9220 2920
rect 9250 2910 9270 2920
rect 9290 2910 9370 2920
rect 9410 2910 9420 2920
rect 9720 2910 9730 2920
rect 9990 2910 9990 2920
rect 2010 2900 2020 2910
rect 3130 2900 3150 2910
rect 4220 2900 4230 2910
rect 4430 2900 4480 2910
rect 4540 2900 4940 2910
rect 5120 2900 5130 2910
rect 5140 2900 5150 2910
rect 6560 2900 6570 2910
rect 8640 2900 8750 2910
rect 8770 2900 8940 2910
rect 9100 2900 9150 2910
rect 9190 2900 9220 2910
rect 9250 2900 9270 2910
rect 9290 2900 9370 2910
rect 2010 2890 2020 2900
rect 3130 2890 3150 2900
rect 3940 2890 3950 2900
rect 4440 2890 4490 2900
rect 4540 2890 4950 2900
rect 4960 2890 5150 2900
rect 8630 2890 8790 2900
rect 8800 2890 8810 2900
rect 8830 2890 8860 2900
rect 8880 2890 8920 2900
rect 8990 2890 9000 2900
rect 9090 2890 9140 2900
rect 9200 2890 9230 2900
rect 9250 2890 9360 2900
rect 9400 2890 9410 2900
rect 9920 2890 9960 2900
rect 2000 2880 2020 2890
rect 3120 2880 3150 2890
rect 4240 2880 4250 2890
rect 4450 2880 5140 2890
rect 8620 2880 8710 2890
rect 8880 2880 8900 2890
rect 8960 2880 8990 2890
rect 9080 2880 9110 2890
rect 9200 2880 9230 2890
rect 9240 2880 9370 2890
rect 9930 2880 9950 2890
rect 2000 2870 2020 2880
rect 3130 2870 3150 2880
rect 3990 2870 4000 2880
rect 4240 2870 4250 2880
rect 4470 2870 5140 2880
rect 8250 2870 8260 2880
rect 8620 2870 8650 2880
rect 8680 2870 8690 2880
rect 8840 2870 8880 2880
rect 8940 2870 8990 2880
rect 9070 2870 9100 2880
rect 9180 2870 9380 2880
rect 9930 2870 9940 2880
rect 9960 2870 9990 2880
rect 2000 2860 2020 2870
rect 4240 2860 4250 2870
rect 4480 2860 5130 2870
rect 8640 2860 8650 2870
rect 8800 2860 8820 2870
rect 8900 2860 8990 2870
rect 9060 2860 9100 2870
rect 9180 2860 9360 2870
rect 9930 2860 9950 2870
rect 2010 2850 2020 2860
rect 3910 2850 3930 2860
rect 3980 2850 3990 2860
rect 4490 2850 5120 2860
rect 6550 2850 6560 2860
rect 7340 2850 7350 2860
rect 7380 2850 7390 2860
rect 8630 2850 8710 2860
rect 8740 2850 8780 2860
rect 8870 2850 8910 2860
rect 8930 2850 8980 2860
rect 9050 2850 9090 2860
rect 9180 2850 9360 2860
rect 9940 2850 9950 2860
rect 2000 2840 2020 2850
rect 3980 2840 3990 2850
rect 4510 2840 4630 2850
rect 4660 2840 5110 2850
rect 8620 2840 8710 2850
rect 8820 2840 8850 2850
rect 8920 2840 8960 2850
rect 9040 2840 9080 2850
rect 9180 2840 9370 2850
rect 9990 2840 9990 2850
rect 2000 2830 2010 2840
rect 4530 2830 4620 2840
rect 4680 2830 5090 2840
rect 8220 2830 8230 2840
rect 8610 2830 8670 2840
rect 8790 2830 8820 2840
rect 8910 2830 8940 2840
rect 9030 2830 9070 2840
rect 9180 2830 9360 2840
rect 9650 2830 9670 2840
rect 9990 2830 9990 2840
rect 2000 2820 2010 2830
rect 4080 2820 4090 2830
rect 4550 2820 4600 2830
rect 4730 2820 5080 2830
rect 8610 2820 8680 2830
rect 8750 2820 8790 2830
rect 8910 2820 8920 2830
rect 9020 2820 9060 2830
rect 9180 2820 9230 2830
rect 9260 2820 9360 2830
rect 9650 2820 9660 2830
rect 9670 2820 9680 2830
rect 9980 2820 9990 2830
rect 2000 2810 2020 2820
rect 3110 2810 3150 2820
rect 3980 2810 3990 2820
rect 4000 2810 4010 2820
rect 4750 2810 5070 2820
rect 7190 2810 7200 2820
rect 8610 2810 8740 2820
rect 8890 2810 8910 2820
rect 9010 2810 9060 2820
rect 9160 2810 9220 2820
rect 9290 2810 9360 2820
rect 9370 2810 9380 2820
rect 9560 2810 9570 2820
rect 9590 2810 9600 2820
rect 9610 2810 9630 2820
rect 9670 2810 9680 2820
rect 2000 2800 2010 2810
rect 3100 2800 3130 2810
rect 3970 2800 3980 2810
rect 4770 2800 5050 2810
rect 8620 2800 8720 2810
rect 8850 2800 8870 2810
rect 9000 2800 9060 2810
rect 9150 2800 9220 2810
rect 9290 2800 9350 2810
rect 9390 2800 9400 2810
rect 9550 2800 9560 2810
rect 9620 2800 9630 2810
rect 9640 2800 9660 2810
rect 9930 2800 9940 2810
rect 2000 2790 2010 2800
rect 3100 2790 3140 2800
rect 3970 2790 3980 2800
rect 4790 2790 5020 2800
rect 5070 2790 5100 2800
rect 7160 2790 7170 2800
rect 7560 2790 7570 2800
rect 8190 2790 8200 2800
rect 8620 2790 8700 2800
rect 8710 2790 8720 2800
rect 8800 2790 8840 2800
rect 8990 2790 9040 2800
rect 9130 2790 9220 2800
rect 9290 2790 9340 2800
rect 9410 2790 9420 2800
rect 9620 2790 9630 2800
rect 9650 2790 9670 2800
rect 9920 2790 9930 2800
rect 2000 2780 2010 2790
rect 3100 2780 3130 2790
rect 4260 2780 4270 2790
rect 4790 2780 4980 2790
rect 5060 2780 5100 2790
rect 8180 2780 8190 2790
rect 8630 2780 8660 2790
rect 8670 2780 8680 2790
rect 8760 2780 8800 2790
rect 8980 2780 9030 2790
rect 9090 2780 9200 2790
rect 9210 2780 9220 2790
rect 9280 2780 9340 2790
rect 9590 2780 9610 2790
rect 9630 2780 9640 2790
rect 9660 2780 9670 2790
rect 9920 2780 9930 2790
rect 1990 2770 2000 2780
rect 3100 2770 3130 2780
rect 3940 2770 3950 2780
rect 4810 2770 4950 2780
rect 5050 2770 5100 2780
rect 7600 2770 7610 2780
rect 8630 2770 8650 2780
rect 8660 2770 8670 2780
rect 8730 2770 8750 2780
rect 8960 2770 9020 2780
rect 9030 2770 9050 2780
rect 9070 2770 9180 2780
rect 9290 2770 9330 2780
rect 9400 2770 9410 2780
rect 9440 2770 9450 2780
rect 9920 2770 9930 2780
rect 9980 2770 9990 2780
rect 1990 2760 2030 2770
rect 3110 2760 3150 2770
rect 3880 2760 3890 2770
rect 4150 2760 4160 2770
rect 4820 2760 4940 2770
rect 5030 2760 5090 2770
rect 5100 2760 5120 2770
rect 6050 2760 6120 2770
rect 8640 2760 8730 2770
rect 8940 2760 9020 2770
rect 9060 2760 9170 2770
rect 9180 2760 9200 2770
rect 9290 2760 9330 2770
rect 9400 2760 9420 2770
rect 9470 2760 9480 2770
rect 9990 2760 9990 2770
rect 2000 2750 2040 2760
rect 3110 2750 3150 2760
rect 3930 2750 3940 2760
rect 4170 2750 4190 2760
rect 4840 2750 4860 2760
rect 4880 2750 4910 2760
rect 5020 2750 5090 2760
rect 5100 2750 5110 2760
rect 6040 2750 6130 2760
rect 8640 2750 8710 2760
rect 8930 2750 9010 2760
rect 9020 2750 9210 2760
rect 9270 2750 9320 2760
rect 9630 2750 9640 2760
rect 2010 2740 2040 2750
rect 3140 2740 3150 2750
rect 3930 2740 3940 2750
rect 4190 2740 4200 2750
rect 5020 2740 5100 2750
rect 5990 2740 6130 2750
rect 8640 2740 8690 2750
rect 8930 2740 8980 2750
rect 9030 2740 9210 2750
rect 9260 2740 9310 2750
rect 9510 2740 9520 2750
rect 9560 2740 9570 2750
rect 2000 2730 2030 2740
rect 3920 2730 3930 2740
rect 5040 2730 5120 2740
rect 5960 2730 5970 2740
rect 5990 2730 6130 2740
rect 7050 2730 7060 2740
rect 8660 2730 8680 2740
rect 8930 2730 8980 2740
rect 9020 2730 9210 2740
rect 9230 2730 9310 2740
rect 9580 2730 9590 2740
rect 9700 2730 9710 2740
rect 9900 2730 9910 2740
rect 2000 2720 2030 2730
rect 3910 2720 3920 2730
rect 3930 2720 3940 2730
rect 5030 2720 5120 2730
rect 5950 2720 6140 2730
rect 7030 2720 7040 2730
rect 8650 2720 8680 2730
rect 8940 2720 8980 2730
rect 9000 2720 9300 2730
rect 9600 2720 9610 2730
rect 9640 2720 9650 2730
rect 9900 2720 9910 2730
rect 2000 2710 2020 2720
rect 3900 2710 3930 2720
rect 5010 2710 5120 2720
rect 5940 2710 6150 2720
rect 7010 2710 7020 2720
rect 8650 2710 8690 2720
rect 8830 2710 8900 2720
rect 8940 2710 8980 2720
rect 8990 2710 9260 2720
rect 9280 2710 9290 2720
rect 9360 2710 9370 2720
rect 9400 2710 9410 2720
rect 9900 2710 9920 2720
rect 2000 2700 2020 2710
rect 3910 2700 3920 2710
rect 5010 2700 5120 2710
rect 5930 2700 6170 2710
rect 8650 2700 8690 2710
rect 8700 2700 8710 2710
rect 8740 2700 8750 2710
rect 8820 2700 8930 2710
rect 8940 2700 9240 2710
rect 9280 2700 9290 2710
rect 9910 2700 9940 2710
rect 2000 2690 2020 2700
rect 2800 2690 2820 2700
rect 3130 2690 3150 2700
rect 4990 2690 5000 2700
rect 5010 2690 5120 2700
rect 5890 2690 6180 2700
rect 8640 2690 8760 2700
rect 8810 2690 8930 2700
rect 9020 2690 9220 2700
rect 9270 2690 9280 2700
rect 9930 2690 9940 2700
rect 1990 2680 2000 2690
rect 2790 2680 2830 2690
rect 3130 2680 3150 2690
rect 3900 2680 3930 2690
rect 4240 2680 4250 2690
rect 5000 2680 5120 2690
rect 5880 2680 6190 2690
rect 8640 2680 8780 2690
rect 8800 2680 8950 2690
rect 9080 2680 9170 2690
rect 9260 2680 9270 2690
rect 9940 2680 9960 2690
rect 1980 2670 2000 2680
rect 2260 2670 2410 2680
rect 2790 2670 2860 2680
rect 2920 2670 2990 2680
rect 3130 2670 3150 2680
rect 3900 2670 3910 2680
rect 5000 2670 5110 2680
rect 5880 2670 6190 2680
rect 8090 2670 8100 2680
rect 8650 2670 8980 2680
rect 9250 2670 9260 2680
rect 9650 2670 9660 2680
rect 9960 2670 9970 2680
rect 1980 2660 1990 2670
rect 2210 2660 2260 2670
rect 2330 2660 2420 2670
rect 2770 2660 2930 2670
rect 3050 2660 3140 2670
rect 4200 2660 4210 2670
rect 4990 2660 5090 2670
rect 5100 2660 5110 2670
rect 5850 2660 6200 2670
rect 8080 2660 8090 2670
rect 8640 2660 8780 2670
rect 8830 2660 9000 2670
rect 9240 2660 9250 2670
rect 9970 2660 9980 2670
rect 1970 2650 1990 2660
rect 2170 2650 2200 2660
rect 2370 2650 2440 2660
rect 2770 2650 2890 2660
rect 3110 2650 3120 2660
rect 3130 2650 3140 2660
rect 3900 2650 3910 2660
rect 4980 2650 5090 2660
rect 5820 2650 5830 2660
rect 5850 2650 6210 2660
rect 8660 2650 8760 2660
rect 8770 2650 8790 2660
rect 8850 2650 9010 2660
rect 9980 2650 9990 2660
rect 1970 2640 1990 2650
rect 2130 2640 2160 2650
rect 2390 2640 2440 2650
rect 2760 2640 2870 2650
rect 3040 2640 3050 2650
rect 3900 2640 3910 2650
rect 4200 2640 4210 2650
rect 4980 2640 5070 2650
rect 5830 2640 6220 2650
rect 6910 2640 6920 2650
rect 7170 2640 7180 2650
rect 8060 2640 8070 2650
rect 8660 2640 8750 2650
rect 8770 2640 8780 2650
rect 8870 2640 9020 2650
rect 9960 2640 9990 2650
rect 1970 2630 1980 2640
rect 2110 2630 2140 2640
rect 2200 2630 2220 2640
rect 2250 2630 2280 2640
rect 2390 2630 2440 2640
rect 2760 2630 2860 2640
rect 2930 2630 2940 2640
rect 3060 2630 3080 2640
rect 3900 2630 3930 2640
rect 4200 2630 4210 2640
rect 4950 2630 5060 2640
rect 5830 2630 6230 2640
rect 6900 2630 6910 2640
rect 8730 2630 8740 2640
rect 8890 2630 9030 2640
rect 9200 2630 9210 2640
rect 9990 2630 9990 2640
rect 1960 2620 1980 2630
rect 2090 2620 2110 2630
rect 2180 2620 2190 2630
rect 2270 2620 2280 2630
rect 2400 2620 2430 2630
rect 2760 2620 2850 2630
rect 2910 2620 2920 2630
rect 2960 2620 2980 2630
rect 2990 2620 3000 2630
rect 3080 2620 3090 2630
rect 3920 2620 3930 2630
rect 4200 2620 4210 2630
rect 4260 2620 4270 2630
rect 4950 2620 5040 2630
rect 5830 2620 5850 2630
rect 5860 2620 6230 2630
rect 6890 2620 6900 2630
rect 8900 2620 9040 2630
rect 9190 2620 9200 2630
rect 9750 2620 9760 2630
rect 1950 2610 1970 2620
rect 2070 2610 2090 2620
rect 2140 2610 2180 2620
rect 2190 2610 2200 2620
rect 2220 2610 2260 2620
rect 2400 2610 2430 2620
rect 2760 2610 2840 2620
rect 2910 2610 2930 2620
rect 3040 2610 3050 2620
rect 3080 2610 3090 2620
rect 3930 2610 3940 2620
rect 4260 2610 4270 2620
rect 4950 2610 4970 2620
rect 5000 2610 5010 2620
rect 5820 2610 5830 2620
rect 5840 2610 6240 2620
rect 8910 2610 9050 2620
rect 9190 2610 9200 2620
rect 9770 2610 9780 2620
rect 9860 2610 9870 2620
rect 1950 2600 1970 2610
rect 2060 2600 2080 2610
rect 2130 2600 2170 2610
rect 2410 2600 2430 2610
rect 2760 2600 2830 2610
rect 3930 2600 3940 2610
rect 5810 2600 5820 2610
rect 5830 2600 5900 2610
rect 5910 2600 6250 2610
rect 7200 2600 7230 2610
rect 8870 2600 8900 2610
rect 8940 2600 9050 2610
rect 9790 2600 9800 2610
rect 9880 2600 9890 2610
rect 1950 2590 1970 2600
rect 2040 2590 2060 2600
rect 2410 2590 2430 2600
rect 2770 2590 2810 2600
rect 2820 2590 2830 2600
rect 3920 2590 3940 2600
rect 4080 2590 4090 2600
rect 5790 2590 5830 2600
rect 5840 2590 5860 2600
rect 5880 2590 6250 2600
rect 7200 2590 7230 2600
rect 8860 2590 8940 2600
rect 8960 2590 9050 2600
rect 9170 2590 9190 2600
rect 9810 2590 9820 2600
rect 9870 2590 9880 2600
rect 9900 2590 9910 2600
rect 1940 2580 1970 2590
rect 2040 2580 2050 2590
rect 2090 2580 2120 2590
rect 2410 2580 2420 2590
rect 2810 2580 2840 2590
rect 3920 2580 3940 2590
rect 4060 2580 4080 2590
rect 4200 2580 4220 2590
rect 4250 2580 4260 2590
rect 5800 2580 5810 2590
rect 5840 2580 5880 2590
rect 5890 2580 6260 2590
rect 7210 2580 7240 2590
rect 7270 2580 7280 2590
rect 8860 2580 8940 2590
rect 8970 2580 9010 2590
rect 9020 2580 9030 2590
rect 9160 2580 9180 2590
rect 9830 2580 9840 2590
rect 9890 2580 9900 2590
rect 9920 2580 9930 2590
rect 1930 2570 1940 2580
rect 2020 2570 2040 2580
rect 2100 2570 2110 2580
rect 2410 2570 2420 2580
rect 2830 2570 2840 2580
rect 3900 2570 3910 2580
rect 4060 2570 4070 2580
rect 4220 2570 4230 2580
rect 4240 2570 4250 2580
rect 5780 2570 5790 2580
rect 5840 2570 6270 2580
rect 7210 2570 7250 2580
rect 7270 2570 7290 2580
rect 7990 2570 8000 2580
rect 8870 2570 8940 2580
rect 9000 2570 9020 2580
rect 9150 2570 9190 2580
rect 9490 2570 9500 2580
rect 9520 2570 9530 2580
rect 9850 2570 9860 2580
rect 9910 2570 9920 2580
rect 9940 2570 9950 2580
rect 1930 2560 1940 2570
rect 2010 2560 2030 2570
rect 2410 2560 2420 2570
rect 2890 2560 2900 2570
rect 4040 2560 4060 2570
rect 4090 2560 4100 2570
rect 4180 2560 4200 2570
rect 4220 2560 4250 2570
rect 5770 2560 5810 2570
rect 5820 2560 6270 2570
rect 7140 2560 7160 2570
rect 7220 2560 7290 2570
rect 8880 2560 8940 2570
rect 8980 2560 9000 2570
rect 9020 2560 9040 2570
rect 9150 2560 9180 2570
rect 9320 2560 9330 2570
rect 9400 2560 9420 2570
rect 9470 2560 9480 2570
rect 9540 2560 9550 2570
rect 9870 2560 9880 2570
rect 9930 2560 9940 2570
rect 1930 2550 1940 2560
rect 2000 2550 2020 2560
rect 2330 2550 2360 2560
rect 2820 2550 2830 2560
rect 2900 2550 2910 2560
rect 4000 2550 4010 2560
rect 4040 2550 4060 2560
rect 4070 2550 4100 2560
rect 4160 2550 4170 2560
rect 4230 2550 4270 2560
rect 5790 2550 6280 2560
rect 7140 2550 7150 2560
rect 7160 2550 7170 2560
rect 7220 2550 7250 2560
rect 7270 2550 7300 2560
rect 8890 2550 8930 2560
rect 8980 2550 9010 2560
rect 9030 2550 9050 2560
rect 9160 2550 9180 2560
rect 9470 2550 9480 2560
rect 9890 2550 9900 2560
rect 9950 2550 9960 2560
rect 1930 2540 1940 2550
rect 1990 2540 2000 2550
rect 2330 2540 2370 2550
rect 2820 2540 2830 2550
rect 2880 2540 2890 2550
rect 2900 2540 2910 2550
rect 3930 2540 3960 2550
rect 4080 2540 4100 2550
rect 5770 2540 6280 2550
rect 7170 2540 7180 2550
rect 7280 2540 7300 2550
rect 8890 2540 8910 2550
rect 8990 2540 9060 2550
rect 9160 2540 9180 2550
rect 9350 2540 9360 2550
rect 9410 2540 9420 2550
rect 9580 2540 9590 2550
rect 9910 2540 9920 2550
rect 9970 2540 9980 2550
rect 1930 2530 1940 2540
rect 1980 2530 1990 2540
rect 2330 2530 2350 2540
rect 2870 2530 2880 2540
rect 2890 2530 2910 2540
rect 2940 2530 2950 2540
rect 3030 2530 3040 2540
rect 3110 2530 3140 2540
rect 3930 2530 3950 2540
rect 4080 2530 4090 2540
rect 4100 2530 4110 2540
rect 4130 2530 4160 2540
rect 5770 2530 6290 2540
rect 7180 2530 7190 2540
rect 7240 2530 7250 2540
rect 7280 2530 7310 2540
rect 8900 2530 8910 2540
rect 8990 2530 9060 2540
rect 9150 2530 9170 2540
rect 9430 2530 9440 2540
rect 9600 2530 9610 2540
rect 9930 2530 9940 2540
rect 1930 2520 1940 2530
rect 1970 2520 1990 2530
rect 2390 2520 2400 2530
rect 2860 2520 2900 2530
rect 3140 2520 3180 2530
rect 4050 2520 4060 2530
rect 4090 2520 4100 2530
rect 4110 2520 4150 2530
rect 5770 2520 6300 2530
rect 7180 2520 7210 2530
rect 7250 2520 7260 2530
rect 7300 2520 7310 2530
rect 7930 2520 7940 2530
rect 8880 2520 8890 2530
rect 8990 2520 9060 2530
rect 9150 2520 9170 2530
rect 9620 2520 9630 2530
rect 9950 2520 9960 2530
rect 1930 2510 1950 2520
rect 1970 2510 1980 2520
rect 2030 2510 2110 2520
rect 2160 2510 2240 2520
rect 2250 2510 2270 2520
rect 2300 2510 2380 2520
rect 3970 2510 3980 2520
rect 4000 2510 4010 2520
rect 4020 2510 4070 2520
rect 4090 2510 4110 2520
rect 4120 2510 4130 2520
rect 5750 2510 5760 2520
rect 5770 2510 6300 2520
rect 7200 2510 7220 2520
rect 7260 2510 7270 2520
rect 7310 2510 7320 2520
rect 8830 2510 8860 2520
rect 8870 2510 8900 2520
rect 8980 2510 9050 2520
rect 9150 2510 9160 2520
rect 9480 2510 9490 2520
rect 1930 2500 1970 2510
rect 2000 2500 2010 2510
rect 2070 2500 2090 2510
rect 2320 2500 2350 2510
rect 3930 2500 3940 2510
rect 3980 2500 4030 2510
rect 4050 2500 4090 2510
rect 4100 2500 4110 2510
rect 5770 2500 6310 2510
rect 7220 2500 7230 2510
rect 7270 2500 7280 2510
rect 7320 2500 7330 2510
rect 8830 2500 8890 2510
rect 8970 2500 9080 2510
rect 9140 2500 9160 2510
rect 9280 2500 9290 2510
rect 9410 2500 9420 2510
rect 9580 2500 9590 2510
rect 9990 2500 9990 2510
rect 1930 2490 1980 2500
rect 3200 2490 3210 2500
rect 3980 2490 3990 2500
rect 4010 2490 4020 2500
rect 4060 2490 4090 2500
rect 5640 2490 5660 2500
rect 5760 2490 6310 2500
rect 7230 2490 7260 2500
rect 7270 2490 7290 2500
rect 7320 2490 7330 2500
rect 7880 2490 7890 2500
rect 8840 2490 8890 2500
rect 8940 2490 9090 2500
rect 9130 2490 9150 2500
rect 9260 2490 9270 2500
rect 9600 2490 9610 2500
rect 9680 2490 9690 2500
rect 1930 2480 1950 2490
rect 4010 2480 4020 2490
rect 5640 2480 5660 2490
rect 5760 2480 6320 2490
rect 7240 2480 7290 2490
rect 7330 2480 7350 2490
rect 7860 2480 7870 2490
rect 8940 2480 9100 2490
rect 9110 2480 9140 2490
rect 9250 2480 9260 2490
rect 9700 2480 9710 2490
rect 1920 2470 1940 2480
rect 5610 2470 5660 2480
rect 5750 2470 6320 2480
rect 7250 2470 7260 2480
rect 7270 2470 7300 2480
rect 7340 2470 7350 2480
rect 8950 2470 9130 2480
rect 1910 2460 1930 2470
rect 3910 2460 3920 2470
rect 5590 2460 5650 2470
rect 5740 2460 6330 2470
rect 7260 2460 7270 2470
rect 7350 2460 7360 2470
rect 8970 2460 9100 2470
rect 9500 2460 9510 2470
rect 1920 2450 1930 2460
rect 3230 2450 3240 2460
rect 5560 2450 5650 2460
rect 5740 2450 6340 2460
rect 9470 2450 9480 2460
rect 1910 2440 1920 2450
rect 2140 2440 2180 2450
rect 5560 2440 5610 2450
rect 5630 2440 5660 2450
rect 5720 2440 5730 2450
rect 5750 2440 6340 2450
rect 6770 2440 6800 2450
rect 7280 2440 7290 2450
rect 7360 2440 7380 2450
rect 9290 2440 9300 2450
rect 9430 2440 9440 2450
rect 9480 2440 9490 2450
rect 9690 2440 9700 2450
rect 9730 2440 9740 2450
rect 9770 2440 9780 2450
rect 1910 2430 1920 2440
rect 2140 2430 2230 2440
rect 3240 2430 3250 2440
rect 4010 2430 4030 2440
rect 5570 2430 5650 2440
rect 5710 2430 6350 2440
rect 6750 2430 6760 2440
rect 6780 2430 6810 2440
rect 7300 2430 7310 2440
rect 7380 2430 7390 2440
rect 7420 2430 7430 2440
rect 9440 2430 9450 2440
rect 9670 2430 9680 2440
rect 9700 2430 9710 2440
rect 1910 2420 1920 2430
rect 3250 2420 3260 2430
rect 5550 2420 5640 2430
rect 5700 2420 6350 2430
rect 6750 2420 6850 2430
rect 7320 2420 7330 2430
rect 7390 2420 7430 2430
rect 9220 2420 9230 2430
rect 9490 2420 9520 2430
rect 9540 2420 9560 2430
rect 9660 2420 9680 2430
rect 3240 2410 3260 2420
rect 5550 2410 5560 2420
rect 5570 2410 5640 2420
rect 5690 2410 6360 2420
rect 6750 2410 6850 2420
rect 7390 2410 7430 2420
rect 9230 2410 9250 2420
rect 9330 2410 9340 2420
rect 9560 2410 9570 2420
rect 9640 2410 9650 2420
rect 9680 2410 9690 2420
rect 3240 2400 3260 2410
rect 5560 2400 5620 2410
rect 5690 2400 6360 2410
rect 6740 2400 6870 2410
rect 7420 2400 7440 2410
rect 8950 2400 8960 2410
rect 9250 2400 9260 2410
rect 9480 2400 9490 2410
rect 9590 2400 9600 2410
rect 9830 2400 9850 2410
rect 5570 2390 5580 2400
rect 5690 2390 6370 2400
rect 6740 2390 6890 2400
rect 7370 2390 7380 2400
rect 7430 2390 7440 2400
rect 9320 2390 9330 2400
rect 9470 2390 9480 2400
rect 9590 2390 9600 2400
rect 9840 2390 9850 2400
rect 1900 2380 1910 2390
rect 3250 2380 3260 2390
rect 5690 2380 6370 2390
rect 6740 2380 6900 2390
rect 7430 2380 7450 2390
rect 9270 2380 9280 2390
rect 9550 2380 9560 2390
rect 9700 2380 9710 2390
rect 1900 2370 1910 2380
rect 3250 2370 3270 2380
rect 5700 2370 6380 2380
rect 6740 2370 6900 2380
rect 7400 2370 7410 2380
rect 7440 2370 7460 2380
rect 8400 2370 8410 2380
rect 9150 2370 9160 2380
rect 9200 2370 9210 2380
rect 9450 2370 9460 2380
rect 9530 2370 9540 2380
rect 9570 2370 9580 2380
rect 9590 2370 9600 2380
rect 9700 2370 9710 2380
rect 1890 2360 1910 2370
rect 3260 2360 3280 2370
rect 5670 2360 6380 2370
rect 6740 2360 6900 2370
rect 7450 2360 7480 2370
rect 8410 2360 8420 2370
rect 9150 2360 9160 2370
rect 9250 2360 9260 2370
rect 9270 2360 9280 2370
rect 9320 2360 9330 2370
rect 9410 2360 9420 2370
rect 9460 2360 9470 2370
rect 9640 2360 9650 2370
rect 9830 2360 9840 2370
rect 1890 2350 1910 2360
rect 3260 2350 3280 2360
rect 5660 2350 6390 2360
rect 6740 2350 6840 2360
rect 6850 2350 6870 2360
rect 6880 2350 6920 2360
rect 7430 2350 7440 2360
rect 7460 2350 7480 2360
rect 8420 2350 8430 2360
rect 8510 2350 8530 2360
rect 9250 2350 9260 2360
rect 9300 2350 9310 2360
rect 9320 2350 9330 2360
rect 9360 2350 9380 2360
rect 9490 2350 9500 2360
rect 9550 2350 9570 2360
rect 9630 2350 9640 2360
rect 9800 2350 9810 2360
rect 9850 2350 9860 2360
rect 1890 2340 1900 2350
rect 3260 2340 3280 2350
rect 5670 2340 6390 2350
rect 6740 2340 6830 2350
rect 6900 2340 6940 2350
rect 7480 2340 7490 2350
rect 8430 2340 8540 2350
rect 9210 2340 9220 2350
rect 9240 2340 9260 2350
rect 9310 2340 9320 2350
rect 9330 2340 9340 2350
rect 9480 2340 9500 2350
rect 9540 2340 9550 2350
rect 9650 2340 9660 2350
rect 9720 2340 9730 2350
rect 9780 2340 9790 2350
rect 9800 2340 9810 2350
rect 1880 2330 1900 2340
rect 3260 2330 3290 2340
rect 5650 2330 6400 2340
rect 6740 2330 6830 2340
rect 6910 2330 6950 2340
rect 6960 2330 7010 2340
rect 7460 2330 7470 2340
rect 7490 2330 7500 2340
rect 8400 2330 8410 2340
rect 8460 2330 8470 2340
rect 8480 2330 8490 2340
rect 8500 2330 8560 2340
rect 9230 2330 9250 2340
rect 9330 2330 9340 2340
rect 9360 2330 9400 2340
rect 9440 2330 9450 2340
rect 9490 2330 9500 2340
rect 9550 2330 9560 2340
rect 9710 2330 9720 2340
rect 9800 2330 9810 2340
rect 9840 2330 9850 2340
rect 1880 2320 1900 2330
rect 3260 2320 3290 2330
rect 5480 2320 5520 2330
rect 5660 2320 6410 2330
rect 6730 2320 6840 2330
rect 6930 2320 7030 2330
rect 7470 2320 7480 2330
rect 7500 2320 7510 2330
rect 8520 2320 8570 2330
rect 9210 2320 9220 2330
rect 9370 2320 9390 2330
rect 9490 2320 9500 2330
rect 9830 2320 9840 2330
rect 1880 2310 1900 2320
rect 3260 2310 3290 2320
rect 5660 2310 6410 2320
rect 6740 2310 6750 2320
rect 6760 2310 6840 2320
rect 6950 2310 7060 2320
rect 7480 2310 7490 2320
rect 7510 2310 7540 2320
rect 8540 2310 8570 2320
rect 9360 2310 9380 2320
rect 9410 2310 9420 2320
rect 1880 2300 1900 2310
rect 3260 2300 3290 2310
rect 5480 2300 5510 2310
rect 5540 2300 5560 2310
rect 5660 2300 6420 2310
rect 6740 2300 6830 2310
rect 6950 2300 7050 2310
rect 7060 2300 7080 2310
rect 7180 2300 7200 2310
rect 7540 2300 7560 2310
rect 8560 2300 8580 2310
rect 9470 2300 9480 2310
rect 1880 2290 1890 2300
rect 3270 2290 3300 2300
rect 5480 2290 5500 2300
rect 5520 2290 5530 2300
rect 5640 2290 6410 2300
rect 6740 2290 6750 2300
rect 6760 2290 6830 2300
rect 6950 2290 7040 2300
rect 7070 2290 7220 2300
rect 7490 2290 7500 2300
rect 7560 2290 7580 2300
rect 8560 2290 8590 2300
rect 9620 2290 9630 2300
rect 9730 2290 9740 2300
rect 9820 2290 9830 2300
rect 1870 2280 1880 2290
rect 3270 2280 3300 2290
rect 5470 2280 5480 2290
rect 5520 2280 5530 2290
rect 5630 2280 5920 2290
rect 5940 2280 6000 2290
rect 6010 2280 6410 2290
rect 6420 2280 6430 2290
rect 6740 2280 6830 2290
rect 6960 2280 7040 2290
rect 7100 2280 7230 2290
rect 7570 2280 7590 2290
rect 8570 2280 8590 2290
rect 1870 2270 1880 2280
rect 3270 2270 3300 2280
rect 4150 2270 4210 2280
rect 4220 2270 4230 2280
rect 4240 2270 4250 2280
rect 5430 2270 5440 2280
rect 5460 2270 5490 2280
rect 5510 2270 5530 2280
rect 5650 2270 6000 2280
rect 6010 2270 6410 2280
rect 6740 2270 6820 2280
rect 6970 2270 7050 2280
rect 7170 2270 7260 2280
rect 7320 2270 7330 2280
rect 7500 2270 7510 2280
rect 7580 2270 7610 2280
rect 8580 2270 8600 2280
rect 9350 2270 9370 2280
rect 9790 2270 9800 2280
rect 1870 2260 1880 2270
rect 3270 2260 3300 2270
rect 5410 2260 5480 2270
rect 5510 2260 5520 2270
rect 5530 2260 5540 2270
rect 5640 2260 6400 2270
rect 6430 2260 6440 2270
rect 6740 2260 6760 2270
rect 6770 2260 6820 2270
rect 6990 2260 7070 2270
rect 7200 2260 7280 2270
rect 7320 2260 7330 2270
rect 7360 2260 7400 2270
rect 7590 2260 7620 2270
rect 8590 2260 8610 2270
rect 9130 2260 9150 2270
rect 9350 2260 9360 2270
rect 1860 2250 1870 2260
rect 3280 2250 3300 2260
rect 5420 2250 5530 2260
rect 5540 2250 5550 2260
rect 5640 2250 6400 2260
rect 6440 2250 6450 2260
rect 6740 2250 6750 2260
rect 6770 2250 6820 2260
rect 7000 2250 7040 2260
rect 7050 2250 7080 2260
rect 7240 2250 7250 2260
rect 7260 2250 7290 2260
rect 7320 2250 7330 2260
rect 7360 2250 7410 2260
rect 7510 2250 7520 2260
rect 7600 2250 7630 2260
rect 8610 2250 8640 2260
rect 9110 2250 9130 2260
rect 1860 2240 1870 2250
rect 3280 2240 3300 2250
rect 5420 2240 5430 2250
rect 5440 2240 5540 2250
rect 5590 2240 6400 2250
rect 6440 2240 6450 2250
rect 6740 2240 6760 2250
rect 6780 2240 6830 2250
rect 7020 2240 7040 2250
rect 7270 2240 7300 2250
rect 7310 2240 7390 2250
rect 7510 2240 7520 2250
rect 7610 2240 7630 2250
rect 8640 2240 8650 2250
rect 9080 2240 9100 2250
rect 9260 2240 9270 2250
rect 1860 2230 1870 2240
rect 3280 2230 3310 2240
rect 5410 2230 5540 2240
rect 5600 2230 6400 2240
rect 6740 2230 6760 2240
rect 6780 2230 6860 2240
rect 7280 2230 7380 2240
rect 7510 2230 7520 2240
rect 7620 2230 7640 2240
rect 8660 2230 8680 2240
rect 8720 2230 8730 2240
rect 8780 2230 8800 2240
rect 9060 2230 9070 2240
rect 9280 2230 9290 2240
rect 1860 2220 1870 2230
rect 3280 2220 3310 2230
rect 5400 2220 5460 2230
rect 5470 2220 5500 2230
rect 5520 2220 5530 2230
rect 5570 2220 5580 2230
rect 5590 2220 6400 2230
rect 6740 2220 6760 2230
rect 6790 2220 6880 2230
rect 7300 2220 7360 2230
rect 7370 2220 7380 2230
rect 7510 2220 7520 2230
rect 7640 2220 7650 2230
rect 8820 2220 8830 2230
rect 9030 2220 9050 2230
rect 9560 2220 9570 2230
rect 1860 2210 1870 2220
rect 2640 2210 2690 2220
rect 3280 2210 3300 2220
rect 5390 2210 5470 2220
rect 5490 2210 5510 2220
rect 5520 2210 5530 2220
rect 5580 2210 5600 2220
rect 5610 2210 6400 2220
rect 6740 2210 6760 2220
rect 6790 2210 6900 2220
rect 7330 2210 7340 2220
rect 7510 2210 7520 2220
rect 7650 2210 7660 2220
rect 8990 2210 9000 2220
rect 9550 2210 9560 2220
rect 9570 2210 9580 2220
rect 1860 2200 1870 2210
rect 2620 2200 2700 2210
rect 3280 2200 3300 2210
rect 5370 2200 5470 2210
rect 5500 2200 5510 2210
rect 5530 2200 5580 2210
rect 5590 2200 6400 2210
rect 6460 2200 6470 2210
rect 6750 2200 6780 2210
rect 6800 2200 6910 2210
rect 7380 2200 7390 2210
rect 7510 2200 7520 2210
rect 7660 2200 7680 2210
rect 8860 2200 8920 2210
rect 9700 2200 9710 2210
rect 9970 2200 9980 2210
rect 1860 2190 1870 2200
rect 2600 2190 2710 2200
rect 2720 2190 2750 2200
rect 3280 2190 3310 2200
rect 5360 2190 5470 2200
rect 5490 2190 5510 2200
rect 5520 2190 5530 2200
rect 5550 2190 6390 2200
rect 6750 2190 6770 2200
rect 6820 2190 6920 2200
rect 7380 2190 7390 2200
rect 7500 2190 7510 2200
rect 7680 2190 7690 2200
rect 9700 2190 9720 2200
rect 9810 2190 9820 2200
rect 9990 2190 9990 2200
rect 2450 2180 2490 2190
rect 2580 2180 2670 2190
rect 2760 2180 2770 2190
rect 2810 2180 2820 2190
rect 3280 2180 3300 2190
rect 5330 2180 5470 2190
rect 5490 2180 5520 2190
rect 5540 2180 6390 2190
rect 6750 2180 6770 2190
rect 6800 2180 6940 2190
rect 7490 2180 7510 2190
rect 7680 2180 7710 2190
rect 9730 2180 9740 2190
rect 9950 2180 9960 2190
rect 9980 2180 9990 2190
rect 1850 2170 1860 2180
rect 2430 2170 2440 2180
rect 2560 2170 2660 2180
rect 2760 2170 2840 2180
rect 3270 2170 3300 2180
rect 5320 2170 5480 2180
rect 5510 2170 6390 2180
rect 6750 2170 6770 2180
rect 6810 2170 6820 2180
rect 6830 2170 6960 2180
rect 7420 2170 7440 2180
rect 7470 2170 7510 2180
rect 7690 2170 7730 2180
rect 8360 2170 8370 2180
rect 9970 2170 9990 2180
rect 1850 2160 1860 2170
rect 2420 2160 2430 2170
rect 2550 2160 2640 2170
rect 2750 2160 2840 2170
rect 3270 2160 3300 2170
rect 5150 2160 5160 2170
rect 5310 2160 6390 2170
rect 6480 2160 6490 2170
rect 6750 2160 6770 2170
rect 6820 2160 6970 2170
rect 7390 2160 7400 2170
rect 7410 2160 7450 2170
rect 7460 2160 7500 2170
rect 7710 2160 7750 2170
rect 9790 2160 9800 2170
rect 1850 2150 1860 2160
rect 2400 2150 2420 2160
rect 2540 2150 2630 2160
rect 2740 2150 2830 2160
rect 3280 2150 3300 2160
rect 5310 2150 6390 2160
rect 6750 2150 6770 2160
rect 6820 2150 6950 2160
rect 7300 2150 7310 2160
rect 7390 2150 7420 2160
rect 7440 2150 7480 2160
rect 7730 2150 7750 2160
rect 9270 2150 9280 2160
rect 9590 2150 9600 2160
rect 9950 2150 9960 2160
rect 1850 2140 1860 2150
rect 2380 2140 2430 2150
rect 2540 2140 2630 2150
rect 2730 2140 2820 2150
rect 3280 2140 3300 2150
rect 5170 2140 5180 2150
rect 5290 2140 6380 2150
rect 6480 2140 6500 2150
rect 6760 2140 6790 2150
rect 6830 2140 6970 2150
rect 6990 2140 7000 2150
rect 7290 2140 7320 2150
rect 7400 2140 7420 2150
rect 7440 2140 7460 2150
rect 7740 2140 7840 2150
rect 8370 2140 8380 2150
rect 9590 2140 9600 2150
rect 9780 2140 9790 2150
rect 1840 2130 1860 2140
rect 2390 2130 2450 2140
rect 2540 2130 2640 2140
rect 2660 2130 2730 2140
rect 2760 2130 2800 2140
rect 3270 2130 3300 2140
rect 5170 2130 5180 2140
rect 5280 2130 6380 2140
rect 6480 2130 6500 2140
rect 6760 2130 6790 2140
rect 6850 2130 6860 2140
rect 6870 2130 6990 2140
rect 7290 2130 7310 2140
rect 7400 2130 7420 2140
rect 7800 2130 7820 2140
rect 7850 2130 7860 2140
rect 9230 2130 9240 2140
rect 9480 2130 9490 2140
rect 9670 2130 9680 2140
rect 1850 2120 1860 2130
rect 2410 2120 2660 2130
rect 3270 2120 3300 2130
rect 5270 2120 5400 2130
rect 5410 2120 6380 2130
rect 6470 2120 6510 2130
rect 6760 2120 6790 2130
rect 6870 2120 7000 2130
rect 7290 2120 7310 2130
rect 7410 2120 7430 2130
rect 7850 2120 7860 2130
rect 1840 2110 1870 2120
rect 2560 2110 2640 2120
rect 3260 2110 3300 2120
rect 5300 2110 6380 2120
rect 6480 2110 6510 2120
rect 6760 2110 6790 2120
rect 6870 2110 7020 2120
rect 7290 2110 7300 2120
rect 7850 2110 7860 2120
rect 9340 2110 9350 2120
rect 9520 2110 9530 2120
rect 9560 2110 9570 2120
rect 9670 2110 9700 2120
rect 1850 2100 1870 2110
rect 2570 2100 2630 2110
rect 3260 2100 3300 2110
rect 5250 2100 5260 2110
rect 5290 2100 6140 2110
rect 6150 2100 6380 2110
rect 6490 2100 6520 2110
rect 6760 2100 6780 2110
rect 6890 2100 7030 2110
rect 7280 2100 7300 2110
rect 7850 2100 7870 2110
rect 8390 2100 8400 2110
rect 9620 2100 9630 2110
rect 1850 2090 1870 2100
rect 2580 2090 2600 2100
rect 3260 2090 3300 2100
rect 5290 2090 6390 2100
rect 6490 2090 6520 2100
rect 6770 2090 6790 2100
rect 6860 2090 6870 2100
rect 6900 2090 7040 2100
rect 7270 2090 7310 2100
rect 8390 2090 8410 2100
rect 9250 2090 9260 2100
rect 9360 2090 9370 2100
rect 9530 2090 9540 2100
rect 1850 2080 1870 2090
rect 3260 2080 3300 2090
rect 5190 2080 5200 2090
rect 5280 2080 6380 2090
rect 6490 2080 6520 2090
rect 6770 2080 6790 2090
rect 6910 2080 7060 2090
rect 7260 2080 7300 2090
rect 7870 2080 7880 2090
rect 8390 2080 8420 2090
rect 9340 2080 9350 2090
rect 9460 2080 9470 2090
rect 9690 2080 9700 2090
rect 1850 2070 1870 2080
rect 3260 2070 3290 2080
rect 5260 2070 6150 2080
rect 6160 2070 6380 2080
rect 6490 2070 6510 2080
rect 6770 2070 6800 2080
rect 6920 2070 7050 2080
rect 7250 2070 7300 2080
rect 7870 2070 7890 2080
rect 8390 2070 8430 2080
rect 9260 2070 9270 2080
rect 9280 2070 9290 2080
rect 9370 2070 9380 2080
rect 9680 2070 9690 2080
rect 1850 2060 1860 2070
rect 3250 2060 3300 2070
rect 5110 2060 5130 2070
rect 5160 2060 5170 2070
rect 5260 2060 6390 2070
rect 6500 2060 6510 2070
rect 6770 2060 6800 2070
rect 6930 2060 7070 2070
rect 7220 2060 7300 2070
rect 7880 2060 7900 2070
rect 8390 2060 8440 2070
rect 9170 2060 9180 2070
rect 9200 2060 9210 2070
rect 9300 2060 9310 2070
rect 9570 2060 9580 2070
rect 9670 2060 9680 2070
rect 1840 2050 1860 2060
rect 3250 2050 3290 2060
rect 5060 2050 5070 2060
rect 5080 2050 5120 2060
rect 5130 2050 5140 2060
rect 5150 2050 5160 2060
rect 5240 2050 5250 2060
rect 5260 2050 6390 2060
rect 6490 2050 6510 2060
rect 6780 2050 6800 2060
rect 6950 2050 7100 2060
rect 7130 2050 7150 2060
rect 7170 2050 7210 2060
rect 7250 2050 7300 2060
rect 7320 2050 7330 2060
rect 7880 2050 7900 2060
rect 7960 2050 8000 2060
rect 8390 2050 8470 2060
rect 8480 2050 8500 2060
rect 9230 2050 9240 2060
rect 9600 2050 9630 2060
rect 9660 2050 9670 2060
rect 1840 2040 1860 2050
rect 3240 2040 3300 2050
rect 5110 2040 5150 2050
rect 5240 2040 6380 2050
rect 6480 2040 6510 2050
rect 6770 2040 6800 2050
rect 6970 2040 7160 2050
rect 7180 2040 7220 2050
rect 7230 2040 7300 2050
rect 7320 2040 7330 2050
rect 7890 2040 8010 2050
rect 8390 2040 8520 2050
rect 9140 2040 9150 2050
rect 9470 2040 9480 2050
rect 1850 2030 1860 2040
rect 3240 2030 3300 2040
rect 5120 2030 5150 2040
rect 5230 2030 5260 2040
rect 5270 2030 6380 2040
rect 6470 2030 6520 2040
rect 6780 2030 6810 2040
rect 6980 2030 7290 2040
rect 7320 2030 7330 2040
rect 7910 2030 7930 2040
rect 7960 2030 7980 2040
rect 8000 2030 8010 2040
rect 8390 2030 8470 2040
rect 8480 2030 8530 2040
rect 9120 2030 9140 2040
rect 1850 2020 1860 2030
rect 3230 2020 3300 2030
rect 5130 2020 5140 2030
rect 5150 2020 5170 2030
rect 5230 2020 5250 2030
rect 5260 2020 6370 2030
rect 6470 2020 6520 2030
rect 6780 2020 6820 2030
rect 6980 2020 7280 2030
rect 8390 2020 8440 2030
rect 8510 2020 8530 2030
rect 9090 2020 9110 2030
rect 9320 2020 9340 2030
rect 9370 2020 9390 2030
rect 1850 2010 1860 2020
rect 3230 2010 3310 2020
rect 5150 2010 5210 2020
rect 5230 2010 6360 2020
rect 6470 2010 6520 2020
rect 6780 2010 6820 2020
rect 7010 2010 7280 2020
rect 8390 2010 8440 2020
rect 8520 2010 8550 2020
rect 9180 2010 9210 2020
rect 9400 2010 9430 2020
rect 1850 2000 1870 2010
rect 3230 2000 3310 2010
rect 5160 2000 5210 2010
rect 5220 2000 6360 2010
rect 6480 2000 6520 2010
rect 6780 2000 6830 2010
rect 7020 2000 7280 2010
rect 7970 2000 7980 2010
rect 8390 2000 8440 2010
rect 8540 2000 8570 2010
rect 1850 1990 1860 2000
rect 3220 1990 3310 2000
rect 5010 1990 5030 2000
rect 5140 1990 5150 2000
rect 5160 1990 6160 2000
rect 6180 1990 6200 2000
rect 6210 1990 6230 2000
rect 6240 1990 6360 2000
rect 6480 1990 6520 2000
rect 6790 1990 6830 2000
rect 7040 1990 7280 2000
rect 7970 1990 7980 2000
rect 8380 1990 8450 2000
rect 8550 1990 8590 2000
rect 9680 1990 9690 2000
rect 1840 1980 1860 1990
rect 3220 1980 3310 1990
rect 4820 1980 4840 1990
rect 5060 1980 5140 1990
rect 5150 1980 6160 1990
rect 6180 1980 6190 1990
rect 6240 1980 6360 1990
rect 6480 1980 6520 1990
rect 6790 1980 6830 1990
rect 7050 1980 7280 1990
rect 7780 1980 7840 1990
rect 8380 1980 8450 1990
rect 8550 1980 8610 1990
rect 9660 1980 9670 1990
rect 1850 1970 1860 1980
rect 3220 1970 3320 1980
rect 4830 1970 4840 1980
rect 4850 1970 4870 1980
rect 4910 1970 4920 1980
rect 4930 1970 4940 1980
rect 5030 1970 6140 1980
rect 6150 1970 6220 1980
rect 6230 1970 6360 1980
rect 6460 1970 6530 1980
rect 6790 1970 6830 1980
rect 7070 1970 7280 1980
rect 7770 1970 7810 1980
rect 7840 1970 7850 1980
rect 8380 1970 8450 1980
rect 8570 1970 8680 1980
rect 9040 1970 9050 1980
rect 1840 1960 1860 1970
rect 3220 1960 3320 1970
rect 4860 1960 4880 1970
rect 4910 1960 4920 1970
rect 4990 1960 5000 1970
rect 5030 1960 6190 1970
rect 6200 1960 6210 1970
rect 6270 1960 6360 1970
rect 6470 1960 6530 1970
rect 6790 1960 6830 1970
rect 7090 1960 7270 1970
rect 7770 1960 7820 1970
rect 7970 1960 7980 1970
rect 8380 1960 8450 1970
rect 8590 1960 8710 1970
rect 8720 1960 8730 1970
rect 8860 1960 8880 1970
rect 9020 1960 9030 1970
rect 9930 1960 9960 1970
rect 1860 1950 1870 1960
rect 3220 1950 3320 1960
rect 5030 1950 6170 1960
rect 6190 1950 6200 1960
rect 6310 1950 6370 1960
rect 6470 1950 6540 1960
rect 6800 1950 6840 1960
rect 7140 1950 7160 1960
rect 7180 1950 7220 1960
rect 7780 1950 7830 1960
rect 7870 1950 7880 1960
rect 7960 1950 7970 1960
rect 8380 1950 8450 1960
rect 8640 1950 8660 1960
rect 8670 1950 8690 1960
rect 8710 1950 8760 1960
rect 8810 1950 8870 1960
rect 8890 1950 8990 1960
rect 9910 1950 9920 1960
rect 1850 1940 1860 1950
rect 3220 1940 3320 1950
rect 5020 1940 6170 1950
rect 6310 1940 6370 1950
rect 6480 1940 6520 1950
rect 6530 1940 6540 1950
rect 6790 1940 6830 1950
rect 7140 1940 7150 1950
rect 7780 1940 7840 1950
rect 7890 1940 7900 1950
rect 7940 1940 7950 1950
rect 8380 1940 8450 1950
rect 8770 1940 8810 1950
rect 9670 1940 9680 1950
rect 9880 1940 9890 1950
rect 9900 1940 9910 1950
rect 1850 1930 1860 1940
rect 3220 1930 3320 1940
rect 4540 1930 4550 1940
rect 4600 1930 4620 1940
rect 4780 1930 4790 1940
rect 4840 1930 4860 1940
rect 4980 1930 6170 1940
rect 6340 1930 6380 1940
rect 6480 1930 6520 1940
rect 6800 1930 6830 1940
rect 7330 1930 7340 1940
rect 7780 1930 7840 1940
rect 8380 1930 8450 1940
rect 9680 1930 9690 1940
rect 9980 1930 9990 1940
rect 1850 1920 1860 1930
rect 3230 1920 3320 1930
rect 4490 1920 4500 1930
rect 4630 1920 4640 1930
rect 4860 1920 4870 1930
rect 4980 1920 6180 1930
rect 6340 1920 6380 1930
rect 6490 1920 6520 1930
rect 6800 1920 6830 1930
rect 7330 1920 7340 1930
rect 7770 1920 7830 1930
rect 8380 1920 8450 1930
rect 9600 1920 9680 1930
rect 9870 1920 9880 1930
rect 9960 1920 9970 1930
rect 1850 1910 1860 1920
rect 2660 1910 2690 1920
rect 3250 1910 3320 1920
rect 4480 1910 4490 1920
rect 4550 1910 4570 1920
rect 4640 1910 4650 1920
rect 4770 1910 4780 1920
rect 4810 1910 4880 1920
rect 4970 1910 4980 1920
rect 5000 1910 5020 1920
rect 5060 1910 6180 1920
rect 6340 1910 6390 1920
rect 6470 1910 6530 1920
rect 6800 1910 6840 1920
rect 7330 1910 7340 1920
rect 7790 1910 7840 1920
rect 8380 1910 8450 1920
rect 9610 1910 9630 1920
rect 9670 1910 9690 1920
rect 1850 1900 1860 1910
rect 2600 1900 2660 1910
rect 2680 1900 2730 1910
rect 3270 1900 3320 1910
rect 4640 1900 4650 1910
rect 4770 1900 4780 1910
rect 4850 1900 4860 1910
rect 5000 1900 5010 1910
rect 5020 1900 5030 1910
rect 5110 1900 6150 1910
rect 6160 1900 6180 1910
rect 6340 1900 6540 1910
rect 6800 1900 6830 1910
rect 7780 1900 7850 1910
rect 8380 1900 8450 1910
rect 9600 1900 9610 1910
rect 9680 1900 9690 1910
rect 1850 1890 1860 1900
rect 2460 1890 2550 1900
rect 2560 1890 2570 1900
rect 2700 1890 2740 1900
rect 3270 1890 3320 1900
rect 4370 1890 4380 1900
rect 4810 1890 4820 1900
rect 4880 1890 4890 1900
rect 4960 1890 4970 1900
rect 5020 1890 5030 1900
rect 5050 1890 5060 1900
rect 5140 1890 6150 1900
rect 6160 1890 6180 1900
rect 6340 1890 6550 1900
rect 6790 1890 6830 1900
rect 7790 1890 7850 1900
rect 8370 1890 8450 1900
rect 9930 1890 9960 1900
rect 9970 1890 9980 1900
rect 1850 1880 1870 1890
rect 2450 1880 2480 1890
rect 2720 1880 2780 1890
rect 2800 1880 2820 1890
rect 3270 1880 3320 1890
rect 4340 1880 4350 1890
rect 4360 1880 4370 1890
rect 4760 1880 4770 1890
rect 4790 1880 4800 1890
rect 4810 1880 4820 1890
rect 4880 1880 4900 1890
rect 4910 1880 4920 1890
rect 4950 1880 4980 1890
rect 5010 1880 5020 1890
rect 5040 1880 5110 1890
rect 5140 1880 6150 1890
rect 6160 1880 6180 1890
rect 6350 1880 6480 1890
rect 6490 1880 6500 1890
rect 6540 1880 6560 1890
rect 6800 1880 6830 1890
rect 7780 1880 7850 1890
rect 8370 1880 8450 1890
rect 9760 1880 9770 1890
rect 2430 1870 2470 1880
rect 2750 1870 2830 1880
rect 3270 1870 3320 1880
rect 4320 1870 4330 1880
rect 4340 1870 4350 1880
rect 4400 1870 4410 1880
rect 4470 1870 4480 1880
rect 4560 1870 4570 1880
rect 4590 1870 4600 1880
rect 4760 1870 4770 1880
rect 4800 1870 4810 1880
rect 4880 1870 4900 1880
rect 4910 1870 4930 1880
rect 4960 1870 4990 1880
rect 5030 1870 5090 1880
rect 5100 1870 5110 1880
rect 5140 1870 6170 1880
rect 6350 1870 6460 1880
rect 6550 1870 6570 1880
rect 6800 1870 6830 1880
rect 7790 1870 7850 1880
rect 8370 1870 8450 1880
rect 9150 1870 9160 1880
rect 9190 1870 9200 1880
rect 9240 1870 9250 1880
rect 9530 1870 9540 1880
rect 1860 1860 1870 1870
rect 2400 1860 2440 1870
rect 2800 1860 2840 1870
rect 3260 1860 3270 1870
rect 3280 1860 3310 1870
rect 4290 1860 4300 1870
rect 4470 1860 4480 1870
rect 4780 1860 4790 1870
rect 4800 1860 4810 1870
rect 4880 1860 4900 1870
rect 4910 1860 4920 1870
rect 4950 1860 5000 1870
rect 5040 1860 5090 1870
rect 5150 1860 5200 1870
rect 5210 1860 5230 1870
rect 5270 1860 6140 1870
rect 6170 1860 6180 1870
rect 6350 1860 6460 1870
rect 6560 1860 6570 1870
rect 6800 1860 6840 1870
rect 7790 1860 7850 1870
rect 8370 1860 8450 1870
rect 9200 1860 9210 1870
rect 9250 1860 9270 1870
rect 9280 1860 9300 1870
rect 9310 1860 9320 1870
rect 9360 1860 9380 1870
rect 1850 1850 1870 1860
rect 2390 1850 2420 1860
rect 2530 1850 2560 1860
rect 2830 1850 2860 1860
rect 2870 1850 2890 1860
rect 3280 1850 3310 1860
rect 4300 1850 4310 1860
rect 4470 1850 4480 1860
rect 4530 1850 4540 1860
rect 4580 1850 4590 1860
rect 4600 1850 4610 1860
rect 4750 1850 4760 1860
rect 4890 1850 4920 1860
rect 4950 1850 5020 1860
rect 5050 1850 5090 1860
rect 5130 1850 5140 1860
rect 5150 1850 5180 1860
rect 5220 1850 5230 1860
rect 5300 1850 6130 1860
rect 6290 1850 6320 1860
rect 6330 1850 6450 1860
rect 6800 1850 6840 1860
rect 7790 1850 7850 1860
rect 8370 1850 8380 1860
rect 8390 1850 8450 1860
rect 9200 1850 9210 1860
rect 9770 1850 9780 1860
rect 1860 1840 1880 1850
rect 2370 1840 2390 1850
rect 2520 1840 2580 1850
rect 2850 1840 2890 1850
rect 3280 1840 3310 1850
rect 4340 1840 4350 1850
rect 4360 1840 4370 1850
rect 4530 1840 4540 1850
rect 4580 1840 4590 1850
rect 4600 1840 4610 1850
rect 4750 1840 4760 1850
rect 4790 1840 4810 1850
rect 4900 1840 4930 1850
rect 4940 1840 5010 1850
rect 5040 1840 5080 1850
rect 5150 1840 5170 1850
rect 5210 1840 5260 1850
rect 5310 1840 6110 1850
rect 6280 1840 6460 1850
rect 6810 1840 6830 1850
rect 7790 1840 7860 1850
rect 8380 1840 8400 1850
rect 8410 1840 8450 1850
rect 9110 1840 9120 1850
rect 9190 1840 9200 1850
rect 9210 1840 9230 1850
rect 9330 1840 9340 1850
rect 1850 1830 1870 1840
rect 2350 1830 2380 1840
rect 2530 1830 2550 1840
rect 2880 1830 2900 1840
rect 3270 1830 3310 1840
rect 4280 1830 4290 1840
rect 4330 1830 4350 1840
rect 4530 1830 4540 1840
rect 4740 1830 4750 1840
rect 4770 1830 4780 1840
rect 4790 1830 4810 1840
rect 4850 1830 4860 1840
rect 4870 1830 4880 1840
rect 4890 1830 4930 1840
rect 4940 1830 5010 1840
rect 5030 1830 5070 1840
rect 5110 1830 5120 1840
rect 5140 1830 5170 1840
rect 5200 1830 5260 1840
rect 5270 1830 5290 1840
rect 5320 1830 6080 1840
rect 6270 1830 6460 1840
rect 6810 1830 6840 1840
rect 7790 1830 7860 1840
rect 8360 1830 8370 1840
rect 8380 1830 8400 1840
rect 8410 1830 8450 1840
rect 9180 1830 9200 1840
rect 9220 1830 9230 1840
rect 9380 1830 9400 1840
rect 1850 1820 1870 1830
rect 2320 1820 2350 1830
rect 2880 1820 2910 1830
rect 3270 1820 3310 1830
rect 4270 1820 4280 1830
rect 4330 1820 4340 1830
rect 4470 1820 4480 1830
rect 4530 1820 4540 1830
rect 4740 1820 4750 1830
rect 4790 1820 4810 1830
rect 4850 1820 4860 1830
rect 4880 1820 4900 1830
rect 4910 1820 5010 1830
rect 5030 1820 5060 1830
rect 5100 1820 5160 1830
rect 5200 1820 5300 1830
rect 5330 1820 6080 1830
rect 6280 1820 6400 1830
rect 6410 1820 6470 1830
rect 6800 1820 6840 1830
rect 7780 1820 7850 1830
rect 8360 1820 8450 1830
rect 9310 1820 9330 1830
rect 1860 1810 1880 1820
rect 2290 1810 2330 1820
rect 2840 1810 2900 1820
rect 3270 1810 3300 1820
rect 4270 1810 4280 1820
rect 4330 1810 4340 1820
rect 4530 1810 4540 1820
rect 4740 1810 4750 1820
rect 4790 1810 4800 1820
rect 4840 1810 4850 1820
rect 4890 1810 4900 1820
rect 4910 1810 4970 1820
rect 5040 1810 5060 1820
rect 5090 1810 5160 1820
rect 5180 1810 5190 1820
rect 5200 1810 5300 1820
rect 5330 1810 6080 1820
rect 6280 1810 6380 1820
rect 6410 1810 6500 1820
rect 6800 1810 6840 1820
rect 7790 1810 7860 1820
rect 8360 1810 8370 1820
rect 8390 1810 8460 1820
rect 9250 1810 9270 1820
rect 9290 1810 9300 1820
rect 9380 1810 9390 1820
rect 9430 1810 9440 1820
rect 9980 1810 9990 1820
rect 1850 1800 1890 1810
rect 2250 1800 2310 1810
rect 2800 1800 2810 1810
rect 3270 1800 3300 1810
rect 4330 1800 4340 1810
rect 4760 1800 4770 1810
rect 4780 1800 4790 1810
rect 4830 1800 4840 1810
rect 4850 1800 4860 1810
rect 4890 1800 4900 1810
rect 4910 1800 4920 1810
rect 4930 1800 4980 1810
rect 5040 1800 5050 1810
rect 5090 1800 5150 1810
rect 5190 1800 5230 1810
rect 5250 1800 5260 1810
rect 5270 1800 5320 1810
rect 5340 1800 6070 1810
rect 6280 1800 6370 1810
rect 6420 1800 6510 1810
rect 6800 1800 6840 1810
rect 7340 1800 7350 1810
rect 7790 1800 7860 1810
rect 8360 1800 8370 1810
rect 8380 1800 8390 1810
rect 8400 1800 8460 1810
rect 9200 1800 9210 1810
rect 9270 1800 9280 1810
rect 9370 1800 9380 1810
rect 1860 1790 1880 1800
rect 2240 1790 2300 1800
rect 2460 1790 2520 1800
rect 2710 1790 2780 1800
rect 3260 1790 3300 1800
rect 4110 1790 4120 1800
rect 4330 1790 4340 1800
rect 4560 1790 4570 1800
rect 4610 1790 4620 1800
rect 4730 1790 4740 1800
rect 4780 1790 4790 1800
rect 4830 1790 4840 1800
rect 4850 1790 4860 1800
rect 4890 1790 4950 1800
rect 4980 1790 5000 1800
rect 5020 1790 5050 1800
rect 5070 1790 5150 1800
rect 5170 1790 5220 1800
rect 5280 1790 5320 1800
rect 5340 1790 6040 1800
rect 6050 1790 6070 1800
rect 6290 1790 6370 1800
rect 6420 1790 6520 1800
rect 6810 1790 6840 1800
rect 7340 1790 7350 1800
rect 7790 1790 7850 1800
rect 8360 1790 8370 1800
rect 8400 1790 8460 1800
rect 9420 1790 9430 1800
rect 9450 1790 9460 1800
rect 9770 1790 9780 1800
rect 9920 1790 9930 1800
rect 9940 1790 9950 1800
rect 1870 1780 1880 1790
rect 2260 1780 2340 1790
rect 2420 1780 2760 1790
rect 3260 1780 3290 1790
rect 4330 1780 4350 1790
rect 4610 1780 4620 1790
rect 4810 1780 4820 1790
rect 4840 1780 4860 1790
rect 4890 1780 4990 1790
rect 5020 1780 5050 1790
rect 5080 1780 5140 1790
rect 5180 1780 5220 1790
rect 5240 1780 5260 1790
rect 5280 1780 5320 1790
rect 5340 1780 6050 1790
rect 6290 1780 6370 1790
rect 6420 1780 6550 1790
rect 6810 1780 6840 1790
rect 7340 1780 7350 1790
rect 7800 1780 7860 1790
rect 8400 1780 8470 1790
rect 9100 1780 9110 1790
rect 9770 1780 9780 1790
rect 9930 1780 9940 1790
rect 1870 1770 1880 1780
rect 2360 1770 2370 1780
rect 2380 1770 2630 1780
rect 2650 1770 2660 1780
rect 3260 1770 3290 1780
rect 4290 1770 4300 1780
rect 4330 1770 4340 1780
rect 4400 1770 4410 1780
rect 4720 1770 4730 1780
rect 4750 1770 4780 1780
rect 4810 1770 4820 1780
rect 4850 1770 4860 1780
rect 4880 1770 4990 1780
rect 5030 1770 5050 1780
rect 5070 1770 5140 1780
rect 5160 1770 5170 1780
rect 5180 1770 5210 1780
rect 5240 1770 5260 1780
rect 5280 1770 5310 1780
rect 5350 1770 5410 1780
rect 5460 1770 6050 1780
rect 6300 1770 6370 1780
rect 6420 1770 6550 1780
rect 6810 1770 6850 1780
rect 7810 1770 7860 1780
rect 8400 1770 8480 1780
rect 9100 1770 9110 1780
rect 9910 1770 9920 1780
rect 1880 1760 1890 1770
rect 2400 1760 2530 1770
rect 3250 1760 3290 1770
rect 4210 1760 4220 1770
rect 4290 1760 4300 1770
rect 4610 1760 4620 1770
rect 4630 1760 4640 1770
rect 4690 1760 4710 1770
rect 4720 1760 4730 1770
rect 4760 1760 4780 1770
rect 4790 1760 4800 1770
rect 4810 1760 4830 1770
rect 4880 1760 4950 1770
rect 4960 1760 4990 1770
rect 5010 1760 5040 1770
rect 5060 1760 5130 1770
rect 5160 1760 5200 1770
rect 5240 1760 5250 1770
rect 5280 1760 5310 1770
rect 5330 1760 5340 1770
rect 5360 1760 5400 1770
rect 5470 1760 6040 1770
rect 6310 1760 6360 1770
rect 6410 1760 6550 1770
rect 6810 1760 6840 1770
rect 7810 1760 7860 1770
rect 8350 1760 8360 1770
rect 8370 1760 8490 1770
rect 8500 1760 8520 1770
rect 9370 1760 9380 1770
rect 9410 1760 9420 1770
rect 1880 1750 1890 1760
rect 2430 1750 2530 1760
rect 3260 1750 3280 1760
rect 4070 1750 4080 1760
rect 4700 1750 4720 1760
rect 4760 1750 4820 1760
rect 4840 1750 4860 1760
rect 4880 1750 4920 1760
rect 4930 1750 4950 1760
rect 4960 1750 4990 1760
rect 5010 1750 5040 1760
rect 5070 1750 5130 1760
rect 5170 1750 5200 1760
rect 5230 1750 5250 1760
rect 5280 1750 5300 1760
rect 5360 1750 5400 1760
rect 5430 1750 5450 1760
rect 5490 1750 6050 1760
rect 6320 1750 6370 1760
rect 6410 1750 6550 1760
rect 6810 1750 6840 1760
rect 7800 1750 7860 1760
rect 8350 1750 8360 1760
rect 8390 1750 8490 1760
rect 9200 1750 9210 1760
rect 9420 1750 9430 1760
rect 9830 1750 9850 1760
rect 1880 1740 1900 1750
rect 2440 1740 2500 1750
rect 3250 1740 3280 1750
rect 4220 1740 4230 1750
rect 4530 1740 4540 1750
rect 4640 1740 4650 1750
rect 4710 1740 4720 1750
rect 4740 1740 4750 1750
rect 4760 1740 4770 1750
rect 4780 1740 4860 1750
rect 4890 1740 4940 1750
rect 4960 1740 4980 1750
rect 5010 1740 5040 1750
rect 5070 1740 5130 1750
rect 5160 1740 5190 1750
rect 5220 1740 5250 1750
rect 5270 1740 5300 1750
rect 5320 1740 5330 1750
rect 5340 1740 5380 1750
rect 5420 1740 5430 1750
rect 5440 1740 5470 1750
rect 5510 1740 6030 1750
rect 6310 1740 6370 1750
rect 6410 1740 6550 1750
rect 6810 1740 6840 1750
rect 7810 1740 7860 1750
rect 8350 1740 8360 1750
rect 8390 1740 8500 1750
rect 9200 1740 9210 1750
rect 1880 1730 1900 1740
rect 3240 1730 3280 1740
rect 4350 1730 4360 1740
rect 4380 1730 4390 1740
rect 4530 1730 4540 1740
rect 4620 1730 4630 1740
rect 4700 1730 4710 1740
rect 4750 1730 4800 1740
rect 4830 1730 4870 1740
rect 4890 1730 4950 1740
rect 4960 1730 4980 1740
rect 5010 1730 5030 1740
rect 5050 1730 5060 1740
rect 5070 1730 5120 1740
rect 5150 1730 5190 1740
rect 5220 1730 5240 1740
rect 5270 1730 5290 1740
rect 5350 1730 5380 1740
rect 5410 1730 5420 1740
rect 5430 1730 5480 1740
rect 5520 1730 6030 1740
rect 6310 1730 6380 1740
rect 6390 1730 6510 1740
rect 6530 1730 6550 1740
rect 6810 1730 6840 1740
rect 7800 1730 7860 1740
rect 8350 1730 8370 1740
rect 8390 1730 8510 1740
rect 9540 1730 9550 1740
rect 9830 1730 9840 1740
rect 9930 1730 9940 1740
rect 1890 1720 1900 1730
rect 3240 1720 3280 1730
rect 4350 1720 4360 1730
rect 4530 1720 4540 1730
rect 4550 1720 4570 1730
rect 4580 1720 4590 1730
rect 4650 1720 4660 1730
rect 4700 1720 4710 1730
rect 4730 1720 4740 1730
rect 4760 1720 4770 1730
rect 4820 1720 4830 1730
rect 4840 1720 4870 1730
rect 4890 1720 4950 1730
rect 4970 1720 4980 1730
rect 5000 1720 5030 1730
rect 5060 1720 5120 1730
rect 5140 1720 5180 1730
rect 5210 1720 5240 1730
rect 5270 1720 5290 1730
rect 5330 1720 5370 1730
rect 5410 1720 5490 1730
rect 5530 1720 5990 1730
rect 6000 1720 6030 1730
rect 6320 1720 6490 1730
rect 6510 1720 6540 1730
rect 6810 1720 6840 1730
rect 7810 1720 7860 1730
rect 8350 1720 8370 1730
rect 8390 1720 8500 1730
rect 1900 1710 1910 1720
rect 3240 1710 3270 1720
rect 3480 1710 3490 1720
rect 4230 1710 4240 1720
rect 4300 1710 4310 1720
rect 4530 1710 4540 1720
rect 4630 1710 4640 1720
rect 4650 1710 4660 1720
rect 4700 1710 4710 1720
rect 4830 1710 4870 1720
rect 4890 1710 4920 1720
rect 4930 1710 4970 1720
rect 5010 1710 5030 1720
rect 5040 1710 5050 1720
rect 5060 1710 5110 1720
rect 5140 1710 5180 1720
rect 5200 1710 5230 1720
rect 5270 1710 5280 1720
rect 5320 1710 5370 1720
rect 5400 1710 5510 1720
rect 5540 1710 5990 1720
rect 6020 1710 6050 1720
rect 6320 1710 6490 1720
rect 6500 1710 6540 1720
rect 6810 1710 6850 1720
rect 7810 1710 7860 1720
rect 8340 1710 8370 1720
rect 8390 1710 8500 1720
rect 9920 1710 9930 1720
rect 1890 1700 1920 1710
rect 2580 1700 2600 1710
rect 3230 1700 3260 1710
rect 4300 1700 4310 1710
rect 4530 1700 4540 1710
rect 4590 1700 4600 1710
rect 4750 1700 4760 1710
rect 4830 1700 4870 1710
rect 4890 1700 4970 1710
rect 4990 1700 5030 1710
rect 5050 1700 5110 1710
rect 5140 1700 5170 1710
rect 5200 1700 5220 1710
rect 5250 1700 5280 1710
rect 5330 1700 5360 1710
rect 5390 1700 5430 1710
rect 5450 1700 5460 1710
rect 5470 1700 5520 1710
rect 5540 1700 6010 1710
rect 6330 1700 6540 1710
rect 6810 1700 6840 1710
rect 7350 1700 7360 1710
rect 7820 1700 7860 1710
rect 8340 1700 8360 1710
rect 8380 1700 8510 1710
rect 9210 1700 9220 1710
rect 9920 1700 9930 1710
rect 1900 1690 1920 1700
rect 2570 1690 2600 1700
rect 3220 1690 3260 1700
rect 4240 1690 4250 1700
rect 4290 1690 4310 1700
rect 4530 1690 4540 1700
rect 4660 1690 4670 1700
rect 4690 1690 4700 1700
rect 4720 1690 4730 1700
rect 4770 1690 4780 1700
rect 4850 1690 4870 1700
rect 4900 1690 4960 1700
rect 5000 1690 5030 1700
rect 5050 1690 5110 1700
rect 5130 1690 5170 1700
rect 5190 1690 5220 1700
rect 5260 1690 5270 1700
rect 5310 1690 5350 1700
rect 5390 1690 5420 1700
rect 5480 1690 5520 1700
rect 5550 1690 6000 1700
rect 6330 1690 6530 1700
rect 6810 1690 6850 1700
rect 7340 1690 7360 1700
rect 7810 1690 7870 1700
rect 8340 1690 8360 1700
rect 8390 1690 8510 1700
rect 9110 1690 9120 1700
rect 9200 1690 9230 1700
rect 1900 1680 1920 1690
rect 2540 1680 2550 1690
rect 2560 1680 2590 1690
rect 3220 1680 3260 1690
rect 4070 1680 4080 1690
rect 4420 1680 4440 1690
rect 4580 1680 4590 1690
rect 4640 1680 4650 1690
rect 4690 1680 4700 1690
rect 4790 1680 4820 1690
rect 4830 1680 4840 1690
rect 4850 1680 4870 1690
rect 4900 1680 4960 1690
rect 4990 1680 5030 1690
rect 5050 1680 5100 1690
rect 5120 1680 5160 1690
rect 5190 1680 5210 1690
rect 5240 1680 5270 1690
rect 5310 1680 5340 1690
rect 5380 1680 5410 1690
rect 5440 1680 5450 1690
rect 5490 1680 5530 1690
rect 5550 1680 5980 1690
rect 6000 1680 6020 1690
rect 6330 1680 6480 1690
rect 6490 1680 6520 1690
rect 6810 1680 6850 1690
rect 7340 1680 7360 1690
rect 7810 1680 7870 1690
rect 8340 1680 8360 1690
rect 8390 1680 8510 1690
rect 9210 1680 9220 1690
rect 9790 1680 9800 1690
rect 9910 1680 9920 1690
rect 1900 1670 1930 1680
rect 2570 1670 2580 1680
rect 2590 1670 2600 1680
rect 3210 1670 3250 1680
rect 4170 1670 4180 1680
rect 4250 1670 4260 1680
rect 4380 1670 4390 1680
rect 4740 1670 4750 1680
rect 4790 1670 4840 1680
rect 4890 1670 4960 1680
rect 4980 1670 5010 1680
rect 5040 1670 5100 1680
rect 5120 1670 5160 1680
rect 5180 1670 5210 1680
rect 5250 1670 5260 1680
rect 5310 1670 5340 1680
rect 5380 1670 5410 1680
rect 5450 1670 5460 1680
rect 5490 1670 5530 1680
rect 5560 1670 6010 1680
rect 6020 1670 6040 1680
rect 6330 1670 6510 1680
rect 6810 1670 6840 1680
rect 7350 1670 7360 1680
rect 7810 1670 7870 1680
rect 8390 1670 8510 1680
rect 9910 1670 9920 1680
rect 1910 1660 1930 1670
rect 3210 1660 3240 1670
rect 4160 1660 4170 1670
rect 4350 1660 4370 1670
rect 4400 1660 4410 1670
rect 4430 1660 4440 1670
rect 4450 1660 4460 1670
rect 4590 1660 4600 1670
rect 4630 1660 4640 1670
rect 4790 1660 4830 1670
rect 4900 1660 4910 1670
rect 4930 1660 4960 1670
rect 4980 1660 5010 1670
rect 5040 1660 5100 1670
rect 5120 1660 5160 1670
rect 5180 1660 5200 1670
rect 5230 1660 5260 1670
rect 5300 1660 5330 1670
rect 5360 1660 5400 1670
rect 5450 1660 5460 1670
rect 5490 1660 5530 1670
rect 5560 1660 5960 1670
rect 5970 1660 5980 1670
rect 5990 1660 6010 1670
rect 6030 1660 6040 1670
rect 6330 1660 6500 1670
rect 6810 1660 6840 1670
rect 7350 1660 7360 1670
rect 7810 1660 7870 1670
rect 8330 1660 8340 1670
rect 8390 1660 8520 1670
rect 9710 1660 9720 1670
rect 9780 1660 9790 1670
rect 9900 1660 9910 1670
rect 1910 1650 1940 1660
rect 3200 1650 3240 1660
rect 4080 1650 4100 1660
rect 4130 1650 4190 1660
rect 4260 1650 4270 1660
rect 4370 1650 4380 1660
rect 4510 1650 4520 1660
rect 4600 1650 4610 1660
rect 4660 1650 4670 1660
rect 4690 1650 4710 1660
rect 4750 1650 4760 1660
rect 4780 1650 4830 1660
rect 4940 1650 4960 1660
rect 4990 1650 5010 1660
rect 5040 1650 5100 1660
rect 5110 1650 5160 1660
rect 5170 1650 5190 1660
rect 5220 1650 5230 1660
rect 5240 1650 5250 1660
rect 5290 1650 5300 1660
rect 5350 1650 5400 1660
rect 5440 1650 5460 1660
rect 5490 1650 5530 1660
rect 5550 1650 5980 1660
rect 6000 1650 6010 1660
rect 6340 1650 6500 1660
rect 6820 1650 6840 1660
rect 7350 1650 7360 1660
rect 7810 1650 7870 1660
rect 8330 1650 8340 1660
rect 8400 1650 8510 1660
rect 9200 1650 9210 1660
rect 9870 1650 9880 1660
rect 9890 1650 9900 1660
rect 9960 1650 9970 1660
rect 1920 1640 1940 1650
rect 3200 1640 3240 1650
rect 4100 1640 4200 1650
rect 4430 1640 4440 1650
rect 4680 1640 4710 1650
rect 4770 1640 4800 1650
rect 4810 1640 4860 1650
rect 4870 1640 4880 1650
rect 4900 1640 4920 1650
rect 4930 1640 4960 1650
rect 4980 1640 5000 1650
rect 5040 1640 5100 1650
rect 5110 1640 5170 1650
rect 5220 1640 5230 1650
rect 5240 1640 5250 1650
rect 5290 1640 5300 1650
rect 5340 1640 5400 1650
rect 5490 1640 5520 1650
rect 5550 1640 5560 1650
rect 5570 1640 5940 1650
rect 5960 1640 5980 1650
rect 6340 1640 6490 1650
rect 6500 1640 6510 1650
rect 6810 1640 6830 1650
rect 7350 1640 7360 1650
rect 7820 1640 7870 1650
rect 8330 1640 8340 1650
rect 8370 1640 8430 1650
rect 8450 1640 8480 1650
rect 8490 1640 8500 1650
rect 1920 1630 1940 1640
rect 3190 1630 3230 1640
rect 4090 1630 4210 1640
rect 4700 1630 4730 1640
rect 4760 1630 4780 1640
rect 4810 1630 4840 1640
rect 4900 1630 4960 1640
rect 5030 1630 5100 1640
rect 5120 1630 5170 1640
rect 5230 1630 5240 1640
rect 5290 1630 5300 1640
rect 5330 1630 5410 1640
rect 5480 1630 5520 1640
rect 5550 1630 5560 1640
rect 5570 1630 5950 1640
rect 5960 1630 6000 1640
rect 6340 1630 6500 1640
rect 6820 1630 6840 1640
rect 7350 1630 7360 1640
rect 7820 1630 7870 1640
rect 8370 1630 8430 1640
rect 8450 1630 8470 1640
rect 9820 1630 9840 1640
rect 9880 1630 9890 1640
rect 9950 1630 9960 1640
rect 1920 1620 1950 1630
rect 3190 1620 3220 1630
rect 4090 1620 4210 1630
rect 4310 1620 4320 1630
rect 4360 1620 4370 1630
rect 4380 1620 4390 1630
rect 4660 1620 4670 1630
rect 4720 1620 4760 1630
rect 4800 1620 4970 1630
rect 4990 1620 5010 1630
rect 5030 1620 5100 1630
rect 5130 1620 5190 1630
rect 5210 1620 5240 1630
rect 5280 1620 5290 1630
rect 5330 1620 5420 1630
rect 5470 1620 5510 1630
rect 5550 1620 5560 1630
rect 5570 1620 5620 1630
rect 5640 1620 5990 1630
rect 6330 1620 6490 1630
rect 6810 1620 6840 1630
rect 7820 1620 7880 1630
rect 8380 1620 8430 1630
rect 9250 1620 9260 1630
rect 9720 1620 9730 1630
rect 9820 1620 9840 1630
rect 9850 1620 9860 1630
rect 1930 1610 1950 1620
rect 3170 1610 3220 1620
rect 4100 1610 4220 1620
rect 4310 1610 4320 1620
rect 4390 1610 4400 1620
rect 4720 1610 4750 1620
rect 4800 1610 4810 1620
rect 4820 1610 4980 1620
rect 5030 1610 5110 1620
rect 5140 1610 5230 1620
rect 5320 1610 5430 1620
rect 5440 1610 5500 1620
rect 5540 1610 5600 1620
rect 5660 1610 5970 1620
rect 6330 1610 6480 1620
rect 6810 1610 6830 1620
rect 7350 1610 7360 1620
rect 7820 1610 7880 1620
rect 8320 1610 8350 1620
rect 8390 1610 8430 1620
rect 9210 1610 9220 1620
rect 9230 1610 9240 1620
rect 9380 1610 9420 1620
rect 9710 1610 9740 1620
rect 9870 1610 9880 1620
rect 1930 1600 1960 1610
rect 3170 1600 3210 1610
rect 4100 1600 4220 1610
rect 4280 1600 4290 1610
rect 4310 1600 4320 1610
rect 4810 1600 5120 1610
rect 5140 1600 5170 1610
rect 5190 1600 5210 1610
rect 5270 1600 5280 1610
rect 5310 1600 5360 1610
rect 5410 1600 5480 1610
rect 5520 1600 5530 1610
rect 5550 1600 5580 1610
rect 5680 1600 5970 1610
rect 6330 1600 6440 1610
rect 6820 1600 6840 1610
rect 7830 1600 7880 1610
rect 8320 1600 8330 1610
rect 8380 1600 8440 1610
rect 9160 1600 9170 1610
rect 9380 1600 9420 1610
rect 1930 1590 1970 1600
rect 3160 1590 3200 1600
rect 4100 1590 4220 1600
rect 4290 1590 4310 1600
rect 4900 1590 5130 1600
rect 5150 1590 5160 1600
rect 5260 1590 5270 1600
rect 5300 1590 5350 1600
rect 5420 1590 5460 1600
rect 5530 1590 5580 1600
rect 5620 1590 5640 1600
rect 5690 1590 5960 1600
rect 6340 1590 6440 1600
rect 6810 1590 6830 1600
rect 7820 1590 7880 1600
rect 8320 1590 8330 1600
rect 8390 1590 8450 1600
rect 9830 1590 9840 1600
rect 1940 1580 1970 1590
rect 3150 1580 3200 1590
rect 4110 1580 4220 1590
rect 4660 1580 4700 1590
rect 4730 1580 4800 1590
rect 4960 1580 5160 1590
rect 5250 1580 5260 1590
rect 5310 1580 5340 1590
rect 5360 1580 5370 1590
rect 5420 1580 5450 1590
rect 5490 1580 5500 1590
rect 5510 1580 5520 1590
rect 5540 1580 5570 1590
rect 5600 1580 5660 1590
rect 5700 1580 5960 1590
rect 6330 1580 6430 1590
rect 6810 1580 6840 1590
rect 7360 1580 7370 1590
rect 7820 1580 7880 1590
rect 8380 1580 8450 1590
rect 9860 1580 9870 1590
rect 9920 1580 9940 1590
rect 1950 1570 1970 1580
rect 3140 1570 3190 1580
rect 4110 1570 4230 1580
rect 4700 1570 4740 1580
rect 4790 1570 4930 1580
rect 5000 1570 5160 1580
rect 5240 1570 5250 1580
rect 5280 1570 5330 1580
rect 5380 1570 5410 1580
rect 5470 1570 5480 1580
rect 5500 1570 5510 1580
rect 5520 1570 5570 1580
rect 5590 1570 5680 1580
rect 5710 1570 5970 1580
rect 6340 1570 6420 1580
rect 6810 1570 6840 1580
rect 7360 1570 7370 1580
rect 7820 1570 7880 1580
rect 8310 1570 8320 1580
rect 8390 1570 8450 1580
rect 9300 1570 9330 1580
rect 9820 1570 9830 1580
rect 9850 1570 9860 1580
rect 1950 1560 1980 1570
rect 3140 1560 3180 1570
rect 4110 1560 4220 1570
rect 4310 1560 4320 1570
rect 4710 1560 4730 1570
rect 4780 1560 4790 1570
rect 4800 1560 4830 1570
rect 4840 1560 4960 1570
rect 4970 1560 4980 1570
rect 5060 1560 5260 1570
rect 5280 1560 5350 1570
rect 5370 1560 5380 1570
rect 5390 1560 5410 1570
rect 5420 1560 5430 1570
rect 5480 1560 5490 1570
rect 5520 1560 5560 1570
rect 5590 1560 5630 1570
rect 5660 1560 5690 1570
rect 5710 1560 5960 1570
rect 6340 1560 6400 1570
rect 6800 1560 6830 1570
rect 7830 1560 7890 1570
rect 8310 1560 8320 1570
rect 8390 1560 8450 1570
rect 9730 1560 9740 1570
rect 9840 1560 9850 1570
rect 1960 1550 1990 1560
rect 3120 1550 3180 1560
rect 4130 1550 4240 1560
rect 4810 1550 4830 1560
rect 4850 1550 4990 1560
rect 5000 1550 5030 1560
rect 5100 1550 5260 1560
rect 5280 1550 5300 1560
rect 5320 1550 5330 1560
rect 5360 1550 5370 1560
rect 5380 1550 5430 1560
rect 5440 1550 5450 1560
rect 5460 1550 5480 1560
rect 5500 1550 5560 1560
rect 5580 1550 5610 1560
rect 5620 1550 5630 1560
rect 5670 1550 5700 1560
rect 5720 1550 5810 1560
rect 5820 1550 5980 1560
rect 6330 1550 6400 1560
rect 6810 1550 6840 1560
rect 7840 1550 7890 1560
rect 8310 1550 8320 1560
rect 8390 1550 8460 1560
rect 9840 1550 9850 1560
rect 1970 1540 2000 1550
rect 3110 1540 3170 1550
rect 4120 1540 4240 1550
rect 4820 1540 4980 1550
rect 5000 1540 5070 1550
rect 5120 1540 5270 1550
rect 5350 1540 5560 1550
rect 5580 1540 5610 1550
rect 5650 1540 5660 1550
rect 5720 1540 5960 1550
rect 6340 1540 6410 1550
rect 6800 1540 6830 1550
rect 7840 1540 7880 1550
rect 8370 1540 8440 1550
rect 9800 1540 9810 1550
rect 9920 1540 9930 1550
rect 1970 1530 2010 1540
rect 3100 1530 3160 1540
rect 4130 1530 4250 1540
rect 4330 1530 4340 1540
rect 4870 1530 4890 1540
rect 4910 1530 4920 1540
rect 4940 1530 4980 1540
rect 5000 1530 5120 1540
rect 5150 1530 5280 1540
rect 5320 1530 5330 1540
rect 5340 1530 5560 1540
rect 5590 1530 5610 1540
rect 5700 1530 5710 1540
rect 5730 1530 5920 1540
rect 5930 1530 5960 1540
rect 5970 1530 5980 1540
rect 6340 1530 6410 1540
rect 6800 1530 6830 1540
rect 7830 1530 7880 1540
rect 8300 1530 8310 1540
rect 8380 1530 8450 1540
rect 9490 1530 9530 1540
rect 9790 1530 9800 1540
rect 9830 1530 9840 1540
rect 9980 1530 9990 1540
rect 1980 1520 2010 1530
rect 3090 1520 3150 1530
rect 4140 1520 4250 1530
rect 4330 1520 4340 1530
rect 4910 1520 4920 1530
rect 4950 1520 4970 1530
rect 5000 1520 5140 1530
rect 5180 1520 5290 1530
rect 5340 1520 5560 1530
rect 5640 1520 5660 1530
rect 5700 1520 5710 1530
rect 5730 1520 5880 1530
rect 5890 1520 5960 1530
rect 5970 1520 5980 1530
rect 5990 1520 6010 1530
rect 6340 1520 6400 1530
rect 6800 1520 6830 1530
rect 7840 1520 7880 1530
rect 8300 1520 8310 1530
rect 8370 1520 8450 1530
rect 9000 1520 9010 1530
rect 9490 1520 9510 1530
rect 9790 1520 9800 1530
rect 9930 1520 9940 1530
rect 9980 1520 9990 1530
rect 1990 1510 2020 1520
rect 3080 1510 3140 1520
rect 4130 1510 4140 1520
rect 4150 1510 4240 1520
rect 4960 1510 4980 1520
rect 5000 1510 5170 1520
rect 5200 1510 5310 1520
rect 5330 1510 5560 1520
rect 5630 1510 5660 1520
rect 5690 1510 5700 1520
rect 5720 1510 5940 1520
rect 5950 1510 5960 1520
rect 6340 1510 6380 1520
rect 6800 1510 6820 1520
rect 7830 1510 7890 1520
rect 8300 1510 8310 1520
rect 8380 1510 8450 1520
rect 9000 1510 9010 1520
rect 9490 1510 9500 1520
rect 9890 1510 9910 1520
rect 9940 1510 9960 1520
rect 9970 1510 9980 1520
rect 1990 1500 2020 1510
rect 3070 1500 3120 1510
rect 4930 1500 4980 1510
rect 5000 1500 5190 1510
rect 5230 1500 5450 1510
rect 5490 1500 5560 1510
rect 5630 1500 5660 1510
rect 5680 1500 5700 1510
rect 5730 1500 5940 1510
rect 6340 1500 6380 1510
rect 6800 1500 6820 1510
rect 7370 1500 7380 1510
rect 7840 1500 7880 1510
rect 8300 1500 8310 1510
rect 8360 1500 8450 1510
rect 9490 1500 9500 1510
rect 9880 1500 9900 1510
rect 9930 1500 9940 1510
rect 9970 1500 9980 1510
rect 2000 1490 2040 1500
rect 3060 1490 3110 1500
rect 4940 1490 4950 1500
rect 4960 1490 4980 1500
rect 5000 1490 5010 1500
rect 5020 1490 5220 1500
rect 5250 1490 5450 1500
rect 5510 1490 5560 1500
rect 5580 1490 5600 1500
rect 5630 1490 5670 1500
rect 5690 1490 5700 1500
rect 5730 1490 5960 1500
rect 6340 1490 6380 1500
rect 6800 1490 6820 1500
rect 7370 1490 7380 1500
rect 7830 1490 7890 1500
rect 8290 1490 8300 1500
rect 8360 1490 8450 1500
rect 9220 1490 9230 1500
rect 9770 1490 9780 1500
rect 9870 1490 9890 1500
rect 2010 1480 2040 1490
rect 2950 1480 2960 1490
rect 2980 1480 3010 1490
rect 3050 1480 3110 1490
rect 4350 1480 4360 1490
rect 4940 1480 4950 1490
rect 4960 1480 4970 1490
rect 4990 1480 5010 1490
rect 5020 1480 5030 1490
rect 5040 1480 5070 1490
rect 5090 1480 5110 1490
rect 5120 1480 5240 1490
rect 5270 1480 5450 1490
rect 5510 1480 5560 1490
rect 5590 1480 5600 1490
rect 5630 1480 5670 1490
rect 5710 1480 5720 1490
rect 5730 1480 5850 1490
rect 5880 1480 5890 1490
rect 5940 1480 5960 1490
rect 6330 1480 6370 1490
rect 6800 1480 6820 1490
rect 7370 1480 7380 1490
rect 7830 1480 7890 1490
rect 8290 1480 8300 1490
rect 8360 1480 8450 1490
rect 9220 1480 9230 1490
rect 9870 1480 9890 1490
rect 9900 1480 9910 1490
rect 9920 1480 9930 1490
rect 2020 1470 2060 1480
rect 2940 1470 3000 1480
rect 3020 1470 3100 1480
rect 4960 1470 4970 1480
rect 4990 1470 5260 1480
rect 5290 1470 5450 1480
rect 5460 1470 5470 1480
rect 5490 1470 5500 1480
rect 5510 1470 5560 1480
rect 5580 1470 5600 1480
rect 5630 1470 5680 1480
rect 5720 1470 5730 1480
rect 5740 1470 5870 1480
rect 5880 1470 5890 1480
rect 6330 1470 6370 1480
rect 6800 1470 6810 1480
rect 7370 1470 7380 1480
rect 7850 1470 7900 1480
rect 8280 1470 8310 1480
rect 8370 1470 8450 1480
rect 9570 1470 9580 1480
rect 9600 1470 9640 1480
rect 9760 1470 9770 1480
rect 9910 1470 9920 1480
rect 910 1460 980 1470
rect 2030 1460 2070 1470
rect 2920 1460 3090 1470
rect 4140 1460 4150 1470
rect 4960 1460 4970 1470
rect 4990 1460 5010 1470
rect 5030 1460 5280 1470
rect 5300 1460 5450 1470
rect 5460 1460 5480 1470
rect 5490 1460 5500 1470
rect 5510 1460 5560 1470
rect 5580 1460 5600 1470
rect 5630 1460 5700 1470
rect 5720 1460 5880 1470
rect 6330 1460 6360 1470
rect 6800 1460 6810 1470
rect 7370 1460 7380 1470
rect 7840 1460 7900 1470
rect 8280 1460 8300 1470
rect 8370 1460 8450 1470
rect 9580 1460 9590 1470
rect 9790 1460 9800 1470
rect 890 1450 900 1460
rect 940 1450 990 1460
rect 2040 1450 2080 1460
rect 2910 1450 3070 1460
rect 4360 1450 4370 1460
rect 4780 1450 4830 1460
rect 4840 1450 4850 1460
rect 4880 1450 4890 1460
rect 4960 1450 4970 1460
rect 4990 1450 5010 1460
rect 5060 1450 5080 1460
rect 5100 1450 5110 1460
rect 5120 1450 5290 1460
rect 5310 1450 5450 1460
rect 5470 1450 5480 1460
rect 5510 1450 5550 1460
rect 5570 1450 5600 1460
rect 5630 1450 5700 1460
rect 5710 1450 5890 1460
rect 6340 1450 6360 1460
rect 6800 1450 6810 1460
rect 7360 1450 7370 1460
rect 7850 1450 7900 1460
rect 8280 1450 8300 1460
rect 8370 1450 8450 1460
rect 870 1440 880 1450
rect 890 1440 920 1450
rect 930 1440 940 1450
rect 970 1440 1000 1450
rect 2040 1440 2080 1450
rect 2910 1440 3060 1450
rect 4830 1440 4840 1450
rect 4890 1440 4900 1450
rect 4950 1440 4970 1450
rect 4990 1440 5010 1450
rect 5020 1440 5030 1450
rect 5050 1440 5140 1450
rect 5170 1440 5220 1450
rect 5230 1440 5300 1450
rect 5320 1440 5450 1450
rect 5470 1440 5490 1450
rect 5510 1440 5550 1450
rect 5570 1440 5580 1450
rect 5630 1440 5900 1450
rect 6330 1440 6350 1450
rect 6800 1440 6810 1450
rect 7840 1440 7900 1450
rect 8280 1440 8300 1450
rect 8360 1440 8440 1450
rect 9370 1440 9380 1450
rect 9580 1440 9590 1450
rect 9700 1440 9710 1450
rect 9740 1440 9750 1450
rect 860 1430 1010 1440
rect 2050 1430 2100 1440
rect 2890 1430 3050 1440
rect 4150 1430 4160 1440
rect 4840 1430 4850 1440
rect 4860 1430 4870 1440
rect 4890 1430 4900 1440
rect 4950 1430 4970 1440
rect 4990 1430 5000 1440
rect 5070 1430 5140 1440
rect 5170 1430 5310 1440
rect 5330 1430 5450 1440
rect 5470 1430 5490 1440
rect 5510 1430 5550 1440
rect 5620 1430 5890 1440
rect 6800 1430 6810 1440
rect 7850 1430 7890 1440
rect 8270 1430 8300 1440
rect 8360 1430 8440 1440
rect 9360 1430 9370 1440
rect 9610 1430 9620 1440
rect 9640 1430 9650 1440
rect 9740 1430 9750 1440
rect 850 1420 860 1430
rect 870 1420 1010 1430
rect 2060 1420 2120 1430
rect 2890 1420 3040 1430
rect 4640 1420 4650 1430
rect 4860 1420 4870 1430
rect 4890 1420 4900 1430
rect 4980 1420 4990 1430
rect 5100 1420 5120 1430
rect 5130 1420 5150 1430
rect 5160 1420 5320 1430
rect 5350 1420 5450 1430
rect 5480 1420 5490 1430
rect 5580 1420 5600 1430
rect 5620 1420 5890 1430
rect 6800 1420 6810 1430
rect 7370 1420 7390 1430
rect 7860 1420 7910 1430
rect 8270 1420 8290 1430
rect 8360 1420 8440 1430
rect 9500 1420 9520 1430
rect 9640 1420 9650 1430
rect 9840 1420 9850 1430
rect 850 1410 1000 1420
rect 2070 1410 2120 1420
rect 2870 1410 3030 1420
rect 4810 1410 4830 1420
rect 4900 1410 4910 1420
rect 4950 1410 4960 1420
rect 4980 1410 5000 1420
rect 5080 1410 5090 1420
rect 5110 1410 5120 1420
rect 5150 1410 5340 1420
rect 5350 1410 5450 1420
rect 5480 1410 5500 1420
rect 5580 1410 5590 1420
rect 5630 1410 5930 1420
rect 6800 1410 6810 1420
rect 7370 1410 7390 1420
rect 7850 1410 7910 1420
rect 8270 1410 8290 1420
rect 8360 1410 8460 1420
rect 9490 1410 9500 1420
rect 9540 1410 9550 1420
rect 9620 1410 9640 1420
rect 9760 1410 9770 1420
rect 850 1400 990 1410
rect 2080 1400 2130 1410
rect 2870 1400 3020 1410
rect 4160 1400 4170 1410
rect 4810 1400 4830 1410
rect 4850 1400 4860 1410
rect 4950 1400 4960 1410
rect 4980 1400 4990 1410
rect 5070 1400 5080 1410
rect 5100 1400 5180 1410
rect 5190 1400 5340 1410
rect 5370 1400 5460 1410
rect 5480 1400 5500 1410
rect 5510 1400 5520 1410
rect 5540 1400 5550 1410
rect 5570 1400 5590 1410
rect 5610 1400 5620 1410
rect 5630 1400 5890 1410
rect 5900 1400 5910 1410
rect 7380 1400 7390 1410
rect 7860 1400 7910 1410
rect 8260 1400 8290 1410
rect 8360 1400 8440 1410
rect 8460 1400 8470 1410
rect 9230 1400 9240 1410
rect 9720 1400 9730 1410
rect 9930 1400 9940 1410
rect 840 1390 990 1400
rect 2090 1390 2150 1400
rect 2860 1390 3000 1400
rect 4380 1390 4390 1400
rect 4680 1390 4710 1400
rect 4810 1390 4820 1400
rect 4850 1390 4860 1400
rect 4930 1390 4940 1400
rect 4980 1390 4990 1400
rect 5090 1390 5110 1400
rect 5120 1390 5170 1400
rect 5190 1390 5350 1400
rect 5380 1390 5460 1400
rect 5490 1390 5510 1400
rect 5560 1390 5580 1400
rect 5620 1390 5890 1400
rect 6810 1390 6820 1400
rect 7380 1390 7390 1400
rect 7860 1390 7910 1400
rect 8260 1390 8280 1400
rect 8360 1390 8440 1400
rect 9220 1390 9230 1400
rect 9250 1390 9260 1400
rect 9290 1390 9300 1400
rect 9710 1390 9720 1400
rect 9750 1390 9760 1400
rect 9930 1390 9940 1400
rect 9950 1390 9990 1400
rect 840 1380 990 1390
rect 2100 1380 2160 1390
rect 2850 1380 2990 1390
rect 4840 1380 4860 1390
rect 4980 1380 4990 1390
rect 5140 1380 5150 1390
rect 5160 1380 5370 1390
rect 5390 1380 5470 1390
rect 5490 1380 5520 1390
rect 5540 1380 5570 1390
rect 5620 1380 5890 1390
rect 6810 1380 6820 1390
rect 7860 1380 7910 1390
rect 8250 1380 8290 1390
rect 8320 1380 8330 1390
rect 8340 1380 8460 1390
rect 9270 1380 9280 1390
rect 9290 1380 9300 1390
rect 9550 1380 9560 1390
rect 9680 1380 9690 1390
rect 9710 1380 9720 1390
rect 9930 1380 9950 1390
rect 9990 1380 9990 1390
rect 840 1370 980 1380
rect 2110 1370 2170 1380
rect 2840 1370 2890 1380
rect 2910 1370 2970 1380
rect 4210 1370 4240 1380
rect 4390 1370 4400 1380
rect 4790 1370 4810 1380
rect 4980 1370 4990 1380
rect 5120 1370 5150 1380
rect 5160 1370 5190 1380
rect 5200 1370 5270 1380
rect 5280 1370 5380 1380
rect 5400 1370 5500 1380
rect 5520 1370 5560 1380
rect 5620 1370 5920 1380
rect 6810 1370 6820 1380
rect 7380 1370 7390 1380
rect 7860 1370 7920 1380
rect 8240 1370 8290 1380
rect 8320 1370 8460 1380
rect 9260 1370 9280 1380
rect 9700 1370 9710 1380
rect 9740 1370 9750 1380
rect 9810 1370 9820 1380
rect 9960 1370 9970 1380
rect 840 1360 960 1370
rect 2120 1360 2180 1370
rect 2820 1360 2860 1370
rect 2900 1360 2950 1370
rect 4200 1360 4260 1370
rect 4820 1360 4830 1370
rect 4910 1360 4920 1370
rect 4950 1360 4960 1370
rect 4980 1360 4990 1370
rect 5120 1360 5250 1370
rect 5260 1360 5270 1370
rect 5290 1360 5400 1370
rect 5420 1360 5490 1370
rect 5610 1360 5920 1370
rect 6810 1360 6820 1370
rect 7860 1360 7920 1370
rect 8230 1360 8280 1370
rect 8340 1360 8440 1370
rect 9700 1360 9710 1370
rect 9800 1360 9810 1370
rect 840 1350 940 1360
rect 2130 1350 2190 1360
rect 2820 1350 2850 1360
rect 2910 1350 2940 1360
rect 3560 1350 3570 1360
rect 4180 1350 4190 1360
rect 4200 1350 4260 1360
rect 4820 1350 4830 1360
rect 4920 1350 4950 1360
rect 5110 1350 5120 1360
rect 5130 1350 5180 1360
rect 5220 1350 5410 1360
rect 5430 1350 5490 1360
rect 5600 1350 5930 1360
rect 5950 1350 5960 1360
rect 6810 1350 6820 1360
rect 7380 1350 7400 1360
rect 7860 1350 7920 1360
rect 8210 1350 8270 1360
rect 8340 1350 8440 1360
rect 9670 1350 9680 1360
rect 9800 1350 9810 1360
rect 840 1340 940 1350
rect 2140 1340 2220 1350
rect 2240 1340 2250 1350
rect 2800 1340 2840 1350
rect 3540 1340 3550 1350
rect 4200 1340 4270 1350
rect 4400 1340 4410 1350
rect 4940 1340 4950 1350
rect 4970 1340 4980 1350
rect 5080 1340 5090 1350
rect 5100 1340 5140 1350
rect 5210 1340 5420 1350
rect 5440 1340 5520 1350
rect 5540 1340 5570 1350
rect 5590 1340 5930 1350
rect 7380 1340 7400 1350
rect 7860 1340 7920 1350
rect 8200 1340 8280 1350
rect 8310 1340 8430 1350
rect 9260 1340 9270 1350
rect 9680 1340 9700 1350
rect 9730 1340 9740 1350
rect 9790 1340 9800 1350
rect 9830 1340 9840 1350
rect 9960 1340 9970 1350
rect 840 1330 930 1340
rect 2150 1330 2220 1340
rect 2790 1330 2820 1340
rect 3640 1330 3650 1340
rect 4220 1330 4270 1340
rect 4970 1330 4980 1340
rect 5100 1330 5200 1340
rect 5210 1330 5220 1340
rect 5250 1330 5380 1340
rect 5390 1330 5430 1340
rect 5450 1330 5530 1340
rect 5570 1330 5930 1340
rect 7380 1330 7400 1340
rect 7860 1330 7910 1340
rect 8190 1330 8440 1340
rect 9670 1330 9690 1340
rect 830 1320 930 1330
rect 2150 1320 2230 1330
rect 2290 1320 2300 1330
rect 2770 1320 2810 1330
rect 4850 1320 4860 1330
rect 4940 1320 4950 1330
rect 4970 1320 4990 1330
rect 5070 1320 5180 1330
rect 5190 1320 5200 1330
rect 5240 1320 5440 1330
rect 5460 1320 5930 1330
rect 7380 1320 7400 1330
rect 7860 1320 7920 1330
rect 8190 1320 8440 1330
rect 9090 1320 9100 1330
rect 9380 1320 9390 1330
rect 9670 1320 9680 1330
rect 9990 1320 9990 1330
rect 830 1310 920 1320
rect 2160 1310 2260 1320
rect 2280 1310 2340 1320
rect 2750 1310 2790 1320
rect 4410 1310 4420 1320
rect 4970 1310 4990 1320
rect 5050 1310 5120 1320
rect 5140 1310 5210 1320
rect 5230 1310 5240 1320
rect 5250 1310 5300 1320
rect 5320 1310 5440 1320
rect 5470 1310 5930 1320
rect 7380 1310 7400 1320
rect 7860 1310 7920 1320
rect 8180 1310 8420 1320
rect 8440 1310 8460 1320
rect 9080 1310 9100 1320
rect 9260 1310 9270 1320
rect 9640 1310 9660 1320
rect 9990 1310 9990 1320
rect 830 1300 920 1310
rect 2170 1300 2270 1310
rect 2280 1300 2360 1310
rect 2720 1300 2790 1310
rect 4970 1300 4980 1310
rect 5030 1300 5110 1310
rect 5160 1300 5210 1310
rect 5260 1300 5300 1310
rect 5310 1300 5450 1310
rect 5470 1300 5520 1310
rect 5600 1300 5920 1310
rect 6820 1300 6830 1310
rect 7380 1300 7400 1310
rect 7870 1300 7920 1310
rect 8180 1300 8420 1310
rect 8430 1300 8440 1310
rect 9080 1300 9120 1310
rect 9670 1300 9680 1310
rect 9820 1300 9840 1310
rect 9990 1300 9990 1310
rect 820 1290 920 1300
rect 2180 1290 2400 1300
rect 2710 1290 2760 1300
rect 3690 1290 3700 1300
rect 4940 1290 4950 1300
rect 4970 1290 4980 1300
rect 5010 1290 5090 1300
rect 5170 1290 5370 1300
rect 5680 1290 5920 1300
rect 7380 1290 7400 1300
rect 7870 1290 7920 1300
rect 8170 1290 8430 1300
rect 9080 1290 9120 1300
rect 9580 1290 9590 1300
rect 9820 1290 9830 1300
rect 9960 1290 9990 1300
rect 820 1280 920 1290
rect 2190 1280 2430 1290
rect 2680 1280 2740 1290
rect 4420 1280 4430 1290
rect 4930 1280 4940 1290
rect 4960 1280 4990 1290
rect 5000 1280 5130 1290
rect 5150 1280 5200 1290
rect 5440 1280 5670 1290
rect 5700 1280 5920 1290
rect 7380 1280 7410 1290
rect 7880 1280 7920 1290
rect 8180 1280 8440 1290
rect 9080 1280 9120 1290
rect 9130 1280 9140 1290
rect 9660 1280 9670 1290
rect 9690 1280 9700 1290
rect 9750 1280 9760 1290
rect 820 1270 920 1280
rect 2200 1270 2440 1280
rect 2490 1270 2500 1280
rect 2660 1270 2720 1280
rect 3500 1270 3510 1280
rect 4930 1270 4940 1280
rect 4960 1270 5120 1280
rect 5290 1270 5680 1280
rect 5700 1270 5930 1280
rect 7380 1270 7400 1280
rect 7880 1270 7920 1280
rect 8170 1270 8450 1280
rect 8990 1270 9000 1280
rect 9070 1270 9120 1280
rect 9480 1270 9490 1280
rect 9650 1270 9660 1280
rect 9830 1270 9840 1280
rect 820 1260 920 1270
rect 2200 1260 2700 1270
rect 3500 1260 3510 1270
rect 4930 1260 4940 1270
rect 4960 1260 5040 1270
rect 5170 1260 5340 1270
rect 5350 1260 5430 1270
rect 5450 1260 5680 1270
rect 5690 1260 5930 1270
rect 7380 1260 7410 1270
rect 7880 1260 7920 1270
rect 8180 1260 8450 1270
rect 9070 1260 9120 1270
rect 9130 1260 9140 1270
rect 9490 1260 9500 1270
rect 9680 1260 9690 1270
rect 9830 1260 9840 1270
rect 9950 1260 9960 1270
rect 9970 1260 9990 1270
rect 820 1250 920 1260
rect 2210 1250 2680 1260
rect 4200 1250 4210 1260
rect 4430 1250 4440 1260
rect 4930 1250 4940 1260
rect 5130 1250 5240 1260
rect 5250 1250 5270 1260
rect 5280 1250 5290 1260
rect 5330 1250 5340 1260
rect 5350 1250 5370 1260
rect 5380 1250 5390 1260
rect 5410 1250 5420 1260
rect 5450 1250 5670 1260
rect 5690 1250 5920 1260
rect 7380 1250 7410 1260
rect 7880 1250 7940 1260
rect 8180 1250 8460 1260
rect 8980 1250 8990 1260
rect 9010 1250 9020 1260
rect 9070 1250 9120 1260
rect 9310 1250 9320 1260
rect 9490 1250 9500 1260
rect 9640 1250 9650 1260
rect 9830 1250 9840 1260
rect 9970 1250 9990 1260
rect 810 1240 910 1250
rect 2200 1240 2210 1250
rect 2220 1240 2650 1250
rect 3750 1240 3760 1250
rect 4200 1240 4210 1250
rect 4430 1240 4440 1250
rect 5050 1240 5150 1250
rect 5160 1240 5190 1250
rect 5200 1240 5210 1250
rect 5220 1240 5240 1250
rect 5250 1240 5270 1250
rect 5280 1240 5290 1250
rect 5330 1240 5340 1250
rect 5350 1240 5370 1250
rect 5410 1240 5420 1250
rect 5440 1240 5680 1250
rect 5690 1240 5910 1250
rect 5930 1240 5940 1250
rect 6770 1240 6790 1250
rect 6820 1240 6830 1250
rect 7380 1240 7400 1250
rect 7880 1240 7940 1250
rect 8180 1240 8460 1250
rect 8900 1240 8910 1250
rect 8940 1240 9000 1250
rect 9010 1240 9020 1250
rect 9070 1240 9120 1250
rect 9630 1240 9640 1250
rect 9670 1240 9680 1250
rect 9970 1240 9990 1250
rect 810 1230 910 1240
rect 2250 1230 2640 1240
rect 3510 1230 3520 1240
rect 3540 1230 3590 1240
rect 4760 1230 4810 1240
rect 5000 1230 5060 1240
rect 5070 1230 5110 1240
rect 5130 1230 5140 1240
rect 5160 1230 5180 1240
rect 5200 1230 5210 1240
rect 5220 1230 5240 1240
rect 5260 1230 5270 1240
rect 5350 1230 5370 1240
rect 5390 1230 5400 1240
rect 5410 1230 5430 1240
rect 5450 1230 5680 1240
rect 5690 1230 5910 1240
rect 5930 1230 5940 1240
rect 6750 1230 6790 1240
rect 6820 1230 6830 1240
rect 7390 1230 7410 1240
rect 7890 1230 7950 1240
rect 8180 1230 8400 1240
rect 8410 1230 8450 1240
rect 8940 1230 9020 1240
rect 9030 1230 9040 1240
rect 9070 1230 9120 1240
rect 9610 1230 9620 1240
rect 9720 1230 9730 1240
rect 810 1220 900 1230
rect 2270 1220 2630 1230
rect 3530 1220 3660 1230
rect 4910 1220 5030 1230
rect 5050 1220 5060 1230
rect 5080 1220 5090 1230
rect 5100 1220 5110 1230
rect 5130 1220 5140 1230
rect 5150 1220 5180 1230
rect 5230 1220 5240 1230
rect 5260 1220 5270 1230
rect 5310 1220 5320 1230
rect 5360 1220 5370 1230
rect 5390 1220 5400 1230
rect 5410 1220 5440 1230
rect 5460 1220 5680 1230
rect 5690 1220 5910 1230
rect 6740 1220 6760 1230
rect 6770 1220 6800 1230
rect 6820 1220 6830 1230
rect 7390 1220 7410 1230
rect 7890 1220 7950 1230
rect 8180 1220 8400 1230
rect 8410 1220 8450 1230
rect 8880 1220 8900 1230
rect 8920 1220 8970 1230
rect 8980 1220 9010 1230
rect 9060 1220 9110 1230
rect 9620 1220 9630 1230
rect 9660 1220 9670 1230
rect 810 1210 900 1220
rect 2140 1210 2160 1220
rect 2230 1210 2240 1220
rect 2300 1210 2630 1220
rect 3520 1210 3530 1220
rect 3540 1210 3660 1220
rect 4830 1210 4840 1220
rect 4850 1210 4880 1220
rect 4900 1210 4950 1220
rect 4970 1210 4980 1220
rect 5010 1210 5020 1220
rect 5040 1210 5060 1220
rect 5070 1210 5080 1220
rect 5130 1210 5140 1220
rect 5160 1210 5190 1220
rect 5230 1210 5240 1220
rect 5260 1210 5270 1220
rect 5420 1210 5430 1220
rect 5460 1210 5680 1220
rect 5690 1210 5890 1220
rect 6730 1210 6740 1220
rect 6790 1210 6800 1220
rect 6820 1210 6830 1220
rect 7380 1210 7410 1220
rect 7890 1210 7950 1220
rect 8180 1210 8410 1220
rect 8430 1210 8440 1220
rect 8900 1210 8950 1220
rect 8980 1210 9000 1220
rect 9070 1210 9110 1220
rect 9320 1210 9330 1220
rect 9650 1210 9660 1220
rect 9710 1210 9720 1220
rect 9820 1210 9830 1220
rect 800 1200 890 1210
rect 2110 1200 2180 1210
rect 2190 1200 2250 1210
rect 2330 1200 2600 1210
rect 2610 1200 2620 1210
rect 3530 1200 3670 1210
rect 4440 1200 4450 1210
rect 4760 1200 4870 1210
rect 4890 1200 4900 1210
rect 4920 1200 4930 1210
rect 4980 1200 4990 1210
rect 5010 1200 5020 1210
rect 5030 1200 5060 1210
rect 5080 1200 5090 1210
rect 5100 1200 5110 1210
rect 5130 1200 5140 1210
rect 5160 1200 5170 1210
rect 5310 1200 5320 1210
rect 5370 1200 5400 1210
rect 5420 1200 5440 1210
rect 5450 1200 5680 1210
rect 5700 1200 5910 1210
rect 6720 1200 6730 1210
rect 6790 1200 6800 1210
rect 6820 1200 6830 1210
rect 7380 1200 7410 1210
rect 7900 1200 7950 1210
rect 8180 1200 8380 1210
rect 8860 1200 8950 1210
rect 8970 1200 8990 1210
rect 9000 1200 9020 1210
rect 9040 1200 9060 1210
rect 9070 1200 9110 1210
rect 9820 1200 9830 1210
rect 9910 1200 9920 1210
rect 9950 1200 9960 1210
rect 800 1190 890 1200
rect 2100 1190 2250 1200
rect 2420 1190 2430 1200
rect 2450 1190 2490 1200
rect 2500 1190 2510 1200
rect 3550 1190 3680 1200
rect 4710 1190 4770 1200
rect 4780 1190 4800 1200
rect 4820 1190 4830 1200
rect 4840 1190 4850 1200
rect 4980 1190 4990 1200
rect 5050 1190 5060 1200
rect 5070 1190 5090 1200
rect 5100 1190 5110 1200
rect 5130 1190 5140 1200
rect 5150 1190 5160 1200
rect 5210 1190 5220 1200
rect 5230 1190 5680 1200
rect 5700 1190 5910 1200
rect 6700 1190 6720 1200
rect 6790 1190 6800 1200
rect 7380 1190 7410 1200
rect 7900 1190 7950 1200
rect 8180 1190 8400 1200
rect 8420 1190 8430 1200
rect 8500 1190 8520 1200
rect 8810 1190 8850 1200
rect 8860 1190 8960 1200
rect 8980 1190 8990 1200
rect 9040 1190 9110 1200
rect 9300 1190 9310 1200
rect 9700 1190 9710 1200
rect 9990 1190 9990 1200
rect 790 1180 870 1190
rect 2100 1180 2250 1190
rect 3560 1180 3700 1190
rect 3840 1180 3850 1190
rect 4210 1180 4220 1190
rect 4670 1180 4690 1190
rect 4700 1180 4720 1190
rect 4780 1180 4800 1190
rect 4840 1180 4850 1190
rect 4860 1180 4870 1190
rect 4890 1180 4900 1190
rect 4980 1180 4990 1190
rect 5020 1180 5030 1190
rect 5050 1180 5060 1190
rect 5080 1180 5090 1190
rect 5130 1180 5170 1190
rect 5180 1180 5210 1190
rect 5300 1180 5680 1190
rect 5700 1180 5880 1190
rect 6690 1180 6710 1190
rect 6790 1180 6800 1190
rect 7380 1180 7420 1190
rect 7900 1180 7950 1190
rect 8180 1180 8380 1190
rect 8410 1180 8430 1190
rect 8470 1180 8480 1190
rect 8550 1180 8570 1190
rect 8750 1180 8770 1190
rect 8810 1180 9000 1190
rect 9020 1180 9110 1190
rect 9310 1180 9320 1190
rect 9640 1180 9650 1190
rect 9970 1180 9980 1190
rect 810 1170 870 1180
rect 2080 1170 2270 1180
rect 3570 1170 3720 1180
rect 4210 1170 4220 1180
rect 4570 1170 4580 1180
rect 4590 1170 4600 1180
rect 4620 1170 4640 1180
rect 4650 1170 4670 1180
rect 4690 1170 4700 1180
rect 4740 1170 4770 1180
rect 4780 1170 4800 1180
rect 4810 1170 4820 1180
rect 4830 1170 4850 1180
rect 4860 1170 4880 1180
rect 4980 1170 4990 1180
rect 5020 1170 5030 1180
rect 5050 1170 5070 1180
rect 5080 1170 5090 1180
rect 5110 1170 5130 1180
rect 5330 1170 5370 1180
rect 5380 1170 5680 1180
rect 5700 1170 5880 1180
rect 6670 1170 6690 1180
rect 6790 1170 6800 1180
rect 7380 1170 7420 1180
rect 7910 1170 7960 1180
rect 8180 1170 8370 1180
rect 8410 1170 8450 1180
rect 8750 1170 8790 1180
rect 8800 1170 9110 1180
rect 9140 1170 9150 1180
rect 9360 1170 9370 1180
rect 9500 1170 9510 1180
rect 9690 1170 9700 1180
rect 9810 1170 9820 1180
rect 780 1160 790 1170
rect 820 1160 870 1170
rect 2070 1160 2280 1170
rect 3580 1160 3730 1170
rect 4560 1160 4570 1170
rect 4580 1160 4600 1170
rect 4610 1160 4650 1170
rect 4680 1160 4700 1170
rect 4740 1160 4750 1170
rect 4760 1160 4770 1170
rect 4790 1160 4800 1170
rect 4810 1160 4820 1170
rect 4840 1160 4850 1170
rect 4860 1160 4890 1170
rect 4900 1160 4910 1170
rect 4980 1160 4990 1170
rect 5000 1160 5050 1170
rect 5390 1160 5420 1170
rect 5430 1160 5680 1170
rect 5700 1160 5880 1170
rect 5890 1160 5900 1170
rect 6660 1160 6670 1170
rect 7380 1160 7420 1170
rect 7910 1160 7960 1170
rect 8170 1160 8380 1170
rect 8410 1160 8430 1170
rect 8520 1160 8530 1170
rect 8540 1160 8550 1170
rect 8730 1160 8770 1170
rect 8790 1160 9110 1170
rect 830 1150 870 1160
rect 2070 1150 2290 1160
rect 3570 1150 3740 1160
rect 4560 1150 4580 1160
rect 4590 1150 4600 1160
rect 4610 1150 4650 1160
rect 4680 1150 4700 1160
rect 4720 1150 4730 1160
rect 4740 1150 4770 1160
rect 4780 1150 4800 1160
rect 4810 1150 4820 1160
rect 4830 1150 4840 1160
rect 4860 1150 4870 1160
rect 4900 1150 4910 1160
rect 5380 1150 5420 1160
rect 5430 1150 5450 1160
rect 5460 1150 5680 1160
rect 5700 1150 5840 1160
rect 5860 1150 5920 1160
rect 6640 1150 6660 1160
rect 6790 1150 6810 1160
rect 7380 1150 7420 1160
rect 7910 1150 7950 1160
rect 8170 1150 8380 1160
rect 8400 1150 8430 1160
rect 8720 1150 8750 1160
rect 8780 1150 9110 1160
rect 9370 1150 9380 1160
rect 9620 1150 9630 1160
rect 770 1140 780 1150
rect 830 1140 880 1150
rect 2050 1140 2330 1150
rect 3580 1140 3740 1150
rect 4560 1140 4580 1150
rect 4590 1140 4600 1150
rect 4620 1140 4640 1150
rect 4650 1140 4660 1150
rect 4680 1140 4700 1150
rect 4720 1140 4730 1150
rect 4740 1140 4750 1150
rect 4760 1140 4770 1150
rect 4790 1140 4800 1150
rect 4830 1140 4840 1150
rect 4860 1140 4880 1150
rect 4890 1140 4900 1150
rect 5400 1140 5430 1150
rect 5440 1140 5450 1150
rect 5460 1140 5620 1150
rect 5670 1140 5680 1150
rect 5700 1140 5890 1150
rect 5900 1140 5920 1150
rect 6630 1140 6640 1150
rect 6800 1140 6810 1150
rect 7380 1140 7420 1150
rect 7910 1140 7950 1150
rect 8170 1140 8380 1150
rect 8510 1140 8520 1150
rect 8710 1140 8760 1150
rect 8770 1140 9110 1150
rect 9150 1140 9160 1150
rect 9320 1140 9330 1150
rect 9380 1140 9390 1150
rect 9540 1140 9550 1150
rect 9580 1140 9590 1150
rect 9920 1140 9930 1150
rect 830 1130 880 1140
rect 2040 1130 2330 1140
rect 3590 1130 3740 1140
rect 4560 1130 4580 1140
rect 4590 1130 4600 1140
rect 4610 1130 4620 1140
rect 4630 1130 4640 1140
rect 4680 1130 4700 1140
rect 4710 1130 4720 1140
rect 4730 1130 4740 1140
rect 4760 1130 4770 1140
rect 4790 1130 4830 1140
rect 5400 1130 5680 1140
rect 5700 1130 5730 1140
rect 5740 1130 5900 1140
rect 5910 1130 5940 1140
rect 6610 1130 6630 1140
rect 6800 1130 6810 1140
rect 7380 1130 7420 1140
rect 7910 1130 7960 1140
rect 8170 1130 8380 1140
rect 8680 1130 9110 1140
rect 9150 1130 9160 1140
rect 9610 1130 9620 1140
rect 9890 1130 9940 1140
rect 9990 1130 9990 1140
rect 830 1120 880 1130
rect 2040 1120 2350 1130
rect 3600 1120 3730 1130
rect 4220 1120 4230 1130
rect 4560 1120 4570 1130
rect 4590 1120 4600 1130
rect 4610 1120 4620 1130
rect 4630 1120 4640 1130
rect 4650 1120 4660 1130
rect 4670 1120 4690 1130
rect 4700 1120 4710 1130
rect 4720 1120 4730 1130
rect 5400 1120 5680 1130
rect 5700 1120 5730 1130
rect 5740 1120 5900 1130
rect 5910 1120 5920 1130
rect 5930 1120 5940 1130
rect 6600 1120 6610 1130
rect 6800 1120 6810 1130
rect 6830 1120 6840 1130
rect 7380 1120 7420 1130
rect 7910 1120 7960 1130
rect 8170 1120 8360 1130
rect 8410 1120 8420 1130
rect 8460 1120 8480 1130
rect 8550 1120 8560 1130
rect 8570 1120 8580 1130
rect 8600 1120 8630 1130
rect 8680 1120 9110 1130
rect 9880 1120 9920 1130
rect 830 1110 880 1120
rect 2030 1110 2350 1120
rect 3610 1110 3720 1120
rect 4220 1110 4230 1120
rect 4560 1110 4570 1120
rect 4580 1110 4590 1120
rect 4600 1110 4610 1120
rect 4620 1110 4630 1120
rect 5400 1110 5410 1120
rect 5440 1110 5520 1120
rect 5530 1110 5620 1120
rect 5630 1110 5680 1120
rect 5700 1110 5800 1120
rect 5810 1110 5900 1120
rect 6580 1110 6590 1120
rect 6800 1110 6810 1120
rect 6830 1110 6840 1120
rect 7380 1110 7420 1120
rect 7910 1110 7960 1120
rect 8160 1110 8350 1120
rect 8460 1110 8470 1120
rect 8480 1110 8490 1120
rect 8540 1110 8550 1120
rect 8680 1110 9110 1120
rect 9880 1110 9900 1120
rect 830 1100 870 1110
rect 1570 1100 1600 1110
rect 2030 1100 2380 1110
rect 2650 1100 2800 1110
rect 3640 1100 3710 1110
rect 4220 1100 4230 1110
rect 5440 1100 5450 1110
rect 5470 1100 5480 1110
rect 5500 1100 5660 1110
rect 5670 1100 5680 1110
rect 5700 1100 5720 1110
rect 5820 1100 5830 1110
rect 5890 1100 5900 1110
rect 6560 1100 6570 1110
rect 6800 1100 6810 1110
rect 6830 1100 6840 1110
rect 7390 1100 7420 1110
rect 7910 1100 7950 1110
rect 8160 1100 8350 1110
rect 8360 1100 8370 1110
rect 8420 1100 8440 1110
rect 8480 1100 8490 1110
rect 8620 1100 8630 1110
rect 8670 1100 9110 1110
rect 9290 1100 9300 1110
rect 9530 1100 9540 1110
rect 9830 1100 9840 1110
rect 9870 1100 9880 1110
rect 9900 1100 9910 1110
rect 830 1090 870 1100
rect 1620 1090 1630 1100
rect 2020 1090 2400 1100
rect 2410 1090 2420 1100
rect 2500 1090 2520 1100
rect 2530 1090 2810 1100
rect 3640 1090 3710 1100
rect 4220 1090 4230 1100
rect 4470 1090 4480 1100
rect 5470 1090 5650 1100
rect 5700 1090 5720 1100
rect 5890 1090 5910 1100
rect 6540 1090 6560 1100
rect 6800 1090 6810 1100
rect 7380 1090 7420 1100
rect 7910 1090 7960 1100
rect 8160 1090 8350 1100
rect 8410 1090 8440 1100
rect 8450 1090 8460 1100
rect 8550 1090 8560 1100
rect 8660 1090 9110 1100
rect 9290 1090 9300 1100
rect 9550 1090 9560 1100
rect 9650 1090 9660 1100
rect 9990 1090 9990 1100
rect 750 1080 760 1090
rect 820 1080 870 1090
rect 1630 1080 1640 1090
rect 2020 1080 2820 1090
rect 3660 1080 3700 1090
rect 5220 1080 5230 1090
rect 5480 1080 5520 1090
rect 5530 1080 5590 1090
rect 5600 1080 5650 1090
rect 5870 1080 5950 1090
rect 6520 1080 6540 1090
rect 6800 1080 6810 1090
rect 6830 1080 6840 1090
rect 7380 1080 7420 1090
rect 7910 1080 7960 1090
rect 8160 1080 8350 1090
rect 8370 1080 8390 1090
rect 8400 1080 8420 1090
rect 8440 1080 8460 1090
rect 8550 1080 8580 1090
rect 8660 1080 9110 1090
rect 9270 1080 9280 1090
rect 9410 1080 9420 1090
rect 9850 1080 9880 1090
rect 9920 1080 9940 1090
rect 750 1070 760 1080
rect 820 1070 860 1080
rect 1630 1070 1640 1080
rect 2020 1070 2160 1080
rect 2180 1070 2840 1080
rect 3660 1070 3670 1080
rect 4000 1070 4010 1080
rect 5200 1070 5210 1080
rect 5440 1070 5450 1080
rect 5470 1070 5490 1080
rect 5520 1070 5590 1080
rect 5670 1070 5680 1080
rect 5700 1070 5710 1080
rect 5850 1070 5870 1080
rect 5880 1070 5990 1080
rect 6010 1070 6030 1080
rect 6500 1070 6520 1080
rect 6800 1070 6810 1080
rect 6830 1070 6840 1080
rect 7390 1070 7420 1080
rect 7920 1070 7960 1080
rect 8160 1070 8360 1080
rect 8370 1070 8380 1080
rect 8390 1070 8400 1080
rect 8410 1070 8430 1080
rect 8440 1070 8460 1080
rect 8500 1070 8520 1080
rect 8550 1070 8570 1080
rect 8590 1070 8610 1080
rect 8660 1070 9110 1080
rect 9260 1070 9270 1080
rect 9410 1070 9420 1080
rect 9540 1070 9550 1080
rect 9840 1070 9850 1080
rect 9860 1070 9880 1080
rect 9890 1070 9920 1080
rect 9940 1070 9950 1080
rect 810 1060 860 1070
rect 1500 1060 1510 1070
rect 1630 1060 1650 1070
rect 2020 1060 2090 1070
rect 2100 1060 2110 1070
rect 2160 1060 2840 1070
rect 3770 1060 3810 1070
rect 4220 1060 4230 1070
rect 5440 1060 5450 1070
rect 5470 1060 5480 1070
rect 5510 1060 5520 1070
rect 5560 1060 5570 1070
rect 5600 1060 5620 1070
rect 5670 1060 5680 1070
rect 5700 1060 5710 1070
rect 5800 1060 5810 1070
rect 5840 1060 5850 1070
rect 5890 1060 5910 1070
rect 5920 1060 5960 1070
rect 6480 1060 6500 1070
rect 6800 1060 6810 1070
rect 6830 1060 6840 1070
rect 7390 1060 7420 1070
rect 7920 1060 7960 1070
rect 8150 1060 8390 1070
rect 8400 1060 8410 1070
rect 8450 1060 8470 1070
rect 8560 1060 8570 1070
rect 8650 1060 9070 1070
rect 9080 1060 9100 1070
rect 9300 1060 9310 1070
rect 9570 1060 9580 1070
rect 9720 1060 9730 1070
rect 9830 1060 9840 1070
rect 9850 1060 9860 1070
rect 9890 1060 9910 1070
rect 810 1050 860 1060
rect 1490 1050 1500 1060
rect 1520 1050 1530 1060
rect 1600 1050 1650 1060
rect 2020 1050 2080 1060
rect 2210 1050 2840 1060
rect 3670 1050 3680 1060
rect 3760 1050 3820 1060
rect 4030 1050 4040 1060
rect 5370 1050 5380 1060
rect 5510 1050 5520 1060
rect 5600 1050 5610 1060
rect 5630 1050 5640 1060
rect 5670 1050 5680 1060
rect 5770 1050 5790 1060
rect 5830 1050 5850 1060
rect 5860 1050 5880 1060
rect 5930 1050 5960 1060
rect 6460 1050 6480 1060
rect 6800 1050 6810 1060
rect 6830 1050 6840 1060
rect 7390 1050 7420 1060
rect 7920 1050 7960 1060
rect 8150 1050 8320 1060
rect 8330 1050 8360 1060
rect 8390 1050 8400 1060
rect 8440 1050 8450 1060
rect 8480 1050 8490 1060
rect 8560 1050 8620 1060
rect 8640 1050 9070 1060
rect 9080 1050 9110 1060
rect 9120 1050 9130 1060
rect 9250 1050 9260 1060
rect 9360 1050 9370 1060
rect 9900 1050 9920 1060
rect 740 1040 750 1050
rect 810 1040 860 1050
rect 1480 1040 1490 1050
rect 1520 1040 1650 1050
rect 2010 1040 2070 1050
rect 2220 1040 2840 1050
rect 3750 1040 3840 1050
rect 4050 1040 4060 1050
rect 4220 1040 4230 1050
rect 4560 1040 4570 1050
rect 5470 1040 5500 1050
rect 5630 1040 5640 1050
rect 5670 1040 5680 1050
rect 5700 1040 5720 1050
rect 5770 1040 5780 1050
rect 5820 1040 5880 1050
rect 5940 1040 5950 1050
rect 6440 1040 6470 1050
rect 6800 1040 6810 1050
rect 6830 1040 6840 1050
rect 7390 1040 7420 1050
rect 7920 1040 7970 1050
rect 8150 1040 8170 1050
rect 8180 1040 8380 1050
rect 8480 1040 8490 1050
rect 8500 1040 8510 1050
rect 8550 1040 8640 1050
rect 8650 1040 9100 1050
rect 9370 1040 9380 1050
rect 9900 1040 9910 1050
rect 9930 1040 9940 1050
rect 9970 1040 9990 1050
rect 810 1030 850 1040
rect 1470 1030 1480 1040
rect 1520 1030 1650 1040
rect 2010 1030 2060 1040
rect 2210 1030 2840 1040
rect 3730 1030 3850 1040
rect 4590 1030 4600 1040
rect 5420 1030 5430 1040
rect 5490 1030 5510 1040
rect 5520 1030 5550 1040
rect 5590 1030 5600 1040
rect 5670 1030 5680 1040
rect 5700 1030 5710 1040
rect 5820 1030 5840 1040
rect 5860 1030 5880 1040
rect 6430 1030 6450 1040
rect 6830 1030 6840 1040
rect 7390 1030 7430 1040
rect 7920 1030 7970 1040
rect 8140 1030 8160 1040
rect 8180 1030 8370 1040
rect 8480 1030 8490 1040
rect 8550 1030 8630 1040
rect 8650 1030 9110 1040
rect 9240 1030 9250 1040
rect 9720 1030 9730 1040
rect 9850 1030 9870 1040
rect 9920 1030 9930 1040
rect 9970 1030 9980 1040
rect 800 1020 840 1030
rect 1460 1020 1470 1030
rect 1510 1020 1610 1030
rect 1640 1020 1650 1030
rect 2010 1020 2050 1030
rect 2220 1020 2250 1030
rect 2260 1020 2840 1030
rect 3700 1020 3710 1030
rect 3730 1020 3850 1030
rect 4620 1020 4630 1030
rect 5490 1020 5550 1030
rect 5570 1020 5610 1030
rect 5620 1020 5640 1030
rect 5670 1020 5680 1030
rect 5700 1020 5710 1030
rect 5790 1020 5810 1030
rect 5980 1020 6000 1030
rect 6410 1020 6450 1030
rect 6830 1020 6840 1030
rect 7390 1020 7430 1030
rect 7930 1020 7970 1030
rect 8140 1020 8150 1030
rect 8180 1020 8350 1030
rect 8480 1020 8490 1030
rect 8550 1020 8630 1030
rect 8650 1020 9060 1030
rect 9070 1020 9100 1030
rect 9940 1020 9950 1030
rect 730 1010 740 1020
rect 800 1010 840 1020
rect 1490 1010 1600 1020
rect 2000 1010 2040 1020
rect 2230 1010 2240 1020
rect 2280 1010 2840 1020
rect 3710 1010 3720 1020
rect 3730 1010 3840 1020
rect 5490 1010 5530 1020
rect 5570 1010 5590 1020
rect 5600 1010 5640 1020
rect 5700 1010 5710 1020
rect 5840 1010 5850 1020
rect 5980 1010 5990 1020
rect 6400 1010 6450 1020
rect 6830 1010 6840 1020
rect 7390 1010 7430 1020
rect 7930 1010 7970 1020
rect 8140 1010 8150 1020
rect 8180 1010 8350 1020
rect 8520 1010 8550 1020
rect 8560 1010 8590 1020
rect 8650 1010 9000 1020
rect 9020 1010 9050 1020
rect 9070 1010 9100 1020
rect 9140 1010 9150 1020
rect 9380 1010 9390 1020
rect 9540 1010 9550 1020
rect 9930 1010 9960 1020
rect 800 1000 830 1010
rect 1440 1000 1450 1010
rect 1490 1000 1580 1010
rect 2000 1000 2030 1010
rect 2040 1000 2050 1010
rect 2290 1000 2840 1010
rect 3720 1000 3730 1010
rect 3740 1000 3830 1010
rect 4110 1000 4120 1010
rect 4210 1000 4220 1010
rect 4680 1000 4690 1010
rect 5380 1000 5390 1010
rect 5470 1000 5530 1010
rect 5620 1000 5630 1010
rect 5670 1000 5680 1010
rect 5700 1000 5710 1010
rect 5850 1000 5860 1010
rect 6280 1000 6290 1010
rect 6410 1000 6460 1010
rect 6830 1000 6840 1010
rect 7400 1000 7430 1010
rect 7930 1000 7970 1010
rect 8140 1000 8150 1010
rect 8190 1000 8340 1010
rect 8500 1000 8530 1010
rect 8540 1000 8550 1010
rect 8560 1000 8600 1010
rect 8660 1000 8990 1010
rect 9030 1000 9050 1010
rect 9070 1000 9100 1010
rect 9140 1000 9150 1010
rect 9400 1000 9410 1010
rect 9500 1000 9510 1010
rect 9930 1000 9960 1010
rect 790 990 820 1000
rect 1480 990 1560 1000
rect 2000 990 2040 1000
rect 2300 990 2460 1000
rect 2480 990 2590 1000
rect 2620 990 2670 1000
rect 2730 990 2820 1000
rect 2830 990 2840 1000
rect 3730 990 3740 1000
rect 3750 990 3830 1000
rect 4130 990 4140 1000
rect 4700 990 4710 1000
rect 5400 990 5420 1000
rect 5450 990 5520 1000
rect 5580 990 5610 1000
rect 5670 990 5680 1000
rect 5700 990 5710 1000
rect 5870 990 5890 1000
rect 5900 990 5910 1000
rect 5920 990 5930 1000
rect 6000 990 6010 1000
rect 6410 990 6460 1000
rect 6810 990 6820 1000
rect 6830 990 6840 1000
rect 7400 990 7430 1000
rect 7930 990 7970 1000
rect 8140 990 8150 1000
rect 8180 990 8340 1000
rect 8360 990 8370 1000
rect 8570 990 8970 1000
rect 9030 990 9040 1000
rect 9080 990 9110 1000
rect 9410 990 9420 1000
rect 790 980 820 990
rect 1470 980 1550 990
rect 2000 980 2030 990
rect 2300 980 2340 990
rect 2390 980 2420 990
rect 2530 980 2560 990
rect 2660 980 2670 990
rect 2740 980 2830 990
rect 3760 980 3820 990
rect 4150 980 4160 990
rect 4190 980 4200 990
rect 4730 980 4740 990
rect 5400 980 5430 990
rect 5450 980 5490 990
rect 5580 980 5640 990
rect 5670 980 5680 990
rect 5700 980 5720 990
rect 5730 980 5740 990
rect 5870 980 5890 990
rect 5900 980 5920 990
rect 6290 980 6300 990
rect 6400 980 6460 990
rect 6810 980 6820 990
rect 6830 980 6840 990
rect 7400 980 7430 990
rect 7940 980 7970 990
rect 8140 980 8150 990
rect 8180 980 8370 990
rect 8560 980 8960 990
rect 9020 980 9040 990
rect 9080 980 9110 990
rect 9750 980 9760 990
rect 9790 980 9830 990
rect 780 970 820 980
rect 1460 970 1540 980
rect 2000 970 2040 980
rect 2740 970 2820 980
rect 3750 970 3760 980
rect 3780 970 3830 980
rect 4750 970 4760 980
rect 5400 970 5470 980
rect 5520 970 5530 980
rect 5560 970 5680 980
rect 5700 970 5720 980
rect 5730 970 5760 980
rect 5850 970 5860 980
rect 5870 970 5920 980
rect 6280 970 6290 980
rect 6400 970 6460 980
rect 6810 970 6820 980
rect 7400 970 7430 980
rect 7940 970 7970 980
rect 8130 970 8150 980
rect 8190 970 8370 980
rect 8570 970 8950 980
rect 9080 970 9100 980
rect 9150 970 9160 980
rect 9520 970 9530 980
rect 9830 970 9840 980
rect 710 960 720 970
rect 780 960 810 970
rect 1460 960 1520 970
rect 2000 960 2030 970
rect 2720 960 2820 970
rect 3800 960 3830 970
rect 4760 960 4770 970
rect 5210 960 5220 970
rect 5300 960 5320 970
rect 5330 960 5380 970
rect 5390 960 5540 970
rect 5550 960 5610 970
rect 5620 960 5640 970
rect 5660 960 5680 970
rect 5720 960 5730 970
rect 5760 960 5800 970
rect 5810 960 5880 970
rect 5990 960 6000 970
rect 6270 960 6300 970
rect 6410 960 6470 970
rect 7390 960 7430 970
rect 7940 960 7970 970
rect 8130 960 8150 970
rect 8190 960 8360 970
rect 8560 960 8950 970
rect 9070 960 9110 970
rect 9750 960 9760 970
rect 9820 960 9830 970
rect 780 950 810 960
rect 1380 950 1390 960
rect 1440 950 1520 960
rect 2000 950 2030 960
rect 2730 950 2820 960
rect 3770 950 3780 960
rect 3790 950 3830 960
rect 4780 950 4790 960
rect 4820 950 4860 960
rect 5220 950 5230 960
rect 5300 950 5320 960
rect 5330 950 5380 960
rect 5400 950 5410 960
rect 5420 950 5430 960
rect 5440 950 5460 960
rect 5480 950 5500 960
rect 5540 950 5550 960
rect 5560 950 5600 960
rect 5630 950 5640 960
rect 5650 950 5680 960
rect 5710 950 5730 960
rect 5740 950 5750 960
rect 5760 950 5770 960
rect 5810 950 5840 960
rect 5850 950 5880 960
rect 5890 950 5970 960
rect 6020 950 6040 960
rect 6270 950 6300 960
rect 6410 950 6470 960
rect 7390 950 7430 960
rect 7940 950 7970 960
rect 8130 950 8140 960
rect 8190 950 8370 960
rect 8540 950 8550 960
rect 8570 950 8940 960
rect 9070 950 9110 960
rect 9750 950 9760 960
rect 780 940 810 950
rect 1420 940 1510 950
rect 2000 940 2030 950
rect 2730 940 2810 950
rect 3780 940 3790 950
rect 4800 940 4840 950
rect 5240 940 5290 950
rect 5310 940 5320 950
rect 5360 940 5370 950
rect 5400 940 5410 950
rect 5450 940 5460 950
rect 5490 940 5500 950
rect 5510 940 5530 950
rect 5540 940 5550 950
rect 5580 940 5590 950
rect 5610 940 5620 950
rect 5630 940 5640 950
rect 5660 940 5690 950
rect 5700 940 5710 950
rect 5720 940 5730 950
rect 5740 940 5750 950
rect 5760 940 5770 950
rect 5780 940 5800 950
rect 5810 940 5870 950
rect 5890 940 5960 950
rect 6030 940 6040 950
rect 6230 940 6240 950
rect 6250 940 6300 950
rect 6410 940 6470 950
rect 7390 940 7430 950
rect 7940 940 7980 950
rect 8120 940 8140 950
rect 8190 940 8370 950
rect 8570 940 8940 950
rect 9070 940 9110 950
rect 770 930 810 940
rect 1410 930 1500 940
rect 2000 930 2030 940
rect 2730 930 2790 940
rect 5250 930 5270 940
rect 5380 930 5410 940
rect 5450 930 5460 940
rect 5470 930 5500 940
rect 5510 930 5530 940
rect 5540 930 5550 940
rect 5560 930 5590 940
rect 5600 930 5620 940
rect 5630 930 5640 940
rect 5670 930 5680 940
rect 5690 930 5710 940
rect 5720 930 5730 940
rect 5740 930 5750 940
rect 5760 930 5780 940
rect 5790 930 5800 940
rect 5810 930 5860 940
rect 5870 930 6020 940
rect 6220 930 6300 940
rect 6420 930 6470 940
rect 6820 930 6850 940
rect 7390 930 7430 940
rect 7950 930 7980 940
rect 8130 930 8140 940
rect 8200 930 8370 940
rect 8420 930 8430 940
rect 8580 930 8930 940
rect 9070 930 9110 940
rect 9460 930 9470 940
rect 780 920 810 930
rect 1340 920 1350 930
rect 1400 920 1480 930
rect 2000 920 2030 930
rect 2730 920 2790 930
rect 3800 920 3810 930
rect 5360 920 5370 930
rect 5390 920 5410 930
rect 5450 920 5460 930
rect 5470 920 5500 930
rect 5510 920 5530 930
rect 5560 920 5580 930
rect 5600 920 5610 930
rect 5630 920 5660 930
rect 5670 920 5690 930
rect 5700 920 5730 930
rect 5740 920 5750 930
rect 5760 920 5780 930
rect 5790 920 5800 930
rect 5810 920 5860 930
rect 5870 920 6020 930
rect 6220 920 6300 930
rect 6420 920 6470 930
rect 6820 920 6850 930
rect 7390 920 7430 930
rect 7950 920 7980 930
rect 8130 920 8150 930
rect 8200 920 8380 930
rect 8400 920 8410 930
rect 8420 920 8430 930
rect 8580 920 8720 930
rect 8740 920 8930 930
rect 9080 920 9110 930
rect 9490 920 9500 930
rect 690 910 700 920
rect 770 910 810 920
rect 1390 910 1470 920
rect 2000 910 2030 920
rect 2720 910 2770 920
rect 4830 910 4840 920
rect 5330 910 5340 920
rect 5350 910 5370 920
rect 5400 910 5410 920
rect 5450 910 5460 920
rect 5510 910 5530 920
rect 5560 910 5590 920
rect 5600 910 5610 920
rect 5620 910 5660 920
rect 5700 910 5710 920
rect 5720 910 5730 920
rect 5760 910 5780 920
rect 5790 910 5850 920
rect 5860 910 6020 920
rect 6030 910 6040 920
rect 6220 910 6290 920
rect 6420 910 6470 920
rect 6820 910 6830 920
rect 6840 910 6850 920
rect 7390 910 7420 920
rect 7960 910 7980 920
rect 8130 910 8150 920
rect 8200 910 8400 920
rect 8520 910 8540 920
rect 8590 910 8710 920
rect 8750 910 8910 920
rect 9080 910 9100 920
rect 9110 910 9120 920
rect 9450 910 9460 920
rect 770 900 810 910
rect 1390 900 1450 910
rect 2000 900 2030 910
rect 2710 900 2760 910
rect 5270 900 5300 910
rect 5330 900 5340 910
rect 5350 900 5370 910
rect 5390 900 5400 910
rect 5450 900 5460 910
rect 5470 900 5480 910
rect 5490 900 5500 910
rect 5510 900 5530 910
rect 5540 900 5550 910
rect 5560 900 5570 910
rect 5580 900 5610 910
rect 5620 900 5640 910
rect 5670 900 5680 910
rect 5720 900 5770 910
rect 5780 900 5790 910
rect 5810 900 5850 910
rect 5860 900 6040 910
rect 6230 900 6290 910
rect 6420 900 6470 910
rect 6840 900 6850 910
rect 7380 900 7430 910
rect 7960 900 7980 910
rect 8130 900 8150 910
rect 8200 900 8410 910
rect 8430 900 8440 910
rect 8590 900 8710 910
rect 8720 900 8900 910
rect 9090 900 9100 910
rect 9110 900 9120 910
rect 9480 900 9490 910
rect 770 890 810 900
rect 840 890 880 900
rect 890 890 910 900
rect 1380 890 1440 900
rect 2000 890 2030 900
rect 2710 890 2750 900
rect 5290 890 5300 900
rect 5330 890 5340 900
rect 5350 890 5370 900
rect 5390 890 5400 900
rect 5450 890 5460 900
rect 5470 890 5480 900
rect 5490 890 5500 900
rect 5520 890 5530 900
rect 5540 890 5550 900
rect 5560 890 5600 900
rect 5630 890 5650 900
rect 5660 890 5680 900
rect 5700 890 5750 900
rect 5780 890 5790 900
rect 5810 890 5910 900
rect 5930 890 6000 900
rect 6010 890 6040 900
rect 6220 890 6290 900
rect 6410 890 6470 900
rect 6840 890 6850 900
rect 7380 890 7420 900
rect 7960 890 7990 900
rect 8130 890 8150 900
rect 8210 890 8430 900
rect 8610 890 8700 900
rect 8720 890 8890 900
rect 9080 890 9100 900
rect 9110 890 9120 900
rect 9540 890 9550 900
rect 770 880 920 890
rect 1290 880 1300 890
rect 1380 880 1420 890
rect 2010 880 2040 890
rect 2700 880 2730 890
rect 4850 880 4860 890
rect 5330 880 5340 890
rect 5360 880 5380 890
rect 5400 880 5410 890
rect 5430 880 5440 890
rect 5450 880 5460 890
rect 5490 880 5530 890
rect 5540 880 5570 890
rect 5580 880 5610 890
rect 5620 880 5680 890
rect 5700 880 5730 890
rect 5810 880 5970 890
rect 5980 880 6050 890
rect 6220 880 6280 890
rect 6420 880 6470 890
rect 6830 880 6850 890
rect 7380 880 7420 890
rect 7960 880 7990 890
rect 8130 880 8150 890
rect 8210 880 8430 890
rect 8650 880 8680 890
rect 8720 880 8870 890
rect 9070 880 9120 890
rect 9430 880 9440 890
rect 9530 880 9560 890
rect 760 870 920 880
rect 1280 870 1290 880
rect 1370 870 1410 880
rect 2010 870 2040 880
rect 2690 870 2720 880
rect 5360 870 5380 880
rect 5400 870 5420 880
rect 5430 870 5440 880
rect 5450 870 5470 880
rect 5480 870 5520 880
rect 5540 870 5570 880
rect 5600 870 5630 880
rect 5660 870 5680 880
rect 5700 870 5710 880
rect 5790 870 5800 880
rect 5810 870 6010 880
rect 6020 870 6050 880
rect 6210 870 6290 880
rect 6420 870 6480 880
rect 6830 870 6860 880
rect 7380 870 7430 880
rect 7960 870 7990 880
rect 8140 870 8150 880
rect 8200 870 8430 880
rect 8640 870 8680 880
rect 8710 870 8870 880
rect 9070 870 9100 880
rect 9110 870 9120 880
rect 9530 870 9550 880
rect 670 860 680 870
rect 760 860 920 870
rect 1360 860 1410 870
rect 2010 860 2040 870
rect 2680 860 2700 870
rect 4570 860 4600 870
rect 5350 860 5430 870
rect 5670 860 5680 870
rect 5700 860 5710 870
rect 5820 860 5960 870
rect 5970 860 6010 870
rect 6020 860 6030 870
rect 6220 860 6290 870
rect 6420 860 6470 870
rect 6840 860 6860 870
rect 7380 860 7420 870
rect 7960 860 7990 870
rect 8140 860 8150 870
rect 8200 860 8450 870
rect 8640 860 8870 870
rect 9070 860 9110 870
rect 9460 860 9470 870
rect 9530 860 9540 870
rect 9560 860 9590 870
rect 760 850 910 860
rect 1250 850 1260 860
rect 1340 850 1410 860
rect 2020 850 2050 860
rect 2660 850 2680 860
rect 4970 850 4980 860
rect 5060 850 5070 860
rect 5370 850 5440 860
rect 5700 850 5710 860
rect 5820 850 5960 860
rect 5980 850 6030 860
rect 6220 850 6280 860
rect 6440 850 6480 860
rect 6840 850 6860 860
rect 7380 850 7420 860
rect 7950 850 7990 860
rect 8140 850 8150 860
rect 8210 850 8460 860
rect 8640 850 8860 860
rect 9080 850 9110 860
rect 9180 850 9190 860
rect 760 840 910 850
rect 1240 840 1250 850
rect 1330 840 1400 850
rect 2020 840 2040 850
rect 2650 840 2660 850
rect 4260 840 4270 850
rect 5370 840 5410 850
rect 5470 840 5490 850
rect 5700 840 5710 850
rect 5770 840 5780 850
rect 5790 840 5820 850
rect 5830 840 5840 850
rect 5860 840 5880 850
rect 5890 840 5920 850
rect 5950 840 6010 850
rect 6210 840 6280 850
rect 6440 840 6480 850
rect 6840 840 6860 850
rect 7370 840 7420 850
rect 7960 840 7990 850
rect 8140 840 8150 850
rect 8220 840 8480 850
rect 8520 840 8530 850
rect 8630 840 8860 850
rect 9080 840 9110 850
rect 760 830 910 840
rect 1230 830 1240 840
rect 1330 830 1400 840
rect 2030 830 2040 840
rect 3970 830 4010 840
rect 4260 830 4280 840
rect 4880 830 4890 840
rect 5250 830 5270 840
rect 5380 830 5430 840
rect 5460 830 5520 840
rect 5530 830 5570 840
rect 5670 830 5680 840
rect 5700 830 5710 840
rect 5760 830 5880 840
rect 5890 830 6000 840
rect 6150 830 6160 840
rect 6200 830 6280 840
rect 6450 830 6480 840
rect 6840 830 6860 840
rect 7370 830 7420 840
rect 7960 830 7990 840
rect 8220 830 8480 840
rect 8520 830 8530 840
rect 8630 830 8850 840
rect 9080 830 9110 840
rect 9440 830 9450 840
rect 660 820 670 830
rect 760 820 880 830
rect 1210 820 1220 830
rect 1310 820 1390 830
rect 2030 820 2040 830
rect 3960 820 4020 830
rect 4270 820 4290 830
rect 5270 820 5280 830
rect 5380 820 5400 830
rect 5420 820 5430 830
rect 5470 820 5480 830
rect 5490 820 5510 830
rect 5560 820 5590 830
rect 5600 820 5680 830
rect 5700 820 5710 830
rect 5770 820 5880 830
rect 5890 820 6020 830
rect 6190 820 6290 830
rect 6450 820 6500 830
rect 6840 820 6860 830
rect 7370 820 7410 830
rect 7960 820 7990 830
rect 8220 820 8540 830
rect 8620 820 8850 830
rect 9080 820 9110 830
rect 760 810 860 820
rect 1200 810 1210 820
rect 1310 810 1380 820
rect 2040 810 2050 820
rect 3950 810 4020 820
rect 4280 810 4300 820
rect 5170 810 5190 820
rect 5280 810 5300 820
rect 5390 810 5420 820
rect 5670 810 5680 820
rect 5770 810 5880 820
rect 5900 810 6050 820
rect 6190 810 6290 820
rect 6460 810 6500 820
rect 6840 810 6860 820
rect 7370 810 7420 820
rect 7970 810 7990 820
rect 8230 810 8550 820
rect 8620 810 8840 820
rect 9080 810 9110 820
rect 9390 810 9400 820
rect 9430 810 9440 820
rect 9820 810 9850 820
rect 9910 810 9920 820
rect 750 800 850 810
rect 1260 800 1360 810
rect 2040 800 2060 810
rect 3920 800 3930 810
rect 3960 800 4020 810
rect 4290 800 4300 810
rect 5300 800 5310 810
rect 5400 800 5420 810
rect 5440 800 5460 810
rect 5470 800 5490 810
rect 5530 800 5550 810
rect 5670 800 5680 810
rect 5780 800 5790 810
rect 5850 800 6040 810
rect 6190 800 6290 810
rect 6460 800 6500 810
rect 6840 800 6860 810
rect 7370 800 7420 810
rect 7970 800 8000 810
rect 8130 800 8140 810
rect 8230 800 8610 810
rect 8630 800 8830 810
rect 9090 800 9100 810
rect 9890 800 9900 810
rect 740 790 830 800
rect 1170 790 1180 800
rect 1240 790 1340 800
rect 2040 790 2060 800
rect 3960 790 4020 800
rect 4300 790 4320 800
rect 4900 790 4910 800
rect 5220 790 5240 800
rect 5310 790 5320 800
rect 5410 790 5430 800
rect 5450 790 5550 800
rect 5700 790 5710 800
rect 5780 790 5790 800
rect 5800 790 5810 800
rect 5820 790 6040 800
rect 6060 790 6070 800
rect 6150 790 6160 800
rect 6190 790 6290 800
rect 6460 790 6510 800
rect 6840 790 6850 800
rect 6860 790 6870 800
rect 7370 790 7410 800
rect 7970 790 8000 800
rect 8230 790 8830 800
rect 9090 790 9100 800
rect 9380 790 9390 800
rect 740 780 820 790
rect 1240 780 1320 790
rect 2040 780 2070 790
rect 2540 780 2550 790
rect 3950 780 3960 790
rect 3980 780 4010 790
rect 4310 780 4320 790
rect 5220 780 5250 790
rect 5320 780 5330 790
rect 5490 780 5520 790
rect 5790 780 5970 790
rect 5980 780 6060 790
rect 6080 780 6090 790
rect 6160 780 6290 790
rect 6460 780 6520 790
rect 6840 780 6850 790
rect 6860 780 6870 790
rect 7360 780 7410 790
rect 7970 780 8000 790
rect 8230 780 8830 790
rect 9090 780 9100 790
rect 730 770 800 780
rect 1140 770 1160 780
rect 1240 770 1310 780
rect 2050 770 2070 780
rect 3670 770 3680 780
rect 3700 770 3730 780
rect 3990 770 4000 780
rect 4320 770 4330 780
rect 4340 770 4350 780
rect 5230 770 5250 780
rect 5420 770 5440 780
rect 5490 770 5520 780
rect 5770 770 5870 780
rect 5880 770 5960 780
rect 5970 770 6090 780
rect 6110 770 6120 780
rect 6180 770 6290 780
rect 6470 770 6510 780
rect 6520 770 6530 780
rect 6860 770 6870 780
rect 7360 770 7420 780
rect 7980 770 8000 780
rect 8130 770 8140 780
rect 8240 770 8810 780
rect 9090 770 9100 780
rect 9370 770 9380 780
rect 640 760 650 770
rect 720 760 780 770
rect 1130 760 1140 770
rect 1240 760 1280 770
rect 2050 760 2070 770
rect 3590 760 3650 770
rect 3670 760 3690 770
rect 3770 760 3790 770
rect 3840 760 3850 770
rect 5280 760 5290 770
rect 5430 760 5440 770
rect 5490 760 5520 770
rect 5700 760 5710 770
rect 5770 760 6040 770
rect 6050 760 6160 770
rect 6170 760 6300 770
rect 6480 760 6530 770
rect 6860 760 6870 770
rect 7360 760 7400 770
rect 7980 760 8010 770
rect 8250 760 8800 770
rect 9080 760 9100 770
rect 720 750 770 760
rect 1120 750 1130 760
rect 1250 750 1290 760
rect 2060 750 2070 760
rect 3540 750 3570 760
rect 3990 750 4000 760
rect 4340 750 4350 760
rect 4910 750 4920 760
rect 5450 750 5460 760
rect 5510 750 5530 760
rect 5770 750 6290 760
rect 6490 750 6530 760
rect 6860 750 6870 760
rect 7360 750 7400 760
rect 7980 750 8010 760
rect 8130 750 8140 760
rect 8250 750 8790 760
rect 9090 750 9110 760
rect 9460 750 9480 760
rect 720 740 760 750
rect 1100 740 1110 750
rect 1240 740 1290 750
rect 2070 740 2080 750
rect 3520 740 3530 750
rect 4910 740 4920 750
rect 5550 740 5560 750
rect 5570 740 5580 750
rect 5770 740 6300 750
rect 6490 740 6530 750
rect 6860 740 6870 750
rect 7360 740 7400 750
rect 7980 740 8010 750
rect 8130 740 8140 750
rect 8250 740 8780 750
rect 9080 740 9100 750
rect 9120 740 9130 750
rect 630 730 640 740
rect 710 730 750 740
rect 1090 730 1100 740
rect 1220 730 1290 740
rect 2070 730 2080 740
rect 3430 730 3510 740
rect 5510 730 5520 740
rect 5740 730 5750 740
rect 5760 730 5850 740
rect 5860 730 6020 740
rect 6040 730 6110 740
rect 6120 730 6300 740
rect 6490 730 6540 740
rect 6860 730 6870 740
rect 7360 730 7400 740
rect 7980 730 8010 740
rect 8130 730 8140 740
rect 8240 730 8770 740
rect 9080 730 9100 740
rect 9690 730 9720 740
rect 710 720 750 730
rect 1080 720 1090 730
rect 1220 720 1290 730
rect 2070 720 2090 730
rect 2440 720 2450 730
rect 3400 720 3420 730
rect 3910 720 3920 730
rect 4780 720 4800 730
rect 5370 720 5380 730
rect 5500 720 5520 730
rect 5640 720 5650 730
rect 5740 720 5760 730
rect 5770 720 5810 730
rect 5820 720 5830 730
rect 5840 720 5980 730
rect 6010 720 6050 730
rect 6060 720 6290 730
rect 6490 720 6540 730
rect 6870 720 6880 730
rect 7360 720 7410 730
rect 7990 720 8020 730
rect 8130 720 8140 730
rect 8230 720 8780 730
rect 9080 720 9100 730
rect 9340 720 9350 730
rect 9380 720 9390 730
rect 700 710 740 720
rect 1060 710 1090 720
rect 1210 710 1300 720
rect 2080 710 2090 720
rect 2420 710 2430 720
rect 4770 710 4790 720
rect 5380 710 5390 720
rect 5490 710 5500 720
rect 5780 710 5970 720
rect 6000 710 6290 720
rect 6490 710 6550 720
rect 6850 710 6860 720
rect 6870 710 6880 720
rect 7350 710 7400 720
rect 7990 710 8020 720
rect 8130 710 8140 720
rect 8250 710 8770 720
rect 9080 710 9100 720
rect 9210 710 9220 720
rect 700 700 730 710
rect 1050 700 1080 710
rect 1210 700 1300 710
rect 2080 700 2100 710
rect 3370 700 3380 710
rect 4160 700 4170 710
rect 4750 700 4790 710
rect 5490 700 5500 710
rect 5510 700 5520 710
rect 5670 700 5680 710
rect 5780 700 5880 710
rect 5890 700 5940 710
rect 5950 700 6290 710
rect 6510 700 6550 710
rect 6870 700 6880 710
rect 7350 700 7400 710
rect 7990 700 8020 710
rect 8130 700 8140 710
rect 8260 700 8770 710
rect 9080 700 9100 710
rect 9110 700 9120 710
rect 9330 700 9340 710
rect 9370 700 9380 710
rect 690 690 730 700
rect 1030 690 1070 700
rect 1210 690 1300 700
rect 2080 690 2100 700
rect 3350 690 3360 700
rect 4130 690 4180 700
rect 4710 690 4770 700
rect 4780 690 4800 700
rect 5500 690 5530 700
rect 5580 690 5590 700
rect 5620 690 5630 700
rect 5650 690 5660 700
rect 5770 690 5780 700
rect 5810 690 5820 700
rect 5840 690 5990 700
rect 6000 690 6160 700
rect 6170 690 6290 700
rect 6520 690 6560 700
rect 7350 690 7400 700
rect 8000 690 8020 700
rect 8130 690 8140 700
rect 8260 690 8750 700
rect 9360 690 9370 700
rect 610 680 620 690
rect 690 680 720 690
rect 1020 680 1060 690
rect 1210 680 1300 690
rect 2090 680 2110 690
rect 2370 680 2380 690
rect 4110 680 4180 690
rect 4710 680 4720 690
rect 4770 680 4810 690
rect 5500 680 5540 690
rect 5550 680 5560 690
rect 5580 680 5610 690
rect 5620 680 5650 690
rect 5780 680 5800 690
rect 5810 680 6290 690
rect 6520 680 6560 690
rect 7340 680 7390 690
rect 8010 680 8030 690
rect 8130 680 8140 690
rect 8280 680 8750 690
rect 9210 680 9220 690
rect 9320 680 9330 690
rect 9690 680 9700 690
rect 690 670 730 680
rect 1010 670 1060 680
rect 1210 670 1300 680
rect 2100 670 2110 680
rect 3320 670 3330 680
rect 4100 670 4170 680
rect 4710 670 4720 680
rect 4770 670 4810 680
rect 5500 670 5540 680
rect 5550 670 5590 680
rect 5600 670 5660 680
rect 5670 670 5680 680
rect 5770 670 5800 680
rect 5810 670 5860 680
rect 5870 670 6290 680
rect 6520 670 6560 680
rect 6880 670 6890 680
rect 7340 670 7390 680
rect 8010 670 8040 680
rect 8130 670 8140 680
rect 8290 670 8740 680
rect 9210 670 9220 680
rect 9350 670 9360 680
rect 9690 670 9710 680
rect 600 660 610 670
rect 690 660 760 670
rect 910 660 930 670
rect 980 660 1040 670
rect 1210 660 1300 670
rect 2100 660 2120 670
rect 3300 660 3310 670
rect 4100 660 4140 670
rect 4710 660 4720 670
rect 4780 660 4820 670
rect 4850 660 4860 670
rect 4920 660 4930 670
rect 5410 660 5420 670
rect 5510 660 5560 670
rect 5570 660 5580 670
rect 5610 660 5680 670
rect 5760 660 5860 670
rect 5880 660 5920 670
rect 5930 660 6290 670
rect 6540 660 6570 670
rect 6860 660 6870 670
rect 6880 660 6890 670
rect 7340 660 7390 670
rect 8010 660 8040 670
rect 8130 660 8140 670
rect 8310 660 8740 670
rect 9340 660 9350 670
rect 9590 660 9600 670
rect 9610 660 9630 670
rect 9700 660 9720 670
rect 590 650 610 660
rect 690 650 820 660
rect 860 650 1050 660
rect 1200 650 1290 660
rect 2100 650 2120 660
rect 2320 650 2330 660
rect 3280 650 3300 660
rect 4090 650 4130 660
rect 4710 650 4720 660
rect 4780 650 4850 660
rect 5410 650 5430 660
rect 5520 650 5580 660
rect 5600 650 5660 660
rect 5670 650 5680 660
rect 5740 650 5780 660
rect 5810 650 6290 660
rect 6540 650 6580 660
rect 6860 650 6870 660
rect 6880 650 6890 660
rect 7340 650 7390 660
rect 8020 650 8050 660
rect 8120 650 8140 660
rect 8320 650 8730 660
rect 9070 650 9080 660
rect 9150 650 9160 660
rect 9620 650 9640 660
rect 9700 650 9730 660
rect 580 640 650 650
rect 670 640 680 650
rect 690 640 1010 650
rect 1030 640 1050 650
rect 1170 640 1290 650
rect 2110 640 2120 650
rect 3260 640 3280 650
rect 4080 640 4110 650
rect 4710 640 4720 650
rect 4830 640 4840 650
rect 5420 640 5430 650
rect 5540 640 5600 650
rect 5610 640 5690 650
rect 5750 640 5820 650
rect 5850 640 6280 650
rect 6530 640 6590 650
rect 6860 640 6870 650
rect 6880 640 6890 650
rect 7330 640 7380 650
rect 8020 640 8060 650
rect 8120 640 8140 650
rect 8330 640 8710 650
rect 9130 640 9140 650
rect 9330 640 9340 650
rect 9620 640 9640 650
rect 520 630 710 640
rect 760 630 980 640
rect 1100 630 1280 640
rect 3240 630 3270 640
rect 4090 630 4110 640
rect 4710 630 4720 640
rect 4810 630 4820 640
rect 5540 630 5590 640
rect 5600 630 5690 640
rect 5780 630 5820 640
rect 5850 630 6280 640
rect 6530 630 6590 640
rect 6880 630 6890 640
rect 7330 630 7380 640
rect 8020 630 8060 640
rect 8120 630 8140 640
rect 8340 630 8690 640
rect 8700 630 8710 640
rect 9130 630 9150 640
rect 9630 630 9640 640
rect 480 620 500 630
rect 610 620 700 630
rect 770 620 960 630
rect 1090 620 1280 630
rect 2120 620 2130 630
rect 2270 620 2280 630
rect 3220 620 3250 630
rect 4560 620 4570 630
rect 4710 620 4720 630
rect 4790 620 4800 630
rect 5550 620 5680 630
rect 5850 620 6290 630
rect 6540 620 6590 630
rect 6890 620 6900 630
rect 7320 620 7380 630
rect 8030 620 8070 630
rect 8110 620 8140 630
rect 8360 620 8690 630
rect 8700 620 8720 630
rect 9140 620 9150 630
rect 9200 620 9210 630
rect 9320 620 9330 630
rect 9630 620 9660 630
rect 9950 620 9980 630
rect 450 610 470 620
rect 630 610 700 620
rect 770 610 930 620
rect 940 610 950 620
rect 1060 610 1260 620
rect 2120 610 2140 620
rect 3150 610 3160 620
rect 3170 610 3210 620
rect 4050 610 4080 620
rect 4550 610 4570 620
rect 4710 610 4720 620
rect 4780 610 4790 620
rect 5560 610 5590 620
rect 5620 610 5630 620
rect 5640 610 5680 620
rect 5820 610 6300 620
rect 6540 610 6610 620
rect 6890 610 6900 620
rect 7310 610 7380 620
rect 8040 610 8090 620
rect 8110 610 8140 620
rect 8360 610 8700 620
rect 9140 610 9150 620
rect 9200 610 9210 620
rect 9220 610 9230 620
rect 9280 610 9290 620
rect 9300 610 9320 620
rect 420 600 430 610
rect 630 600 700 610
rect 770 600 930 610
rect 1060 600 1250 610
rect 1320 600 1390 610
rect 1400 600 1410 610
rect 2120 600 2150 610
rect 2240 600 2250 610
rect 4050 600 4080 610
rect 4550 600 4560 610
rect 4710 600 4720 610
rect 4770 600 4780 610
rect 5570 600 5680 610
rect 5850 600 6300 610
rect 6550 600 6610 610
rect 6870 600 6880 610
rect 6890 600 6910 610
rect 7310 600 7380 610
rect 8050 600 8100 610
rect 8110 600 8140 610
rect 8370 600 8670 610
rect 9120 600 9140 610
rect 9200 600 9210 610
rect 9300 600 9310 610
rect 9700 600 9710 610
rect 390 590 410 600
rect 640 590 710 600
rect 770 590 910 600
rect 920 590 930 600
rect 1060 590 1250 600
rect 1300 590 1420 600
rect 2120 590 2150 600
rect 2210 590 2230 600
rect 4540 590 4550 600
rect 4710 590 4720 600
rect 4760 590 4770 600
rect 5590 590 5680 600
rect 5850 590 6310 600
rect 6560 590 6620 600
rect 6890 590 6910 600
rect 7300 590 7380 600
rect 8060 590 8140 600
rect 8390 590 8650 600
rect 9050 590 9070 600
rect 9100 590 9110 600
rect 9220 590 9230 600
rect 9270 590 9280 600
rect 9300 590 9310 600
rect 9680 590 9700 600
rect 370 580 380 590
rect 650 580 720 590
rect 730 580 740 590
rect 750 580 910 590
rect 1050 580 1230 590
rect 1290 580 1400 590
rect 1420 580 1430 590
rect 2130 580 2160 590
rect 2180 580 2210 590
rect 4530 580 4550 590
rect 4690 580 4710 590
rect 4760 580 4770 590
rect 5590 580 5680 590
rect 5880 580 6320 590
rect 6570 580 6640 590
rect 6900 580 6910 590
rect 7300 580 7380 590
rect 8060 580 8140 590
rect 8400 580 8650 590
rect 9050 580 9090 590
rect 9130 580 9140 590
rect 9170 580 9200 590
rect 9220 580 9240 590
rect 9260 580 9270 590
rect 350 570 360 580
rect 650 570 910 580
rect 1050 570 1210 580
rect 1280 570 1310 580
rect 1320 570 1330 580
rect 1340 570 1380 580
rect 1430 570 1440 580
rect 2130 570 2170 580
rect 2190 570 2200 580
rect 3050 570 3110 580
rect 4080 570 4090 580
rect 4530 570 4540 580
rect 4690 570 4710 580
rect 4750 570 4760 580
rect 4940 570 4950 580
rect 5590 570 5600 580
rect 5610 570 5680 580
rect 5880 570 6320 580
rect 6570 570 6640 580
rect 6880 570 6890 580
rect 6900 570 6910 580
rect 7310 570 7370 580
rect 8070 570 8140 580
rect 8430 570 8570 580
rect 8590 570 8650 580
rect 9050 570 9090 580
rect 9100 570 9140 580
rect 9170 570 9220 580
rect 9230 570 9240 580
rect 9290 570 9300 580
rect 330 560 340 570
rect 650 560 920 570
rect 1050 560 1190 570
rect 1260 560 1280 570
rect 1440 560 1450 570
rect 2130 560 2180 570
rect 3030 560 3040 570
rect 4460 560 4470 570
rect 4510 560 4530 570
rect 4550 560 4560 570
rect 4670 560 4700 570
rect 4750 560 4770 570
rect 5610 560 5680 570
rect 5850 560 5910 570
rect 5930 560 6320 570
rect 6580 560 6650 570
rect 6880 560 6890 570
rect 6900 560 6910 570
rect 7300 560 7370 570
rect 8080 560 8130 570
rect 8440 560 8570 570
rect 8600 560 8610 570
rect 9040 560 9100 570
rect 9120 560 9140 570
rect 9170 560 9180 570
rect 9190 560 9230 570
rect 9250 560 9260 570
rect 310 550 330 560
rect 650 550 930 560
rect 1050 550 1160 560
rect 1250 550 1260 560
rect 1450 550 1460 560
rect 4430 550 4460 560
rect 4480 550 4510 560
rect 4670 550 4700 560
rect 4750 550 4770 560
rect 5630 550 5680 560
rect 5850 550 5880 560
rect 5910 550 5920 560
rect 5930 550 6320 560
rect 6580 550 6660 560
rect 6900 550 6910 560
rect 7310 550 7370 560
rect 8090 550 8110 560
rect 8440 550 8450 560
rect 8460 550 8470 560
rect 8480 550 8560 560
rect 9040 550 9100 560
rect 9180 550 9190 560
rect 9940 550 9960 560
rect 290 540 330 550
rect 650 540 930 550
rect 1050 540 1140 550
rect 1240 540 1250 550
rect 2990 540 3000 550
rect 4470 540 4500 550
rect 4540 540 4550 550
rect 4660 540 4680 550
rect 4750 540 4770 550
rect 5630 540 5680 550
rect 5840 540 5850 550
rect 5930 540 6320 550
rect 6580 540 6660 550
rect 6900 540 6930 550
rect 7300 540 7360 550
rect 8470 540 8500 550
rect 8520 540 8530 550
rect 9170 540 9190 550
rect 9960 540 9980 550
rect 260 530 340 540
rect 640 530 670 540
rect 700 530 940 540
rect 1050 530 1100 540
rect 1230 530 1240 540
rect 4450 530 4480 540
rect 4540 530 4550 540
rect 4650 530 4680 540
rect 4740 530 4770 540
rect 5630 530 5670 540
rect 5890 530 5900 540
rect 5930 530 5940 540
rect 5950 530 6000 540
rect 6010 530 6320 540
rect 6590 530 6660 540
rect 6890 530 6900 540
rect 6910 530 6920 540
rect 7300 530 7360 540
rect 9040 530 9060 540
rect 9170 530 9210 540
rect 9270 530 9280 540
rect 9990 530 9990 540
rect 230 520 340 530
rect 630 520 670 530
rect 710 520 750 530
rect 780 520 830 530
rect 870 520 950 530
rect 1040 520 1090 530
rect 1220 520 1230 530
rect 1490 520 1500 530
rect 2960 520 2970 530
rect 4360 520 4470 530
rect 4540 520 4560 530
rect 4640 520 4690 530
rect 4740 520 4770 530
rect 4950 520 4960 530
rect 5640 520 5670 530
rect 5970 520 6330 530
rect 6600 520 6660 530
rect 6890 520 6940 530
rect 7300 520 7370 530
rect 9040 520 9070 530
rect 9170 520 9210 530
rect 9940 520 9950 530
rect 210 510 320 520
rect 340 510 350 520
rect 580 510 660 520
rect 880 510 990 520
rect 1030 510 1090 520
rect 1210 510 1220 520
rect 2930 510 2950 520
rect 4280 510 4440 520
rect 4540 510 4610 520
rect 4630 510 4690 520
rect 4740 510 4760 520
rect 5650 510 5670 520
rect 5870 510 5890 520
rect 5930 510 6320 520
rect 6600 510 6660 520
rect 6900 510 6940 520
rect 7290 510 7360 520
rect 9050 510 9070 520
rect 9180 510 9190 520
rect 9220 510 9230 520
rect 9260 510 9270 520
rect 190 500 200 510
rect 250 500 320 510
rect 350 500 360 510
rect 530 500 660 510
rect 890 500 1090 510
rect 1190 500 1200 510
rect 1500 500 1510 510
rect 2880 500 2910 510
rect 4260 500 4410 510
rect 4540 500 4690 510
rect 4740 500 4770 510
rect 5660 500 5670 510
rect 5870 500 5880 510
rect 5930 500 5950 510
rect 5960 500 6310 510
rect 6610 500 6660 510
rect 6900 500 6940 510
rect 7280 500 7370 510
rect 9050 500 9070 510
rect 9140 500 9150 510
rect 9180 500 9190 510
rect 9910 500 9920 510
rect 170 490 180 500
rect 290 490 340 500
rect 360 490 370 500
rect 520 490 650 500
rect 900 490 1090 500
rect 1180 490 1190 500
rect 1490 490 1520 500
rect 2860 490 2870 500
rect 4260 490 4400 500
rect 4540 490 4690 500
rect 4740 490 4770 500
rect 5800 490 5820 500
rect 5850 490 5860 500
rect 5870 490 5900 500
rect 5920 490 6310 500
rect 6620 490 6670 500
rect 6900 490 6940 500
rect 7280 490 7350 500
rect 9130 490 9140 500
rect 9910 490 9920 500
rect 9980 490 9990 500
rect 310 480 350 490
rect 370 480 380 490
rect 500 480 650 490
rect 900 480 1090 490
rect 1490 480 1510 490
rect 2830 480 2850 490
rect 4250 480 4310 490
rect 4550 480 4690 490
rect 4740 480 4760 490
rect 5810 480 5830 490
rect 5880 480 5890 490
rect 5910 480 5920 490
rect 5940 480 6320 490
rect 6620 480 6690 490
rect 6910 480 6950 490
rect 7280 480 7350 490
rect 9060 480 9070 490
rect 9900 480 9910 490
rect 320 470 350 480
rect 380 470 390 480
rect 490 470 560 480
rect 650 470 660 480
rect 920 470 1090 480
rect 2790 470 2810 480
rect 4240 470 4260 480
rect 4280 470 4290 480
rect 4550 470 4690 480
rect 4740 470 4760 480
rect 5800 470 5840 480
rect 5940 470 6300 480
rect 6620 470 6700 480
rect 6910 470 6940 480
rect 7280 470 7350 480
rect 9060 470 9080 480
rect 9110 470 9130 480
rect 9200 470 9210 480
rect 9240 470 9250 480
rect 9850 470 9860 480
rect 9900 470 9910 480
rect 9920 470 9930 480
rect 330 460 360 470
rect 470 460 550 470
rect 640 460 670 470
rect 940 460 1080 470
rect 2120 460 2140 470
rect 2760 460 2780 470
rect 4230 460 4260 470
rect 4550 460 4690 470
rect 4740 460 4760 470
rect 4960 460 4970 470
rect 5810 460 5830 470
rect 5840 460 5860 470
rect 5940 460 5950 470
rect 5970 460 6290 470
rect 6620 460 6690 470
rect 6940 460 6950 470
rect 7280 460 7350 470
rect 9040 460 9080 470
rect 9090 460 9130 470
rect 9850 460 9860 470
rect 340 450 370 460
rect 470 450 550 460
rect 630 450 660 460
rect 950 450 1060 460
rect 2070 450 2080 460
rect 2190 450 2200 460
rect 2710 450 2730 460
rect 4220 450 4270 460
rect 4560 450 4690 460
rect 4740 450 4760 460
rect 4960 450 4970 460
rect 5810 450 5870 460
rect 5950 450 6270 460
rect 6630 450 6700 460
rect 7270 450 7350 460
rect 9050 450 9070 460
rect 9100 450 9110 460
rect 9190 450 9200 460
rect 9860 450 9870 460
rect 350 440 380 450
rect 410 440 420 450
rect 460 440 560 450
rect 630 440 670 450
rect 1010 440 1020 450
rect 1130 440 1140 450
rect 2250 440 2260 450
rect 2670 440 2690 450
rect 4210 440 4290 450
rect 4480 440 4490 450
rect 4570 440 4690 450
rect 4720 440 4750 450
rect 5810 440 5820 450
rect 5830 440 5870 450
rect 5950 440 6280 450
rect 6640 440 6700 450
rect 7260 440 7350 450
rect 9000 440 9020 450
rect 9050 440 9060 450
rect 9090 440 9120 450
rect 9130 440 9160 450
rect 9290 440 9320 450
rect 350 430 380 440
rect 410 430 420 440
rect 460 430 560 440
rect 610 430 670 440
rect 1120 430 1130 440
rect 2280 430 2290 440
rect 2640 430 2650 440
rect 4210 430 4290 440
rect 4480 430 4490 440
rect 4590 430 4630 440
rect 4720 430 4740 440
rect 5840 430 5860 440
rect 5970 430 6280 440
rect 6650 430 6720 440
rect 7250 430 7350 440
rect 8990 430 9010 440
rect 9020 430 9030 440
rect 9050 430 9060 440
rect 9080 430 9090 440
rect 9100 430 9150 440
rect 9210 430 9220 440
rect 9290 430 9330 440
rect 370 420 390 430
rect 420 420 430 430
rect 460 420 550 430
rect 560 420 570 430
rect 600 420 670 430
rect 1710 420 1720 430
rect 4200 420 4270 430
rect 4670 420 4680 430
rect 4720 420 4740 430
rect 5810 420 5860 430
rect 5980 420 6270 430
rect 6650 420 6720 430
rect 7240 420 7350 430
rect 8990 420 9020 430
rect 9030 420 9060 430
rect 9080 420 9090 430
rect 9130 420 9140 430
rect 9170 420 9180 430
rect 9290 420 9300 430
rect 370 410 400 420
rect 420 410 430 420
rect 470 410 560 420
rect 590 410 670 420
rect 2350 410 2360 420
rect 2520 410 2530 420
rect 4190 410 4260 420
rect 4480 410 4490 420
rect 4720 410 4740 420
rect 5820 410 5850 420
rect 5980 410 6270 420
rect 6670 410 6730 420
rect 7240 410 7350 420
rect 8990 410 9030 420
rect 9040 410 9090 420
rect 9130 410 9140 420
rect 9340 410 9390 420
rect 80 400 90 410
rect 380 400 400 410
rect 430 400 440 410
rect 480 400 560 410
rect 570 400 670 410
rect 4190 400 4250 410
rect 4340 400 4350 410
rect 4440 400 4450 410
rect 4460 400 4490 410
rect 4720 400 4730 410
rect 5990 400 6000 410
rect 6010 400 6280 410
rect 6680 400 6730 410
rect 7240 400 7340 410
rect 9010 400 9060 410
rect 9080 400 9090 410
rect 9120 400 9140 410
rect 9160 400 9170 410
rect 9330 400 9390 410
rect 390 390 400 400
rect 430 390 450 400
rect 470 390 670 400
rect 4190 390 4260 400
rect 4320 390 4360 400
rect 4460 390 4470 400
rect 4560 390 4570 400
rect 4720 390 4730 400
rect 6000 390 6270 400
rect 6690 390 6740 400
rect 7230 390 7330 400
rect 8980 390 9060 400
rect 9110 390 9130 400
rect 9320 390 9330 400
rect 9350 390 9380 400
rect 390 380 400 390
rect 440 380 450 390
rect 470 380 670 390
rect 4190 380 4250 390
rect 4310 380 4370 390
rect 4560 380 4580 390
rect 4720 380 4730 390
rect 6010 380 6290 390
rect 6700 380 6760 390
rect 7220 380 7330 390
rect 8970 380 9060 390
rect 9090 380 9120 390
rect 9260 380 9280 390
rect 9320 380 9330 390
rect 9390 380 9410 390
rect 9990 380 9990 390
rect 60 370 70 380
rect 390 370 410 380
rect 440 370 450 380
rect 480 370 670 380
rect 1080 370 1090 380
rect 1240 370 1250 380
rect 4190 370 4250 380
rect 4300 370 4380 380
rect 4550 370 4590 380
rect 4720 370 4730 380
rect 6000 370 6290 380
rect 6700 370 6770 380
rect 7220 370 7330 380
rect 8840 370 8860 380
rect 8980 370 9060 380
rect 9100 370 9110 380
rect 9180 370 9190 380
rect 9250 370 9320 380
rect 9400 370 9430 380
rect 380 360 410 370
rect 440 360 450 370
rect 470 360 560 370
rect 570 360 580 370
rect 600 360 610 370
rect 650 360 670 370
rect 1230 360 1250 370
rect 4190 360 4240 370
rect 4290 360 4300 370
rect 4320 360 4340 370
rect 4350 360 4390 370
rect 4550 360 4600 370
rect 4720 360 4740 370
rect 5810 360 5840 370
rect 6000 360 6280 370
rect 6710 360 6780 370
rect 7220 360 7330 370
rect 8830 360 8860 370
rect 8980 360 9000 370
rect 9030 360 9060 370
rect 9090 360 9110 370
rect 9140 360 9150 370
rect 9290 360 9310 370
rect 9320 360 9330 370
rect 9400 360 9430 370
rect 9970 360 9990 370
rect 50 350 60 360
rect 380 350 410 360
rect 460 350 530 360
rect 650 350 660 360
rect 4190 350 4230 360
rect 4240 350 4250 360
rect 4350 350 4400 360
rect 4560 350 4610 360
rect 4720 350 4740 360
rect 4970 350 4980 360
rect 5790 350 5840 360
rect 6010 350 6280 360
rect 6720 350 6780 360
rect 7210 350 7330 360
rect 8810 350 8850 360
rect 8980 350 9000 360
rect 9080 350 9110 360
rect 9240 350 9250 360
rect 9260 350 9290 360
rect 9310 350 9320 360
rect 9970 350 9980 360
rect 380 340 420 350
rect 450 340 510 350
rect 550 340 680 350
rect 4180 340 4260 350
rect 4270 340 4280 350
rect 4360 340 4470 350
rect 4510 340 4530 350
rect 4560 340 4620 350
rect 4690 340 4710 350
rect 4720 340 4740 350
rect 5800 340 5850 350
rect 6000 340 6280 350
rect 6720 340 6790 350
rect 7200 340 7330 350
rect 8800 340 8850 350
rect 8980 340 9020 350
rect 9160 340 9170 350
rect 9270 340 9300 350
rect 9420 340 9430 350
rect 9970 340 9990 350
rect 390 330 420 340
rect 450 330 530 340
rect 690 330 700 340
rect 1050 330 1060 340
rect 4170 330 4220 340
rect 4230 330 4250 340
rect 4360 330 4470 340
rect 4500 330 4540 340
rect 4570 330 4600 340
rect 4680 330 4750 340
rect 5820 330 5860 340
rect 6010 330 6270 340
rect 6740 330 6800 340
rect 7210 330 7320 340
rect 8800 330 8850 340
rect 8880 330 8900 340
rect 8990 330 9030 340
rect 9090 330 9100 340
rect 9150 330 9160 340
rect 9220 330 9230 340
rect 9280 330 9300 340
rect 9490 330 9500 340
rect 30 320 40 330
rect 390 320 420 330
rect 480 320 500 330
rect 700 320 730 330
rect 4220 320 4250 330
rect 4370 320 4480 330
rect 4490 320 4550 330
rect 4660 320 4750 330
rect 5680 320 5690 330
rect 5830 320 5860 330
rect 6010 320 6280 330
rect 6740 320 6820 330
rect 7170 320 7320 330
rect 8800 320 8810 330
rect 8880 320 8890 330
rect 9000 320 9040 330
rect 400 310 420 320
rect 470 310 480 320
rect 720 310 790 320
rect 4220 310 4240 320
rect 4390 310 4410 320
rect 4420 310 4430 320
rect 4460 310 4480 320
rect 4490 310 4500 320
rect 4530 310 4560 320
rect 4660 310 4750 320
rect 5850 310 5860 320
rect 6010 310 6260 320
rect 6750 310 6840 320
rect 7120 310 7320 320
rect 8940 310 8950 320
rect 9000 310 9030 320
rect 9140 310 9150 320
rect 9210 310 9220 320
rect 400 300 430 310
rect 790 300 820 310
rect 930 300 940 310
rect 4140 300 4150 310
rect 4180 300 4240 310
rect 4460 300 4490 310
rect 4530 300 4560 310
rect 4660 300 4740 310
rect 5800 300 5810 310
rect 6000 300 6270 310
rect 6770 300 6860 310
rect 7110 300 7320 310
rect 8900 300 8940 310
rect 9010 300 9050 310
rect 9070 300 9080 310
rect 9210 300 9220 310
rect 9410 300 9420 310
rect 20 290 30 300
rect 400 290 430 300
rect 820 290 990 300
rect 1030 290 1040 300
rect 4120 290 4230 300
rect 4470 290 4490 300
rect 4530 290 4560 300
rect 4650 290 4710 300
rect 5990 290 6280 300
rect 6780 290 6890 300
rect 7050 290 7080 300
rect 7090 290 7100 300
rect 7110 290 7320 300
rect 8900 290 8930 300
rect 9020 290 9050 300
rect 9060 290 9070 300
rect 9130 290 9140 300
rect 9420 290 9430 300
rect 9700 290 9720 300
rect 9750 290 9760 300
rect 20 280 30 290
rect 400 280 430 290
rect 650 280 680 290
rect 850 280 1010 290
rect 1030 280 1040 290
rect 4120 280 4220 290
rect 4470 280 4480 290
rect 4530 280 4570 290
rect 4590 280 4620 290
rect 4650 280 4680 290
rect 5990 280 6070 290
rect 6130 280 6270 290
rect 6790 280 6900 290
rect 6920 280 6930 290
rect 6970 280 7000 290
rect 7030 280 7050 290
rect 7060 280 7320 290
rect 8910 280 8930 290
rect 9030 280 9060 290
rect 9090 280 9100 290
rect 9210 280 9220 290
rect 9420 280 9440 290
rect 400 270 430 280
rect 440 270 450 280
rect 640 270 680 280
rect 860 270 1000 280
rect 1290 270 1300 280
rect 4110 270 4210 280
rect 4530 270 4570 280
rect 4590 270 4630 280
rect 4650 270 4670 280
rect 4980 270 4990 280
rect 5780 270 5790 280
rect 6000 270 6040 280
rect 6130 270 6280 280
rect 6790 270 6990 280
rect 7010 270 7050 280
rect 7070 270 7330 280
rect 8900 270 8930 280
rect 9050 270 9060 280
rect 9120 270 9130 280
rect 9200 270 9210 280
rect 9290 270 9310 280
rect 9430 270 9450 280
rect 9570 270 9580 280
rect 10 260 20 270
rect 400 260 420 270
rect 640 260 680 270
rect 870 260 1000 270
rect 1020 260 1030 270
rect 1280 260 1290 270
rect 4110 260 4200 270
rect 4540 260 4580 270
rect 4590 260 4630 270
rect 4650 260 4660 270
rect 6130 260 6280 270
rect 6810 260 6990 270
rect 7010 260 7050 270
rect 7060 260 7320 270
rect 8890 260 8930 270
rect 9080 260 9090 270
rect 9270 260 9300 270
rect 9390 260 9410 270
rect 9430 260 9440 270
rect 9990 260 9990 270
rect 10 250 20 260
rect 130 250 190 260
rect 390 250 420 260
rect 430 250 440 260
rect 630 250 680 260
rect 870 250 1010 260
rect 1020 250 1030 260
rect 1230 250 1240 260
rect 1270 250 1280 260
rect 4110 250 4190 260
rect 4540 250 4550 260
rect 4570 250 4580 260
rect 4590 250 4600 260
rect 4610 250 4660 260
rect 6130 250 6270 260
rect 6810 250 7330 260
rect 8880 250 8900 260
rect 8930 250 8940 260
rect 9110 250 9120 260
rect 9260 250 9280 260
rect 9340 250 9350 260
rect 9370 250 9390 260
rect 9430 250 9440 260
rect 10 240 20 250
rect 120 240 200 250
rect 380 240 410 250
rect 430 240 440 250
rect 630 240 680 250
rect 870 240 1020 250
rect 1230 240 1270 250
rect 4110 240 4180 250
rect 4540 240 4550 250
rect 4560 240 4580 250
rect 4590 240 4600 250
rect 4620 240 4660 250
rect 4840 240 4850 250
rect 6120 240 6280 250
rect 6830 240 7320 250
rect 8880 240 8890 250
rect 8950 240 8960 250
rect 9070 240 9080 250
rect 9170 240 9180 250
rect 9190 240 9200 250
rect 9240 240 9290 250
rect 9360 240 9380 250
rect 9410 240 9440 250
rect 9830 240 9850 250
rect 10 230 20 240
rect 120 230 210 240
rect 380 230 410 240
rect 420 230 430 240
rect 630 230 680 240
rect 870 230 1020 240
rect 4110 230 4170 240
rect 4210 230 4220 240
rect 4530 230 4550 240
rect 4570 230 4590 240
rect 4620 230 4660 240
rect 4840 230 4870 240
rect 4880 230 4890 240
rect 4990 230 5000 240
rect 6110 230 6290 240
rect 6830 230 6840 240
rect 6850 230 7320 240
rect 8870 230 8880 240
rect 9100 230 9110 240
rect 9190 230 9300 240
rect 9360 230 9400 240
rect 9430 230 9450 240
rect 9810 230 9830 240
rect 9840 230 9850 240
rect 90 220 210 230
rect 370 220 400 230
rect 420 220 430 230
rect 620 220 680 230
rect 870 220 1020 230
rect 4130 220 4160 230
rect 4200 220 4220 230
rect 4230 220 4240 230
rect 4540 220 4550 230
rect 4560 220 4590 230
rect 4630 220 4650 230
rect 4850 220 4890 230
rect 6110 220 6290 230
rect 6850 220 7320 230
rect 8870 220 8880 230
rect 8960 220 8970 230
rect 9160 220 9170 230
rect 9200 220 9300 230
rect 9370 220 9400 230
rect 9500 220 9510 230
rect 9790 220 9800 230
rect 9810 220 9820 230
rect 9830 220 9850 230
rect 60 210 160 220
rect 200 210 210 220
rect 360 210 400 220
rect 420 210 430 220
rect 620 210 680 220
rect 880 210 1020 220
rect 4130 210 4160 220
rect 4180 210 4250 220
rect 4330 210 4350 220
rect 4560 210 4590 220
rect 4630 210 4650 220
rect 4850 210 4880 220
rect 6110 210 6290 220
rect 6850 210 6860 220
rect 6870 210 7310 220
rect 8860 210 8880 220
rect 9160 210 9170 220
rect 9190 210 9310 220
rect 9360 210 9400 220
rect 9780 210 9810 220
rect 9840 210 9850 220
rect 9940 210 9950 220
rect 60 200 140 210
rect 210 200 220 210
rect 340 200 390 210
rect 420 200 430 210
rect 610 200 680 210
rect 860 200 1000 210
rect 1010 200 1020 210
rect 4150 200 4250 210
rect 4320 200 4380 210
rect 4520 200 4540 210
rect 4560 200 4590 210
rect 4630 200 4640 210
rect 6100 200 6300 210
rect 6880 200 7310 210
rect 8700 200 8710 210
rect 8860 200 8870 210
rect 8930 200 8940 210
rect 9080 200 9090 210
rect 9180 200 9240 210
rect 9280 200 9300 210
rect 9800 200 9810 210
rect 9840 200 9850 210
rect 9960 200 9970 210
rect 0 190 10 200
rect 70 190 110 200
rect 210 190 220 200
rect 330 190 380 200
rect 420 190 450 200
rect 610 190 690 200
rect 860 190 1020 200
rect 4150 190 4250 200
rect 4290 190 4400 200
rect 4420 190 4440 200
rect 4490 190 4540 200
rect 4560 190 4580 200
rect 6090 190 6310 200
rect 6900 190 6910 200
rect 6920 190 7320 200
rect 8600 190 8630 200
rect 8650 190 8670 200
rect 8690 190 8740 200
rect 9140 190 9150 200
rect 9170 190 9180 200
rect 9190 190 9230 200
rect 9290 190 9300 200
rect 9760 190 9790 200
rect 9920 190 9930 200
rect 9950 190 9990 200
rect 0 180 10 190
rect 80 180 120 190
rect 210 180 220 190
rect 320 180 380 190
rect 430 180 470 190
rect 600 180 690 190
rect 840 180 1020 190
rect 4160 180 4540 190
rect 4560 180 4580 190
rect 6090 180 6310 190
rect 6930 180 7330 190
rect 8570 180 8680 190
rect 8690 180 8760 190
rect 8840 180 8860 190
rect 9000 180 9010 190
rect 9070 180 9080 190
rect 9180 180 9210 190
rect 9790 180 9800 190
rect 9830 180 9840 190
rect 9850 180 9860 190
rect 9910 180 9920 190
rect 9950 180 9960 190
rect 9990 180 9990 190
rect 0 170 10 180
rect 100 170 140 180
rect 220 170 230 180
rect 250 170 260 180
rect 310 170 370 180
rect 430 170 490 180
rect 580 170 700 180
rect 830 170 1020 180
rect 4160 170 4540 180
rect 4550 170 4580 180
rect 5000 170 5010 180
rect 6080 170 6310 180
rect 6940 170 7320 180
rect 8580 170 8750 180
rect 8840 170 8860 180
rect 8890 170 8910 180
rect 9030 170 9040 180
rect 9190 170 9200 180
rect 9720 170 9730 180
rect 9850 170 9860 180
rect 0 160 10 170
rect 110 160 140 170
rect 220 160 250 170
rect 280 160 360 170
rect 440 160 510 170
rect 550 160 710 170
rect 810 160 1010 170
rect 4170 160 4540 170
rect 4550 160 4580 170
rect 4820 160 4900 170
rect 6070 160 6080 170
rect 6090 160 6320 170
rect 6960 160 6970 170
rect 6980 160 7320 170
rect 8580 160 8750 170
rect 8830 160 8850 170
rect 8860 160 8900 170
rect 9070 160 9080 170
rect 9710 160 9720 170
rect 9840 160 9850 170
rect 9940 160 9950 170
rect 9970 160 9980 170
rect 110 150 150 160
rect 230 150 250 160
rect 260 150 350 160
rect 450 150 460 160
rect 500 150 720 160
rect 780 150 1010 160
rect 4180 150 4360 160
rect 4380 150 4580 160
rect 4820 150 4920 160
rect 6040 150 6070 160
rect 6100 150 6330 160
rect 6990 150 7330 160
rect 8570 150 8730 160
rect 8830 150 8840 160
rect 8880 150 8890 160
rect 9130 150 9140 160
rect 9150 150 9160 160
rect 9170 150 9180 160
rect 9880 150 9890 160
rect 9940 150 9950 160
rect 9990 150 9990 160
rect 110 140 150 150
rect 230 140 340 150
rect 570 140 1010 150
rect 4190 140 4340 150
rect 4400 140 4570 150
rect 4810 140 4940 150
rect 5010 140 5020 150
rect 6030 140 6050 150
rect 6100 140 6330 150
rect 6990 140 7320 150
rect 8570 140 8730 150
rect 8830 140 8840 150
rect 8900 140 8910 150
rect 9080 140 9090 150
rect 9150 140 9160 150
rect 9190 140 9210 150
rect 9570 140 9580 150
rect 9610 140 9620 150
rect 9940 140 9950 150
rect 110 130 160 140
rect 240 130 330 140
rect 580 130 1010 140
rect 4200 130 4320 140
rect 4430 130 4570 140
rect 4610 130 4630 140
rect 4700 130 4730 140
rect 4800 130 4960 140
rect 6010 130 6040 140
rect 6100 130 6320 140
rect 7000 130 7330 140
rect 8570 130 8740 140
rect 9090 130 9100 140
rect 9140 130 9150 140
rect 9190 130 9220 140
rect 9610 130 9620 140
rect 9710 130 9720 140
rect 9950 130 9970 140
rect 100 120 160 130
rect 250 120 320 130
rect 560 120 1010 130
rect 4210 120 4290 130
rect 4460 120 4570 130
rect 4600 120 4630 130
rect 4690 120 4740 130
rect 4800 120 4900 130
rect 4940 120 4970 130
rect 5990 120 6010 130
rect 6100 120 6320 130
rect 7030 120 7320 130
rect 8570 120 8730 130
rect 9150 120 9160 130
rect 9190 120 9210 130
rect 9370 120 9380 130
rect 9920 120 9930 130
rect 100 110 150 120
rect 250 110 320 120
rect 560 110 1010 120
rect 4220 110 4280 120
rect 4470 110 4570 120
rect 4590 110 4630 120
rect 4680 110 4740 120
rect 4780 110 4880 120
rect 4940 110 4960 120
rect 5840 110 5890 120
rect 5900 110 6020 120
rect 6100 110 6330 120
rect 7030 110 7320 120
rect 8570 110 8730 120
rect 9040 110 9060 120
rect 9150 110 9160 120
rect 9180 110 9210 120
rect 9370 110 9380 120
rect 9400 110 9410 120
rect 9470 110 9490 120
rect 9730 110 9740 120
rect 9850 110 9860 120
rect 100 100 160 110
rect 260 100 320 110
rect 570 100 760 110
rect 780 100 790 110
rect 800 100 1020 110
rect 4240 100 4280 110
rect 4490 100 4560 110
rect 4580 100 4640 110
rect 4660 100 4750 110
rect 4770 100 4850 110
rect 4920 100 4950 110
rect 5830 100 6020 110
rect 6100 100 6330 110
rect 7030 100 7320 110
rect 8570 100 8720 110
rect 8800 100 8830 110
rect 9040 100 9060 110
rect 9150 100 9160 110
rect 9180 100 9220 110
rect 9380 100 9390 110
rect 9480 100 9490 110
rect 9850 100 9860 110
rect 9910 100 9920 110
rect 9940 100 9950 110
rect 9960 100 9980 110
rect 90 90 160 100
rect 260 90 330 100
rect 580 90 730 100
rect 800 90 810 100
rect 840 90 1020 100
rect 4250 90 4280 100
rect 4490 90 4840 100
rect 4920 90 4950 100
rect 5850 90 6020 100
rect 6100 90 6360 100
rect 7040 90 7320 100
rect 8590 90 8720 100
rect 8790 90 8800 100
rect 9140 90 9150 100
rect 9190 90 9240 100
rect 9560 90 9570 100
rect 9890 90 9900 100
rect 9970 90 9980 100
rect 100 80 160 90
rect 260 80 320 90
rect 610 80 630 90
rect 640 80 690 90
rect 860 80 1020 90
rect 4260 80 4280 90
rect 4490 80 4520 90
rect 4530 80 4820 90
rect 4910 80 4940 90
rect 5030 80 5040 90
rect 5890 80 6000 90
rect 6100 80 6360 90
rect 6370 80 6380 90
rect 7050 80 7320 90
rect 8600 80 8710 90
rect 8770 80 8790 90
rect 9060 80 9070 90
rect 9080 80 9090 90
rect 9140 80 9150 90
rect 9180 80 9250 90
rect 9440 80 9450 90
rect 9880 80 9900 90
rect 100 70 160 80
rect 260 70 320 80
rect 860 70 1020 80
rect 4270 70 4310 80
rect 4530 70 4820 80
rect 4890 70 4940 80
rect 5890 70 5970 80
rect 6100 70 6400 80
rect 7060 70 7320 80
rect 8600 70 8710 80
rect 8770 70 8780 80
rect 8930 70 8940 80
rect 8960 70 8970 80
rect 9020 70 9030 80
rect 9070 70 9080 80
rect 9180 70 9230 80
rect 9450 70 9460 80
rect 9560 70 9570 80
rect 9680 70 9700 80
rect 9890 70 9900 80
rect 9910 70 9920 80
rect 9960 70 9970 80
rect 9990 70 9990 80
rect 100 60 150 70
rect 270 60 320 70
rect 860 60 1020 70
rect 4290 60 4320 70
rect 4530 60 4590 70
rect 4610 60 4810 70
rect 4870 60 4940 70
rect 6100 60 6410 70
rect 7070 60 7080 70
rect 7090 60 7320 70
rect 8610 60 8700 70
rect 8900 60 8920 70
rect 8940 60 8960 70
rect 9660 60 9670 70
rect 9700 60 9710 70
rect 9920 60 9930 70
rect 100 50 160 60
rect 270 50 310 60
rect 880 50 1020 60
rect 4310 50 4340 60
rect 4520 50 4570 60
rect 4610 50 4800 60
rect 4850 50 4940 60
rect 6090 50 6420 60
rect 7100 50 7110 60
rect 7120 50 7320 60
rect 8620 50 8690 60
rect 8760 50 8770 60
rect 8950 50 8960 60
rect 9080 50 9090 60
rect 9160 50 9170 60
rect 9280 50 9290 60
rect 9490 50 9500 60
rect 9530 50 9540 60
rect 9550 50 9560 60
rect 9590 50 9610 60
rect 9710 50 9720 60
rect 9900 50 9910 60
rect 9920 50 9930 60
rect 9960 50 9970 60
rect 100 40 170 50
rect 270 40 310 50
rect 880 40 1020 50
rect 4330 40 4340 50
rect 4520 40 4560 50
rect 4600 40 4790 50
rect 4840 40 4940 50
rect 6090 40 6420 50
rect 7130 40 7320 50
rect 8750 40 8760 50
rect 8930 40 8940 50
rect 9080 40 9100 50
rect 9160 40 9170 50
rect 9270 40 9290 50
rect 9510 40 9530 50
rect 9570 40 9590 50
rect 9710 40 9720 50
rect 9750 40 9760 50
rect 100 30 170 40
rect 280 30 310 40
rect 700 30 710 40
rect 890 30 1020 40
rect 4340 30 4360 40
rect 4600 30 4780 40
rect 4830 30 4950 40
rect 6080 30 6430 40
rect 7120 30 7310 40
rect 8740 30 8750 40
rect 9090 30 9100 40
rect 9570 30 9600 40
rect 9690 30 9700 40
rect 9710 30 9720 40
rect 9770 30 9780 40
rect 100 20 160 30
rect 280 20 310 30
rect 690 20 730 30
rect 900 20 1020 30
rect 4350 20 4380 30
rect 4600 20 4940 30
rect 6090 20 6430 30
rect 7120 20 7310 30
rect 8580 20 8590 30
rect 8720 20 8730 30
rect 9090 20 9100 30
rect 9520 20 9530 30
rect 9590 20 9610 30
rect 9680 20 9710 30
rect 9780 20 9790 30
rect 9920 20 9930 30
rect 90 10 170 20
rect 290 10 310 20
rect 680 10 730 20
rect 900 10 1020 20
rect 1290 10 1310 20
rect 4360 10 4380 20
rect 4590 10 4930 20
rect 6090 10 6440 20
rect 7140 10 7300 20
rect 8710 10 8720 20
rect 8910 10 8920 20
rect 9000 10 9040 20
rect 9090 10 9100 20
rect 9170 10 9180 20
rect 9600 10 9630 20
rect 90 0 170 10
rect 290 0 310 10
rect 680 0 730 10
rect 910 0 1010 10
rect 1290 0 1310 10
rect 4370 0 4400 10
rect 4580 0 4660 10
rect 4710 0 4910 10
rect 5930 0 5940 10
rect 6090 0 6440 10
rect 7160 0 7290 10
rect 8580 0 8590 10
rect 8710 0 8720 10
rect 8900 0 8910 10
rect 9090 0 9100 10
rect 9610 0 9640 10
rect 9670 0 9680 10
rect 9710 0 9720 10
rect 9780 0 9790 10
<< metal3 >>
rect 2160 7490 2180 7500
rect 3750 7490 3770 7500
rect 3790 7490 3810 7500
rect 5020 7490 5110 7500
rect 9530 7490 9760 7500
rect 2150 7480 2170 7490
rect 3750 7480 3780 7490
rect 3800 7480 3820 7490
rect 5030 7480 5120 7490
rect 9540 7480 9760 7490
rect 2140 7470 2160 7480
rect 3330 7470 3340 7480
rect 3730 7470 3740 7480
rect 3760 7470 3780 7480
rect 3810 7470 3820 7480
rect 5040 7470 5130 7480
rect 9500 7470 9510 7480
rect 9540 7470 9680 7480
rect 9690 7470 9760 7480
rect 2120 7460 2150 7470
rect 3760 7460 3790 7470
rect 3810 7460 3830 7470
rect 5070 7460 5130 7470
rect 9500 7460 9510 7470
rect 9540 7460 9640 7470
rect 9670 7460 9680 7470
rect 9690 7460 9760 7470
rect 2120 7450 2140 7460
rect 3660 7450 3670 7460
rect 3780 7450 3790 7460
rect 3820 7450 3830 7460
rect 5060 7450 5140 7460
rect 9500 7450 9510 7460
rect 9540 7450 9640 7460
rect 9680 7450 9750 7460
rect 2100 7440 2130 7450
rect 3820 7440 3840 7450
rect 5060 7440 5070 7450
rect 5080 7440 5140 7450
rect 9540 7440 9640 7450
rect 9720 7440 9730 7450
rect 2100 7430 2110 7440
rect 3830 7430 3850 7440
rect 5090 7430 5140 7440
rect 9540 7430 9640 7440
rect 2090 7420 2110 7430
rect 3830 7420 3850 7430
rect 5080 7420 5090 7430
rect 5100 7420 5150 7430
rect 9540 7420 9640 7430
rect 2080 7410 2100 7420
rect 3810 7410 3820 7420
rect 3840 7410 3850 7420
rect 5080 7410 5090 7420
rect 5110 7410 5170 7420
rect 9540 7410 9640 7420
rect 2070 7400 2090 7410
rect 3330 7400 3340 7410
rect 3780 7400 3790 7410
rect 3820 7400 3830 7410
rect 3850 7400 3860 7410
rect 5090 7400 5100 7410
rect 5120 7400 5170 7410
rect 9540 7400 9640 7410
rect 2070 7390 2090 7400
rect 3600 7390 3610 7400
rect 3830 7390 3840 7400
rect 3850 7390 3860 7400
rect 5120 7390 5180 7400
rect 9540 7390 9640 7400
rect 2060 7380 2070 7390
rect 3850 7380 3870 7390
rect 5120 7380 5150 7390
rect 5160 7380 5180 7390
rect 9500 7380 9510 7390
rect 9540 7380 9640 7390
rect 2050 7370 2080 7380
rect 3840 7370 3850 7380
rect 3860 7370 3880 7380
rect 5170 7370 5180 7380
rect 9500 7370 9510 7380
rect 9540 7370 9640 7380
rect 2040 7360 2050 7370
rect 3860 7360 3880 7370
rect 5160 7360 5180 7370
rect 9540 7360 9640 7370
rect 2030 7350 2060 7360
rect 3850 7350 3860 7360
rect 3870 7350 3880 7360
rect 5160 7350 5170 7360
rect 5190 7350 5200 7360
rect 9550 7350 9630 7360
rect 2020 7340 2040 7350
rect 3860 7340 3890 7350
rect 5140 7340 5150 7350
rect 9550 7340 9630 7350
rect 2010 7330 2040 7340
rect 3360 7330 3370 7340
rect 3860 7330 3890 7340
rect 5190 7330 5210 7340
rect 9510 7330 9520 7340
rect 9550 7330 9620 7340
rect 9860 7330 9870 7340
rect 2010 7320 2020 7330
rect 3840 7320 3850 7330
rect 3870 7320 3890 7330
rect 9510 7320 9520 7330
rect 9550 7320 9630 7330
rect 9870 7320 9880 7330
rect 2000 7310 2020 7320
rect 3360 7310 3370 7320
rect 3380 7310 3390 7320
rect 3870 7310 3900 7320
rect 5200 7310 5230 7320
rect 9510 7310 9520 7320
rect 9550 7310 9640 7320
rect 2000 7300 2030 7310
rect 3360 7300 3370 7310
rect 3380 7300 3390 7310
rect 3400 7300 3410 7310
rect 3820 7300 3830 7310
rect 3870 7300 3900 7310
rect 5210 7300 5230 7310
rect 9550 7300 9640 7310
rect 9850 7300 9860 7310
rect 1990 7290 2030 7300
rect 3820 7290 3830 7300
rect 3840 7290 3860 7300
rect 3880 7290 3910 7300
rect 5210 7290 5220 7300
rect 5230 7290 5250 7300
rect 9550 7290 9640 7300
rect 1990 7280 2010 7290
rect 3380 7280 3390 7290
rect 3880 7280 3910 7290
rect 5200 7280 5210 7290
rect 5230 7280 5240 7290
rect 9550 7280 9560 7290
rect 9570 7280 9640 7290
rect 9850 7280 9860 7290
rect 1980 7270 2010 7280
rect 3380 7270 3390 7280
rect 3860 7270 3870 7280
rect 3880 7270 3920 7280
rect 9300 7270 9330 7280
rect 9550 7270 9650 7280
rect 9850 7270 9860 7280
rect 1980 7260 1990 7270
rect 3370 7260 3380 7270
rect 3430 7260 3440 7270
rect 3890 7260 3910 7270
rect 6550 7260 6590 7270
rect 9290 7260 9340 7270
rect 9550 7260 9640 7270
rect 9850 7260 9860 7270
rect 1980 7250 1990 7260
rect 3380 7250 3390 7260
rect 3820 7250 3830 7260
rect 3890 7250 3920 7260
rect 6540 7250 6600 7260
rect 9260 7250 9350 7260
rect 9550 7250 9650 7260
rect 9760 7250 9780 7260
rect 9850 7250 9860 7260
rect 1970 7240 1980 7250
rect 3390 7240 3410 7250
rect 3880 7240 3920 7250
rect 6540 7240 6600 7250
rect 9260 7240 9370 7250
rect 9550 7240 9570 7250
rect 9580 7240 9640 7250
rect 9750 7240 9780 7250
rect 1960 7230 1980 7240
rect 3380 7230 3390 7240
rect 3870 7230 3930 7240
rect 6480 7230 6490 7240
rect 6500 7230 6510 7240
rect 6530 7230 6590 7240
rect 8970 7230 8990 7240
rect 9260 7230 9370 7240
rect 9560 7230 9650 7240
rect 9750 7230 9770 7240
rect 9860 7230 9880 7240
rect 1960 7220 1980 7230
rect 3400 7220 3420 7230
rect 3440 7220 3450 7230
rect 3870 7220 3880 7230
rect 3890 7220 3930 7230
rect 6490 7220 6580 7230
rect 8970 7220 9030 7230
rect 9300 7220 9360 7230
rect 9570 7220 9610 7230
rect 9620 7220 9640 7230
rect 1950 7210 1970 7220
rect 3390 7210 3410 7220
rect 3890 7210 3900 7220
rect 3910 7210 3930 7220
rect 6490 7210 6560 7220
rect 8970 7210 9010 7220
rect 9020 7210 9030 7220
rect 9310 7210 9360 7220
rect 9570 7210 9610 7220
rect 1940 7200 1970 7210
rect 3410 7200 3430 7210
rect 3910 7200 3940 7210
rect 6500 7200 6560 7210
rect 6600 7200 6650 7210
rect 8970 7200 9020 7210
rect 9040 7200 9060 7210
rect 9320 7200 9370 7210
rect 9570 7200 9620 7210
rect 1930 7190 1960 7200
rect 3400 7190 3430 7200
rect 3810 7190 3830 7200
rect 3920 7190 3940 7200
rect 6500 7190 6560 7200
rect 6580 7190 6650 7200
rect 8980 7190 9010 7200
rect 9330 7190 9370 7200
rect 9580 7190 9610 7200
rect 1930 7180 1950 7190
rect 3420 7180 3440 7190
rect 3740 7180 3750 7190
rect 3810 7180 3830 7190
rect 3920 7180 3940 7190
rect 6510 7180 6560 7190
rect 6580 7180 6660 7190
rect 6690 7180 6710 7190
rect 9330 7180 9380 7190
rect 9580 7180 9600 7190
rect 1930 7170 1940 7180
rect 3730 7170 3740 7180
rect 3810 7170 3830 7180
rect 3920 7170 3950 7180
rect 6510 7170 6560 7180
rect 6570 7170 6720 7180
rect 9030 7170 9050 7180
rect 9350 7170 9380 7180
rect 9580 7170 9600 7180
rect 3350 7160 3360 7170
rect 3390 7160 3400 7170
rect 3810 7160 3820 7170
rect 3930 7160 3950 7170
rect 5280 7160 5300 7170
rect 6520 7160 6720 7170
rect 9580 7160 9600 7170
rect 1920 7150 1930 7160
rect 3800 7150 3810 7160
rect 3930 7150 3950 7160
rect 5290 7150 5300 7160
rect 6530 7150 6720 7160
rect 8940 7150 8950 7160
rect 9570 7150 9600 7160
rect 1910 7140 1920 7150
rect 3360 7140 3370 7150
rect 3730 7140 3740 7150
rect 3790 7140 3810 7150
rect 3930 7140 3950 7150
rect 6460 7140 6470 7150
rect 6530 7140 6720 7150
rect 8860 7140 8880 7150
rect 8930 7140 8940 7150
rect 9570 7140 9590 7150
rect 1910 7130 1920 7140
rect 3490 7130 3500 7140
rect 3700 7130 3710 7140
rect 3730 7130 3750 7140
rect 3780 7130 3810 7140
rect 3930 7130 3950 7140
rect 6540 7130 6610 7140
rect 6620 7130 6720 7140
rect 8860 7130 8880 7140
rect 8930 7130 8940 7140
rect 9570 7130 9590 7140
rect 1910 7120 1930 7130
rect 3420 7120 3430 7130
rect 3450 7120 3460 7130
rect 3730 7120 3750 7130
rect 3790 7120 3820 7130
rect 3930 7120 3950 7130
rect 6540 7120 6590 7130
rect 6620 7120 6710 7130
rect 9560 7120 9590 7130
rect 1910 7110 1920 7120
rect 3630 7110 3640 7120
rect 3730 7110 3750 7120
rect 3760 7110 3770 7120
rect 3790 7110 3820 7120
rect 3930 7110 3950 7120
rect 6540 7110 6580 7120
rect 6620 7110 6700 7120
rect 8960 7110 8990 7120
rect 9380 7110 9390 7120
rect 9570 7110 9580 7120
rect 1900 7100 1920 7110
rect 3490 7100 3500 7110
rect 3790 7100 3820 7110
rect 3930 7100 3960 7110
rect 6550 7100 6570 7110
rect 6620 7100 6700 7110
rect 9380 7100 9400 7110
rect 9500 7100 9530 7110
rect 1900 7090 1910 7100
rect 3500 7090 3510 7100
rect 3740 7090 3760 7100
rect 3800 7090 3820 7100
rect 3930 7090 3970 7100
rect 6560 7090 6570 7100
rect 6620 7090 6690 7100
rect 9390 7090 9410 7100
rect 9490 7090 9530 7100
rect 1900 7080 1910 7090
rect 3790 7080 3820 7090
rect 3940 7080 3970 7090
rect 6550 7080 6560 7090
rect 6610 7080 6680 7090
rect 8950 7080 8970 7090
rect 9400 7080 9420 7090
rect 9510 7080 9520 7090
rect 2070 7070 2090 7080
rect 3710 7070 3730 7080
rect 3790 7070 3820 7080
rect 3940 7070 3970 7080
rect 6610 7070 6680 7080
rect 8960 7070 8970 7080
rect 1900 7060 1910 7070
rect 2060 7060 2090 7070
rect 3550 7060 3560 7070
rect 3580 7060 3590 7070
rect 3710 7060 3740 7070
rect 3790 7060 3820 7070
rect 3940 7060 3970 7070
rect 6540 7060 6560 7070
rect 6600 7060 6670 7070
rect 8870 7060 8890 7070
rect 9490 7060 9500 7070
rect 1890 7050 1910 7060
rect 2050 7050 2070 7060
rect 3710 7050 3730 7060
rect 3790 7050 3800 7060
rect 3810 7050 3820 7060
rect 3940 7050 3980 7060
rect 6550 7050 6670 7060
rect 8860 7050 8890 7060
rect 9530 7050 9540 7060
rect 1890 7040 1900 7050
rect 2020 7040 2070 7050
rect 3530 7040 3540 7050
rect 3700 7040 3710 7050
rect 3720 7040 3750 7050
rect 3780 7040 3790 7050
rect 3810 7040 3820 7050
rect 3940 7040 3970 7050
rect 6530 7040 6560 7050
rect 6570 7040 6680 7050
rect 6710 7040 6720 7050
rect 1890 7030 1900 7040
rect 1950 7030 1970 7040
rect 2030 7030 2050 7040
rect 3550 7030 3560 7040
rect 3700 7030 3720 7040
rect 3730 7030 3750 7040
rect 3760 7030 3770 7040
rect 3810 7030 3830 7040
rect 3940 7030 3980 7040
rect 6520 7030 6550 7040
rect 6570 7030 6690 7040
rect 6700 7030 6720 7040
rect 9570 7030 9580 7040
rect 1880 7020 1900 7030
rect 1930 7020 1940 7030
rect 1950 7020 1960 7030
rect 2030 7020 2050 7030
rect 3710 7020 3770 7030
rect 3790 7020 3800 7030
rect 3820 7020 3830 7030
rect 3940 7020 3990 7030
rect 6510 7020 6550 7030
rect 6580 7020 6620 7030
rect 6660 7020 6720 7030
rect 1880 7010 1910 7020
rect 1920 7010 1930 7020
rect 1940 7010 1950 7020
rect 3580 7010 3590 7020
rect 3600 7010 3620 7020
rect 3730 7010 3760 7020
rect 3800 7010 3810 7020
rect 3930 7010 3990 7020
rect 6500 7010 6540 7020
rect 6570 7010 6620 7020
rect 6700 7010 6720 7020
rect 8940 7010 8960 7020
rect 1880 7000 1920 7010
rect 1940 7000 1950 7010
rect 2000 7000 2020 7010
rect 3600 7000 3610 7010
rect 3650 7000 3660 7010
rect 3730 7000 3740 7010
rect 3750 7000 3770 7010
rect 3800 7000 3810 7010
rect 3930 7000 3990 7010
rect 6320 7000 6330 7010
rect 6500 7000 6530 7010
rect 6570 7000 6600 7010
rect 8950 7000 8960 7010
rect 9580 7000 9600 7010
rect 1880 6990 1890 7000
rect 1910 6990 1920 7000
rect 1930 6990 1950 7000
rect 1980 6990 2010 7000
rect 3150 6990 3160 7000
rect 3170 6990 3190 7000
rect 3730 6990 3750 7000
rect 3810 6990 3820 7000
rect 3930 6990 3990 7000
rect 6500 6990 6520 7000
rect 6580 6990 6600 7000
rect 9580 6990 9610 7000
rect 1940 6980 1950 6990
rect 1980 6980 1990 6990
rect 3160 6980 3170 6990
rect 3180 6980 3230 6990
rect 3630 6980 3640 6990
rect 3690 6980 3700 6990
rect 3730 6980 3740 6990
rect 3810 6980 3830 6990
rect 3910 6980 4000 6990
rect 6500 6980 6510 6990
rect 6580 6980 6590 6990
rect 9580 6980 9610 6990
rect 1960 6970 1970 6980
rect 3170 6970 3260 6980
rect 3680 6970 3700 6980
rect 3800 6970 3820 6980
rect 3830 6970 3840 6980
rect 3910 6970 4000 6980
rect 9580 6970 9610 6980
rect 1950 6960 1960 6970
rect 3170 6960 3290 6970
rect 3710 6960 3720 6970
rect 3730 6960 3750 6970
rect 3800 6960 3850 6970
rect 3910 6960 3990 6970
rect 8880 6960 8890 6970
rect 9580 6960 9610 6970
rect 1930 6950 1940 6960
rect 2450 6950 2460 6960
rect 2480 6950 2490 6960
rect 3180 6950 3290 6960
rect 3300 6950 3310 6960
rect 3700 6950 3710 6960
rect 3810 6950 3860 6960
rect 3910 6950 3990 6960
rect 8610 6950 8630 6960
rect 8910 6950 8920 6960
rect 9580 6950 9620 6960
rect 1910 6940 1920 6950
rect 1930 6940 1940 6950
rect 2440 6940 2460 6950
rect 2470 6940 2500 6950
rect 3180 6940 3340 6950
rect 3780 6940 3800 6950
rect 3810 6940 3870 6950
rect 3910 6940 3990 6950
rect 5470 6940 5480 6950
rect 8600 6940 8630 6950
rect 8850 6940 8880 6950
rect 8920 6940 8930 6950
rect 9590 6940 9630 6950
rect 1900 6930 1940 6940
rect 2450 6930 2520 6940
rect 3190 6930 3350 6940
rect 3360 6930 3370 6940
rect 3790 6930 3870 6940
rect 3910 6930 3980 6940
rect 8560 6930 8570 6940
rect 8580 6930 8610 6940
rect 8620 6930 8650 6940
rect 8850 6930 8860 6940
rect 8910 6930 8920 6940
rect 9590 6930 9630 6940
rect 1890 6920 1920 6930
rect 2470 6920 2480 6930
rect 2490 6920 2540 6930
rect 3200 6920 3350 6930
rect 3390 6920 3400 6930
rect 3780 6920 3790 6930
rect 3810 6920 3870 6930
rect 3890 6920 3980 6930
rect 5480 6920 5500 6930
rect 8440 6920 8450 6930
rect 8550 6920 8560 6930
rect 8570 6920 8590 6930
rect 8620 6920 8640 6930
rect 9590 6920 9630 6930
rect 1880 6910 1890 6920
rect 2480 6910 2560 6920
rect 2890 6910 2900 6920
rect 3040 6910 3060 6920
rect 3090 6910 3100 6920
rect 3220 6910 3360 6920
rect 3410 6910 3420 6920
rect 3790 6910 3800 6920
rect 3810 6910 3850 6920
rect 3860 6910 3870 6920
rect 3890 6910 3990 6920
rect 5490 6910 5510 6920
rect 9590 6910 9610 6920
rect 1870 6900 1890 6910
rect 2510 6900 2580 6910
rect 2910 6900 2920 6910
rect 3030 6900 3060 6910
rect 3100 6900 3120 6910
rect 3230 6900 3380 6910
rect 3440 6900 3450 6910
rect 3820 6900 3870 6910
rect 3900 6900 3990 6910
rect 5490 6900 5520 6910
rect 8550 6900 8560 6910
rect 1870 6890 1880 6900
rect 2510 6890 2600 6900
rect 2830 6890 2850 6900
rect 2920 6890 2950 6900
rect 3000 6890 3020 6900
rect 3070 6890 3090 6900
rect 3120 6890 3140 6900
rect 3230 6890 3380 6900
rect 3460 6890 3470 6900
rect 3810 6890 3820 6900
rect 3840 6890 3880 6900
rect 3900 6890 4000 6900
rect 5500 6890 5520 6900
rect 8550 6890 8560 6900
rect 9070 6890 9080 6900
rect 1870 6880 1880 6890
rect 2520 6880 2610 6890
rect 2880 6880 2890 6890
rect 2940 6880 2990 6890
rect 3110 6880 3120 6890
rect 3160 6880 3170 6890
rect 3240 6880 3250 6890
rect 3260 6880 3380 6890
rect 3480 6880 3490 6890
rect 3850 6880 3870 6890
rect 3880 6880 3890 6890
rect 3900 6880 4000 6890
rect 5500 6880 5510 6890
rect 8480 6880 8490 6890
rect 9060 6880 9100 6890
rect 9580 6880 9590 6890
rect 1870 6870 1880 6880
rect 2520 6870 2640 6880
rect 2710 6870 2740 6880
rect 2890 6870 2940 6880
rect 2980 6870 3020 6880
rect 3030 6870 3040 6880
rect 3070 6870 3080 6880
rect 3090 6870 3120 6880
rect 3160 6870 3250 6880
rect 3260 6870 3400 6880
rect 3880 6870 4000 6880
rect 5510 6870 5520 6880
rect 5530 6870 5540 6880
rect 8480 6870 8490 6880
rect 8690 6870 8710 6880
rect 9060 6870 9080 6880
rect 9580 6870 9590 6880
rect 2540 6860 2670 6870
rect 2720 6860 2750 6870
rect 2840 6860 2850 6870
rect 2920 6860 2970 6870
rect 2990 6860 3060 6870
rect 3080 6860 3130 6870
rect 3150 6860 3400 6870
rect 3520 6860 3530 6870
rect 3880 6860 3990 6870
rect 5520 6860 5530 6870
rect 8470 6860 8500 6870
rect 8600 6860 8610 6870
rect 8700 6860 8710 6870
rect 8760 6860 8770 6870
rect 8790 6860 8810 6870
rect 9040 6860 9050 6870
rect 9580 6860 9590 6870
rect 1870 6850 1900 6860
rect 2560 6850 2670 6860
rect 2680 6850 2690 6860
rect 2750 6850 2770 6860
rect 2910 6850 2920 6860
rect 2960 6850 2970 6860
rect 3050 6850 3420 6860
rect 3540 6850 3550 6860
rect 3830 6850 3880 6860
rect 3890 6850 3990 6860
rect 5530 6850 5560 6860
rect 6770 6850 6790 6860
rect 8590 6850 8620 6860
rect 9040 6850 9050 6860
rect 9520 6850 9540 6860
rect 1880 6840 1890 6850
rect 2560 6840 2690 6850
rect 2700 6840 2730 6850
rect 2900 6840 2950 6850
rect 3040 6840 3060 6850
rect 3070 6840 3430 6850
rect 3560 6840 3570 6850
rect 3840 6840 3990 6850
rect 5530 6840 5570 6850
rect 8710 6840 8720 6850
rect 9010 6840 9050 6850
rect 1880 6830 1890 6840
rect 2590 6830 2730 6840
rect 2760 6830 2780 6840
rect 2940 6830 2950 6840
rect 3070 6830 3120 6840
rect 3130 6830 3300 6840
rect 3330 6830 3430 6840
rect 3580 6830 3590 6840
rect 3890 6830 3970 6840
rect 5540 6830 5590 6840
rect 8720 6830 8730 6840
rect 9030 6830 9050 6840
rect 1880 6820 1890 6830
rect 2620 6820 2780 6830
rect 2790 6820 2830 6830
rect 2870 6820 2920 6830
rect 2990 6820 3020 6830
rect 3080 6820 3140 6830
rect 3160 6820 3290 6830
rect 3360 6820 3370 6830
rect 3380 6820 3430 6830
rect 3890 6820 3970 6830
rect 5550 6820 5560 6830
rect 5570 6820 5600 6830
rect 9030 6820 9040 6830
rect 1840 6810 1850 6820
rect 1870 6810 1890 6820
rect 2690 6810 2800 6820
rect 2840 6810 2900 6820
rect 2930 6810 3000 6820
rect 3010 6810 3040 6820
rect 3060 6810 3290 6820
rect 3410 6810 3460 6820
rect 3480 6810 3490 6820
rect 3890 6810 3960 6820
rect 5560 6810 5620 6820
rect 2740 6800 2880 6810
rect 2890 6800 3290 6810
rect 3430 6800 3480 6810
rect 3630 6800 3640 6810
rect 3900 6800 3960 6810
rect 5570 6800 5610 6810
rect 2790 6790 2940 6800
rect 2980 6790 3300 6800
rect 3460 6790 3480 6800
rect 3490 6790 3500 6800
rect 3900 6790 3960 6800
rect 5570 6790 5600 6800
rect 9590 6790 9600 6800
rect 1860 6780 1870 6790
rect 1880 6780 1890 6790
rect 2830 6780 3000 6790
rect 3040 6780 3350 6790
rect 3660 6780 3670 6790
rect 3910 6780 3960 6790
rect 5580 6780 5590 6790
rect 9590 6780 9600 6790
rect 1860 6770 1870 6780
rect 2880 6770 3070 6780
rect 3080 6770 3090 6780
rect 3150 6770 3380 6780
rect 3900 6770 3910 6780
rect 3920 6770 3960 6780
rect 9590 6770 9600 6780
rect 2980 6760 3130 6770
rect 3210 6760 3400 6770
rect 3690 6760 3700 6770
rect 3920 6760 3960 6770
rect 5630 6760 5650 6770
rect 9570 6760 9580 6770
rect 1870 6750 1880 6760
rect 1960 6750 1970 6760
rect 2400 6750 2420 6760
rect 3060 6750 3190 6760
rect 3300 6750 3370 6760
rect 3380 6750 3410 6760
rect 3920 6750 3960 6760
rect 5630 6750 5650 6760
rect 9550 6750 9560 6760
rect 1860 6740 1870 6750
rect 1970 6740 1980 6750
rect 2360 6740 2440 6750
rect 3140 6740 3250 6750
rect 3350 6740 3360 6750
rect 3380 6740 3400 6750
rect 3410 6740 3420 6750
rect 3720 6740 3730 6750
rect 3930 6740 3960 6750
rect 5620 6740 5640 6750
rect 5650 6740 5660 6750
rect 9590 6740 9600 6750
rect 1850 6730 1860 6740
rect 2340 6730 2460 6740
rect 3230 6730 3310 6740
rect 3420 6730 3450 6740
rect 3930 6730 3970 6740
rect 9540 6730 9550 6740
rect 9590 6730 9600 6740
rect 1850 6720 1870 6730
rect 2310 6720 2480 6730
rect 3260 6720 3350 6730
rect 3460 6720 3480 6730
rect 3940 6720 3970 6730
rect 8980 6720 8990 6730
rect 9590 6720 9600 6730
rect 1830 6710 1840 6720
rect 1870 6710 1880 6720
rect 2300 6710 2390 6720
rect 2430 6710 2500 6720
rect 3310 6710 3320 6720
rect 3330 6710 3390 6720
rect 3480 6710 3510 6720
rect 3760 6710 3770 6720
rect 3940 6710 3970 6720
rect 9530 6710 9540 6720
rect 9590 6710 9600 6720
rect 1840 6700 1850 6710
rect 2290 6700 2330 6710
rect 2340 6700 2350 6710
rect 2450 6700 2500 6710
rect 3360 6700 3430 6710
rect 3770 6700 3780 6710
rect 3940 6700 3970 6710
rect 9570 6700 9580 6710
rect 9590 6700 9600 6710
rect 1810 6690 1840 6700
rect 1850 6690 1860 6700
rect 2270 6690 2310 6700
rect 2480 6690 2510 6700
rect 2540 6690 2560 6700
rect 3420 6690 3470 6700
rect 3810 6690 3820 6700
rect 3940 6690 3970 6700
rect 9570 6690 9580 6700
rect 1790 6680 1800 6690
rect 1830 6680 1840 6690
rect 2260 6680 2280 6690
rect 2480 6680 2520 6690
rect 3440 6680 3490 6690
rect 3930 6680 3970 6690
rect 9570 6680 9580 6690
rect 1770 6670 1780 6680
rect 1800 6670 1810 6680
rect 1820 6670 1840 6680
rect 1850 6670 1900 6680
rect 2250 6670 2270 6680
rect 2480 6670 2550 6680
rect 3470 6670 3540 6680
rect 3950 6670 3980 6680
rect 8930 6670 8940 6680
rect 9550 6670 9580 6680
rect 9950 6670 9960 6680
rect 1750 6660 1760 6670
rect 1860 6660 1870 6670
rect 2250 6660 2270 6670
rect 2480 6660 2550 6670
rect 3490 6660 3550 6670
rect 3820 6660 3830 6670
rect 3950 6660 3980 6670
rect 8930 6660 8940 6670
rect 9550 6660 9570 6670
rect 9600 6660 9610 6670
rect 9910 6660 9920 6670
rect 2240 6650 2270 6660
rect 2490 6650 2560 6660
rect 3550 6650 3570 6660
rect 3960 6650 3980 6660
rect 8570 6650 8580 6660
rect 9540 6650 9570 6660
rect 9600 6650 9610 6660
rect 1710 6640 1730 6650
rect 1800 6640 1840 6650
rect 2230 6640 2260 6650
rect 2510 6640 2560 6650
rect 3570 6640 3600 6650
rect 3960 6640 3990 6650
rect 9540 6640 9560 6650
rect 9850 6640 9860 6650
rect 1750 6630 1760 6640
rect 2220 6630 2250 6640
rect 2520 6630 2570 6640
rect 3610 6630 3620 6640
rect 3970 6630 3990 6640
rect 9480 6630 9490 6640
rect 9540 6630 9550 6640
rect 9820 6630 9830 6640
rect 1660 6620 1740 6630
rect 2220 6620 2250 6630
rect 2540 6620 2570 6630
rect 3630 6620 3650 6630
rect 3970 6620 3990 6630
rect 8510 6620 8520 6630
rect 9520 6620 9540 6630
rect 9790 6620 9800 6630
rect 1610 6610 1620 6620
rect 1720 6610 1740 6620
rect 1750 6610 1760 6620
rect 2220 6610 2240 6620
rect 2540 6610 2580 6620
rect 3650 6610 3680 6620
rect 3970 6610 3990 6620
rect 8500 6610 8510 6620
rect 9520 6610 9560 6620
rect 9760 6610 9770 6620
rect 1590 6600 1600 6610
rect 1750 6600 1760 6610
rect 2210 6600 2240 6610
rect 2540 6600 2580 6610
rect 3680 6600 3690 6610
rect 3970 6600 3990 6610
rect 6040 6600 6050 6610
rect 6070 6600 6090 6610
rect 8760 6600 8780 6610
rect 9520 6600 9580 6610
rect 1580 6590 1590 6600
rect 1640 6590 1670 6600
rect 1740 6590 1760 6600
rect 2200 6590 2240 6600
rect 2550 6590 2590 6600
rect 3690 6590 3730 6600
rect 3980 6590 3990 6600
rect 6070 6590 6080 6600
rect 6220 6590 6260 6600
rect 6270 6590 6300 6600
rect 8760 6590 8770 6600
rect 9520 6590 9590 6600
rect 9680 6590 9690 6600
rect 1340 6580 1350 6590
rect 1470 6580 1480 6590
rect 1550 6580 1570 6590
rect 1620 6580 1630 6590
rect 1640 6580 1650 6590
rect 1750 6580 1770 6590
rect 2190 6580 2230 6590
rect 2540 6580 2590 6590
rect 3730 6580 3740 6590
rect 3990 6580 4000 6590
rect 5940 6580 5950 6590
rect 6060 6580 6080 6590
rect 6090 6580 6110 6590
rect 6120 6580 6130 6590
rect 6210 6580 6260 6590
rect 6270 6580 6320 6590
rect 6340 6580 6350 6590
rect 8540 6580 8570 6590
rect 8690 6580 8700 6590
rect 8870 6580 8890 6590
rect 9480 6580 9490 6590
rect 9560 6580 9610 6590
rect 9670 6580 9680 6590
rect 1350 6570 1360 6580
rect 1530 6570 1550 6580
rect 1610 6570 1640 6580
rect 1760 6570 1780 6580
rect 2080 6570 2090 6580
rect 2110 6570 2120 6580
rect 2190 6570 2210 6580
rect 2540 6570 2600 6580
rect 3740 6570 3760 6580
rect 4000 6570 4010 6580
rect 5940 6570 5960 6580
rect 6010 6570 6020 6580
rect 6050 6570 6130 6580
rect 6210 6570 6270 6580
rect 6280 6570 6360 6580
rect 6380 6570 6390 6580
rect 8550 6570 8560 6580
rect 8600 6570 8610 6580
rect 8750 6570 8760 6580
rect 8870 6570 8880 6580
rect 9520 6570 9530 6580
rect 9570 6570 9630 6580
rect 9640 6570 9680 6580
rect 1350 6560 1360 6570
rect 1370 6560 1380 6570
rect 1490 6560 1540 6570
rect 1610 6560 1630 6570
rect 1760 6560 1790 6570
rect 2080 6560 2090 6570
rect 2150 6560 2160 6570
rect 2550 6560 2600 6570
rect 3760 6560 3770 6570
rect 4000 6560 4010 6570
rect 5940 6560 5970 6570
rect 6000 6560 6010 6570
rect 6020 6560 6040 6570
rect 6050 6560 6070 6570
rect 6090 6560 6140 6570
rect 6170 6560 6220 6570
rect 6230 6560 6260 6570
rect 6270 6560 6410 6570
rect 6430 6560 6460 6570
rect 6560 6560 6580 6570
rect 8750 6560 8760 6570
rect 9490 6560 9500 6570
rect 9580 6560 9590 6570
rect 9640 6560 9680 6570
rect 1350 6550 1360 6560
rect 1380 6550 1390 6560
rect 1480 6550 1520 6560
rect 1610 6550 1620 6560
rect 1630 6550 1750 6560
rect 1770 6550 1780 6560
rect 2010 6550 2030 6560
rect 2040 6550 2060 6560
rect 2560 6550 2590 6560
rect 3780 6550 3790 6560
rect 4000 6550 4010 6560
rect 5950 6550 5980 6560
rect 6000 6550 6010 6560
rect 6030 6550 6080 6560
rect 6090 6550 6130 6560
rect 6140 6550 6220 6560
rect 6240 6550 6470 6560
rect 6510 6550 6600 6560
rect 9490 6550 9500 6560
rect 9510 6550 9520 6560
rect 1350 6540 1360 6550
rect 1390 6540 1400 6550
rect 1450 6540 1460 6550
rect 1490 6540 1500 6550
rect 1750 6540 1760 6550
rect 1770 6540 1800 6550
rect 2050 6540 2060 6550
rect 2570 6540 2600 6550
rect 3790 6540 3800 6550
rect 4000 6540 4020 6550
rect 5950 6540 5970 6550
rect 5980 6540 5990 6550
rect 6010 6540 6030 6550
rect 6040 6540 6060 6550
rect 6070 6540 6080 6550
rect 6100 6540 6220 6550
rect 6240 6540 6250 6550
rect 6270 6540 6360 6550
rect 6380 6540 6420 6550
rect 6450 6540 6470 6550
rect 6480 6540 6540 6550
rect 6560 6540 6610 6550
rect 8020 6540 8040 6550
rect 8730 6540 8750 6550
rect 9500 6540 9510 6550
rect 1370 6530 1440 6540
rect 1770 6530 1800 6540
rect 2050 6530 2090 6540
rect 2570 6530 2580 6540
rect 3820 6530 3830 6540
rect 5810 6530 5820 6540
rect 5960 6530 6010 6540
rect 6020 6530 6030 6540
rect 6050 6530 6090 6540
rect 6110 6530 6220 6540
rect 6240 6530 6250 6540
rect 6270 6530 6350 6540
rect 6460 6530 6480 6540
rect 6490 6530 6510 6540
rect 6570 6530 6600 6540
rect 6620 6530 6670 6540
rect 8720 6530 8740 6540
rect 9550 6530 9560 6540
rect 1330 6520 1420 6530
rect 1780 6520 1800 6530
rect 2050 6520 2060 6530
rect 2070 6520 2090 6530
rect 2220 6520 2260 6530
rect 2560 6520 2570 6530
rect 3840 6520 3850 6530
rect 3950 6520 3960 6530
rect 4010 6520 4020 6530
rect 5810 6520 5830 6530
rect 5840 6520 5880 6530
rect 5970 6520 6000 6530
rect 6020 6520 6040 6530
rect 6050 6520 6060 6530
rect 6080 6520 6090 6530
rect 6120 6520 6230 6530
rect 6240 6520 6260 6530
rect 6280 6520 6310 6530
rect 6340 6520 6360 6530
rect 6450 6520 6460 6530
rect 6560 6520 6620 6530
rect 6630 6520 6670 6530
rect 8710 6520 8740 6530
rect 9970 6520 9980 6530
rect 1300 6510 1320 6520
rect 2070 6510 2090 6520
rect 2230 6510 2280 6520
rect 2530 6510 2540 6520
rect 3850 6510 3870 6520
rect 4010 6510 4020 6520
rect 5820 6510 5840 6520
rect 5850 6510 5890 6520
rect 5970 6510 6010 6520
rect 6030 6510 6050 6520
rect 6080 6510 6090 6520
rect 6100 6510 6170 6520
rect 6210 6510 6270 6520
rect 6280 6510 6310 6520
rect 6560 6510 6580 6520
rect 6630 6510 6660 6520
rect 8710 6510 8730 6520
rect 9190 6510 9200 6520
rect 9410 6510 9420 6520
rect 9940 6510 9950 6520
rect 1270 6500 1290 6510
rect 2240 6500 2250 6510
rect 2270 6500 2280 6510
rect 2410 6500 2420 6510
rect 2490 6500 2500 6510
rect 3870 6500 3890 6510
rect 4010 6500 4030 6510
rect 5800 6500 5840 6510
rect 5870 6500 5890 6510
rect 5940 6500 5960 6510
rect 5980 6500 6000 6510
rect 6010 6500 6020 6510
rect 6030 6500 6060 6510
rect 6090 6500 6110 6510
rect 6240 6500 6270 6510
rect 6310 6500 6330 6510
rect 6600 6500 6610 6510
rect 6620 6500 6660 6510
rect 8020 6500 8050 6510
rect 8700 6500 8720 6510
rect 9410 6500 9420 6510
rect 1270 6490 1300 6500
rect 2250 6490 2260 6500
rect 2270 6490 2280 6500
rect 3880 6490 3900 6500
rect 5800 6490 5810 6500
rect 5820 6490 5860 6500
rect 5930 6490 6070 6500
rect 6240 6490 6250 6500
rect 6320 6490 6340 6500
rect 6610 6490 6690 6500
rect 8020 6490 8050 6500
rect 8690 6490 8720 6500
rect 1260 6480 1270 6490
rect 1810 6480 1820 6490
rect 2130 6480 2140 6490
rect 3900 6480 3920 6490
rect 4020 6480 4030 6490
rect 5740 6480 5750 6490
rect 5760 6480 5770 6490
rect 5790 6480 5800 6490
rect 5810 6480 5880 6490
rect 5930 6480 5990 6490
rect 6000 6480 6080 6490
rect 6340 6480 6360 6490
rect 6620 6480 6720 6490
rect 8030 6480 8050 6490
rect 8690 6480 8710 6490
rect 9680 6480 9690 6490
rect 9850 6480 9860 6490
rect 1320 6470 1340 6480
rect 1810 6470 1830 6480
rect 2150 6470 2160 6480
rect 2270 6470 2290 6480
rect 3920 6470 3930 6480
rect 4020 6470 4030 6480
rect 5770 6470 5910 6480
rect 5950 6470 5960 6480
rect 6010 6470 6090 6480
rect 6350 6470 6360 6480
rect 6610 6470 6730 6480
rect 8030 6470 8040 6480
rect 8680 6470 8700 6480
rect 9800 6470 9810 6480
rect 1230 6460 1240 6470
rect 1360 6460 1370 6470
rect 1690 6460 1720 6470
rect 1820 6460 1830 6470
rect 2150 6460 2170 6470
rect 2200 6460 2210 6470
rect 2270 6460 2290 6470
rect 2560 6460 2570 6470
rect 3930 6460 3950 6470
rect 4030 6460 4040 6470
rect 5780 6460 5820 6470
rect 5840 6460 5910 6470
rect 6020 6460 6100 6470
rect 6590 6460 6730 6470
rect 8680 6460 8700 6470
rect 9760 6460 9770 6470
rect 1670 6450 1730 6460
rect 1820 6450 1830 6460
rect 2150 6450 2170 6460
rect 2220 6450 2290 6460
rect 2300 6450 2310 6460
rect 3950 6450 3960 6460
rect 4010 6450 4020 6460
rect 5720 6450 5730 6460
rect 5870 6450 5910 6460
rect 5950 6450 6000 6460
rect 6030 6450 6100 6460
rect 6600 6450 6750 6460
rect 8670 6450 8690 6460
rect 9680 6450 9740 6460
rect 1300 6440 1340 6450
rect 1660 6440 1740 6450
rect 1820 6440 1830 6450
rect 2150 6440 2160 6450
rect 2250 6440 2260 6450
rect 2290 6440 2320 6450
rect 2380 6440 2390 6450
rect 4030 6440 4040 6450
rect 5680 6440 5700 6450
rect 5720 6440 5790 6450
rect 5810 6440 5840 6450
rect 5870 6440 6000 6450
rect 6030 6440 6090 6450
rect 6610 6440 6660 6450
rect 6670 6440 6780 6450
rect 8670 6440 8680 6450
rect 1220 6430 1240 6440
rect 1290 6430 1300 6440
rect 1320 6430 1330 6440
rect 1650 6430 1670 6440
rect 1690 6430 1740 6440
rect 1820 6430 1830 6440
rect 1870 6430 1890 6440
rect 1920 6430 1930 6440
rect 2130 6430 2150 6440
rect 2280 6430 2290 6440
rect 2330 6430 2340 6440
rect 2370 6430 2380 6440
rect 3980 6430 3990 6440
rect 5680 6430 5810 6440
rect 5970 6430 6080 6440
rect 6630 6430 6670 6440
rect 6680 6430 6790 6440
rect 8660 6430 8680 6440
rect 9580 6430 9600 6440
rect 1220 6420 1250 6430
rect 1290 6420 1300 6430
rect 1320 6420 1330 6430
rect 1650 6420 1670 6430
rect 1690 6420 1740 6430
rect 1820 6420 1830 6430
rect 1870 6420 1940 6430
rect 2110 6420 2140 6430
rect 2310 6420 2320 6430
rect 5690 6420 5810 6430
rect 5960 6420 6100 6430
rect 6640 6420 6690 6430
rect 6700 6420 6800 6430
rect 8650 6420 8670 6430
rect 9580 6420 9600 6430
rect 9640 6420 9650 6430
rect 1220 6410 1230 6420
rect 1280 6410 1330 6420
rect 1450 6410 1460 6420
rect 1640 6410 1670 6420
rect 1690 6410 1750 6420
rect 1800 6410 1840 6420
rect 1850 6410 1940 6420
rect 2060 6410 2120 6420
rect 2350 6410 2370 6420
rect 4010 6410 4020 6420
rect 5690 6410 5820 6420
rect 5880 6410 5900 6420
rect 5980 6410 6100 6420
rect 6660 6410 6690 6420
rect 6720 6410 6810 6420
rect 8660 6410 8670 6420
rect 9590 6410 9600 6420
rect 9630 6410 9640 6420
rect 1200 6400 1210 6410
rect 1220 6400 1230 6410
rect 1240 6400 1250 6410
rect 1270 6400 1320 6410
rect 1430 6400 1460 6410
rect 1640 6400 1650 6410
rect 1820 6400 1940 6410
rect 2060 6400 2080 6410
rect 2090 6400 2110 6410
rect 5720 6400 5760 6410
rect 5770 6400 5780 6410
rect 5800 6400 5840 6410
rect 5990 6400 6000 6410
rect 6010 6400 6050 6410
rect 6090 6400 6110 6410
rect 6670 6400 6690 6410
rect 6720 6400 6770 6410
rect 6780 6400 6830 6410
rect 8640 6400 8660 6410
rect 9630 6400 9640 6410
rect 1200 6390 1220 6400
rect 1230 6390 1250 6400
rect 1260 6390 1300 6400
rect 1330 6390 1370 6400
rect 1400 6390 1450 6400
rect 1630 6390 1640 6400
rect 1780 6390 1810 6400
rect 1830 6390 1970 6400
rect 2050 6390 2080 6400
rect 2090 6390 2100 6400
rect 4040 6390 4050 6400
rect 5670 6390 5700 6400
rect 5870 6390 6070 6400
rect 6090 6390 6110 6400
rect 6780 6390 6830 6400
rect 8640 6390 8660 6400
rect 9630 6390 9640 6400
rect 1230 6380 1240 6390
rect 1260 6380 1340 6390
rect 1400 6380 1410 6390
rect 1430 6380 1460 6390
rect 1630 6380 1640 6390
rect 1680 6380 1700 6390
rect 1730 6380 1760 6390
rect 1820 6380 1900 6390
rect 1930 6380 1970 6390
rect 2010 6380 2090 6390
rect 2390 6380 2400 6390
rect 5660 6380 5720 6390
rect 5840 6380 5890 6390
rect 5930 6380 5960 6390
rect 6010 6380 6120 6390
rect 6280 6380 6310 6390
rect 6800 6380 6830 6390
rect 8630 6380 8650 6390
rect 1210 6370 1240 6380
rect 1340 6370 1360 6380
rect 1430 6370 1440 6380
rect 1620 6370 1630 6380
rect 1670 6370 1730 6380
rect 1840 6370 1890 6380
rect 1950 6370 2060 6380
rect 5650 6370 5670 6380
rect 5700 6370 5800 6380
rect 5930 6370 5960 6380
rect 5990 6370 6140 6380
rect 6260 6370 6350 6380
rect 6800 6370 6820 6380
rect 7500 6370 7510 6380
rect 8630 6370 8650 6380
rect 9610 6370 9630 6380
rect 1220 6360 1230 6370
rect 1390 6360 1400 6370
rect 1610 6360 1620 6370
rect 1670 6360 1710 6370
rect 1840 6360 1880 6370
rect 1970 6360 2020 6370
rect 4080 6360 4090 6370
rect 5660 6360 5790 6370
rect 5910 6360 6290 6370
rect 6300 6360 6350 6370
rect 6810 6360 6830 6370
rect 8620 6360 8640 6370
rect 9480 6360 9490 6370
rect 9610 6360 9630 6370
rect 1260 6350 1270 6360
rect 1400 6350 1410 6360
rect 1610 6350 1620 6360
rect 1660 6350 1680 6360
rect 1840 6350 1880 6360
rect 1970 6350 2020 6360
rect 4090 6350 4100 6360
rect 5660 6350 5750 6360
rect 5880 6350 5980 6360
rect 6030 6350 6270 6360
rect 6340 6350 6360 6360
rect 6830 6350 6840 6360
rect 8050 6350 8060 6360
rect 8620 6350 8630 6360
rect 9450 6350 9460 6360
rect 9470 6350 9490 6360
rect 1240 6340 1250 6350
rect 1270 6340 1280 6350
rect 1370 6340 1380 6350
rect 1400 6340 1410 6350
rect 1600 6340 1610 6350
rect 1640 6340 1670 6350
rect 1840 6340 1850 6350
rect 1970 6340 2020 6350
rect 2400 6340 2410 6350
rect 5570 6340 5730 6350
rect 5820 6340 5900 6350
rect 6050 6340 6080 6350
rect 6350 6340 6380 6350
rect 6810 6340 6840 6350
rect 8050 6340 8070 6350
rect 8610 6340 8630 6350
rect 9420 6340 9430 6350
rect 9450 6340 9460 6350
rect 1210 6330 1220 6340
rect 1260 6330 1290 6340
rect 1390 6330 1410 6340
rect 1600 6330 1610 6340
rect 1630 6330 1660 6340
rect 1840 6330 1870 6340
rect 1900 6330 1910 6340
rect 1970 6330 2020 6340
rect 2380 6330 2420 6340
rect 5480 6330 5560 6340
rect 5670 6330 5690 6340
rect 5700 6330 5710 6340
rect 5820 6330 5860 6340
rect 6360 6330 6400 6340
rect 6810 6330 6850 6340
rect 7590 6330 7600 6340
rect 8050 6330 8060 6340
rect 8610 6330 8620 6340
rect 9380 6330 9400 6340
rect 9410 6330 9420 6340
rect 9630 6330 9640 6340
rect 1270 6320 1280 6330
rect 1290 6320 1300 6330
rect 1390 6320 1410 6330
rect 1590 6320 1650 6330
rect 1840 6320 1900 6330
rect 1970 6320 2020 6330
rect 2390 6320 2400 6330
rect 2410 6320 2420 6330
rect 2450 6320 2460 6330
rect 5430 6320 5480 6330
rect 5650 6320 5690 6330
rect 5820 6320 5850 6330
rect 6370 6320 6430 6330
rect 6800 6320 6860 6330
rect 7590 6320 7610 6330
rect 8600 6320 8620 6330
rect 9350 6320 9380 6330
rect 9410 6320 9420 6330
rect 9460 6320 9470 6330
rect 9500 6320 9510 6330
rect 1200 6310 1240 6320
rect 1270 6310 1290 6320
rect 1300 6310 1310 6320
rect 1390 6310 1410 6320
rect 1590 6310 1630 6320
rect 1840 6310 1890 6320
rect 2010 6310 2020 6320
rect 2390 6310 2400 6320
rect 2450 6310 2460 6320
rect 5400 6310 5440 6320
rect 5480 6310 5500 6320
rect 5630 6310 5660 6320
rect 5820 6310 5840 6320
rect 6400 6310 6440 6320
rect 6800 6310 6860 6320
rect 7590 6310 7610 6320
rect 8600 6310 8610 6320
rect 9320 6310 9330 6320
rect 9340 6310 9380 6320
rect 9390 6310 9400 6320
rect 9410 6310 9420 6320
rect 9460 6310 9470 6320
rect 9590 6310 9600 6320
rect 1200 6300 1240 6310
rect 1250 6300 1260 6310
rect 1280 6300 1300 6310
rect 1310 6300 1320 6310
rect 1390 6300 1410 6310
rect 1590 6300 1620 6310
rect 1840 6300 1880 6310
rect 2410 6300 2420 6310
rect 2450 6300 2470 6310
rect 4150 6300 4160 6310
rect 5380 6300 5390 6310
rect 5620 6300 5640 6310
rect 5810 6300 5840 6310
rect 6420 6300 6460 6310
rect 6770 6300 6870 6310
rect 7590 6300 7610 6310
rect 8590 6300 8610 6310
rect 9290 6300 9300 6310
rect 9330 6300 9370 6310
rect 9500 6300 9510 6310
rect 9590 6300 9600 6310
rect 9630 6300 9640 6310
rect 1210 6290 1230 6300
rect 1250 6290 1270 6300
rect 1390 6290 1400 6300
rect 1590 6290 1620 6300
rect 1830 6290 1860 6300
rect 2400 6290 2420 6300
rect 4160 6290 4170 6300
rect 5360 6290 5370 6300
rect 5710 6290 5820 6300
rect 6450 6290 6490 6300
rect 6780 6290 6840 6300
rect 8580 6290 8590 6300
rect 9280 6290 9350 6300
rect 9420 6290 9430 6300
rect 9470 6290 9480 6300
rect 9610 6290 9620 6300
rect 9630 6290 9640 6300
rect 9970 6290 9990 6300
rect 1210 6280 1230 6290
rect 1270 6280 1310 6290
rect 1320 6280 1330 6290
rect 1390 6280 1410 6290
rect 1590 6280 1610 6290
rect 1830 6280 1860 6290
rect 2400 6280 2420 6290
rect 4170 6280 4180 6290
rect 5360 6280 5380 6290
rect 5680 6280 5710 6290
rect 6460 6280 6520 6290
rect 6780 6280 6800 6290
rect 6820 6280 6840 6290
rect 7390 6280 7400 6290
rect 8580 6280 8590 6290
rect 9300 6280 9330 6290
rect 9470 6280 9480 6290
rect 9500 6280 9510 6290
rect 9960 6280 9990 6290
rect 1200 6270 1240 6280
rect 1280 6270 1290 6280
rect 1400 6270 1410 6280
rect 1590 6270 1600 6280
rect 1830 6270 1850 6280
rect 2400 6270 2420 6280
rect 4180 6270 4190 6280
rect 5630 6270 5690 6280
rect 6460 6270 6530 6280
rect 6830 6270 6840 6280
rect 8070 6270 8080 6280
rect 8580 6270 8590 6280
rect 9270 6270 9280 6280
rect 9320 6270 9330 6280
rect 9470 6270 9480 6280
rect 9500 6270 9520 6280
rect 9880 6270 9890 6280
rect 9970 6270 9980 6280
rect 1200 6260 1240 6270
rect 1290 6260 1300 6270
rect 1330 6260 1340 6270
rect 1400 6260 1410 6270
rect 1820 6260 1830 6270
rect 2390 6260 2400 6270
rect 2410 6260 2420 6270
rect 4190 6260 4200 6270
rect 5620 6260 5680 6270
rect 6470 6260 6540 6270
rect 6790 6260 6810 6270
rect 6840 6260 6850 6270
rect 7430 6260 7450 6270
rect 8070 6260 8080 6270
rect 8580 6260 8590 6270
rect 9320 6260 9340 6270
rect 9400 6260 9410 6270
rect 9500 6260 9530 6270
rect 9560 6260 9570 6270
rect 9610 6260 9620 6270
rect 9870 6260 9880 6270
rect 9900 6260 9910 6270
rect 9950 6260 9960 6270
rect 9980 6260 9990 6270
rect 1200 6250 1250 6260
rect 1260 6250 1320 6260
rect 1360 6250 1370 6260
rect 1390 6250 1410 6260
rect 1810 6250 1820 6260
rect 2400 6250 2420 6260
rect 4200 6250 4210 6260
rect 5320 6250 5330 6260
rect 5610 6250 5650 6260
rect 6480 6250 6540 6260
rect 6800 6250 6810 6260
rect 6850 6250 6860 6260
rect 7430 6250 7440 6260
rect 8070 6250 8080 6260
rect 8570 6250 8590 6260
rect 9310 6250 9320 6260
rect 9400 6250 9410 6260
rect 9420 6250 9440 6260
rect 9480 6250 9540 6260
rect 9830 6250 9860 6260
rect 9870 6250 9880 6260
rect 9900 6250 9920 6260
rect 9930 6250 9950 6260
rect 1180 6240 1230 6250
rect 1260 6240 1380 6250
rect 1400 6240 1410 6250
rect 2400 6240 2420 6250
rect 2450 6240 2460 6250
rect 4210 6240 4220 6250
rect 5370 6240 5380 6250
rect 5590 6240 5630 6250
rect 6510 6240 6560 6250
rect 6840 6240 6870 6250
rect 7620 6240 7630 6250
rect 8070 6240 8090 6250
rect 9250 6240 9260 6250
rect 9300 6240 9310 6250
rect 9490 6240 9510 6250
rect 9640 6240 9650 6250
rect 9810 6240 9820 6250
rect 9870 6240 9890 6250
rect 9940 6240 9950 6250
rect 1180 6230 1330 6240
rect 1350 6230 1380 6240
rect 1390 6230 1410 6240
rect 1800 6230 1810 6240
rect 2400 6230 2420 6240
rect 2450 6230 2460 6240
rect 4220 6230 4230 6240
rect 5300 6230 5310 6240
rect 5350 6230 5370 6240
rect 5580 6230 5620 6240
rect 6520 6230 6570 6240
rect 6850 6230 6880 6240
rect 7450 6230 7470 6240
rect 8070 6230 8080 6240
rect 9260 6230 9300 6240
rect 9370 6230 9380 6240
rect 9440 6230 9450 6240
rect 9470 6230 9480 6240
rect 9610 6230 9630 6240
rect 9640 6230 9650 6240
rect 9810 6230 9820 6240
rect 9940 6230 9980 6240
rect 1180 6220 1300 6230
rect 1320 6220 1330 6230
rect 1360 6220 1370 6230
rect 1390 6220 1420 6230
rect 2400 6220 2420 6230
rect 5300 6220 5310 6230
rect 5340 6220 5360 6230
rect 5550 6220 5600 6230
rect 6540 6220 6570 6230
rect 6780 6220 6800 6230
rect 6850 6220 6890 6230
rect 8070 6220 8080 6230
rect 9240 6220 9250 6230
rect 9290 6220 9300 6230
rect 9360 6220 9380 6230
rect 9640 6220 9650 6230
rect 9920 6220 9940 6230
rect 9980 6220 9990 6230
rect 1170 6210 1280 6220
rect 1290 6210 1300 6220
rect 1320 6210 1330 6220
rect 1400 6210 1420 6220
rect 1790 6210 1800 6220
rect 2400 6210 2420 6220
rect 5320 6210 5340 6220
rect 5540 6210 5590 6220
rect 6550 6210 6590 6220
rect 6780 6210 6820 6220
rect 6860 6210 6900 6220
rect 8070 6210 8090 6220
rect 9290 6210 9320 6220
rect 9350 6210 9380 6220
rect 9640 6210 9650 6220
rect 9900 6210 9910 6220
rect 9920 6210 9940 6220
rect 9950 6210 9960 6220
rect 9990 6210 9990 6220
rect 1180 6200 1280 6210
rect 1300 6200 1340 6210
rect 1370 6200 1380 6210
rect 1400 6200 1420 6210
rect 1780 6200 1790 6210
rect 2400 6200 2420 6210
rect 4240 6200 4250 6210
rect 5280 6200 5290 6210
rect 5310 6200 5320 6210
rect 5520 6200 5570 6210
rect 6550 6200 6610 6210
rect 6780 6200 6840 6210
rect 6870 6200 6910 6210
rect 7630 6200 7650 6210
rect 8070 6200 8100 6210
rect 9230 6200 9240 6210
rect 9280 6200 9290 6210
rect 9300 6200 9310 6210
rect 9320 6200 9330 6210
rect 9350 6200 9360 6210
rect 9370 6200 9380 6210
rect 9910 6200 9930 6210
rect 9940 6200 9950 6210
rect 1170 6190 1290 6200
rect 1310 6190 1320 6200
rect 1330 6190 1340 6200
rect 1370 6190 1380 6200
rect 1400 6190 1420 6200
rect 1780 6190 1790 6200
rect 2400 6190 2420 6200
rect 5270 6190 5280 6200
rect 5290 6190 5300 6200
rect 5510 6190 5550 6200
rect 6560 6190 6630 6200
rect 6800 6190 6830 6200
rect 6880 6190 6920 6200
rect 7630 6190 7650 6200
rect 9300 6190 9310 6200
rect 9670 6190 9680 6200
rect 1170 6180 1260 6190
rect 1280 6180 1290 6190
rect 1310 6180 1320 6190
rect 1330 6180 1340 6190
rect 1370 6180 1380 6190
rect 1400 6180 1420 6190
rect 1780 6180 1790 6190
rect 2370 6180 2390 6190
rect 2400 6180 2420 6190
rect 5260 6180 5290 6190
rect 5490 6180 5540 6190
rect 6570 6180 6650 6190
rect 6810 6180 6820 6190
rect 6890 6180 6940 6190
rect 9210 6180 9220 6190
rect 9230 6180 9240 6190
rect 9250 6180 9280 6190
rect 9290 6180 9300 6190
rect 9940 6180 9950 6190
rect 9990 6180 9990 6190
rect 1170 6170 1220 6180
rect 1240 6170 1260 6180
rect 1280 6170 1300 6180
rect 1340 6170 1350 6180
rect 1400 6170 1420 6180
rect 1600 6170 1620 6180
rect 1780 6170 1790 6180
rect 2370 6170 2420 6180
rect 5250 6170 5280 6180
rect 5470 6170 5510 6180
rect 6610 6170 6650 6180
rect 6900 6170 6960 6180
rect 7480 6170 7500 6180
rect 7660 6170 7670 6180
rect 9210 6170 9220 6180
rect 9240 6170 9260 6180
rect 9280 6170 9290 6180
rect 9930 6170 9950 6180
rect 1170 6160 1180 6170
rect 1210 6160 1230 6170
rect 1240 6160 1260 6170
rect 1290 6160 1300 6170
rect 1330 6160 1350 6170
rect 1380 6160 1420 6170
rect 1610 6160 1630 6170
rect 1750 6160 1770 6170
rect 1780 6160 1790 6170
rect 2380 6160 2420 6170
rect 4270 6160 4280 6170
rect 5260 6160 5270 6170
rect 5280 6160 5300 6170
rect 5460 6160 5490 6170
rect 6620 6160 6660 6170
rect 6900 6160 6960 6170
rect 7480 6160 7490 6170
rect 7590 6160 7610 6170
rect 7660 6160 7670 6170
rect 9210 6160 9230 6170
rect 9240 6160 9260 6170
rect 9640 6160 9650 6170
rect 9940 6160 9950 6170
rect 1150 6150 1160 6160
rect 1170 6150 1180 6160
rect 1210 6150 1230 6160
rect 1240 6150 1270 6160
rect 1340 6150 1350 6160
rect 1390 6150 1430 6160
rect 1630 6150 1640 6160
rect 1740 6150 1780 6160
rect 2380 6150 2420 6160
rect 4280 6150 4290 6160
rect 5250 6150 5260 6160
rect 5290 6150 5300 6160
rect 5440 6150 5470 6160
rect 5480 6150 5490 6160
rect 6630 6150 6660 6160
rect 6900 6150 6970 6160
rect 7620 6150 7630 6160
rect 7980 6150 7990 6160
rect 8110 6150 8120 6160
rect 9220 6150 9230 6160
rect 9940 6150 9960 6160
rect 9990 6150 9990 6160
rect 1130 6140 1170 6150
rect 1210 6140 1270 6150
rect 1310 6140 1320 6150
rect 1330 6140 1360 6150
rect 1390 6140 1400 6150
rect 1420 6140 1430 6150
rect 1650 6140 1680 6150
rect 1740 6140 1790 6150
rect 2410 6140 2420 6150
rect 5240 6140 5250 6150
rect 5280 6140 5290 6150
rect 5430 6140 5470 6150
rect 6640 6140 6670 6150
rect 6900 6140 6980 6150
rect 7630 6140 7650 6150
rect 7910 6140 7930 6150
rect 8080 6140 8120 6150
rect 8510 6140 8520 6150
rect 9200 6140 9210 6150
rect 9940 6140 9960 6150
rect 1140 6130 1160 6140
rect 1220 6130 1230 6140
rect 1240 6130 1280 6140
rect 1310 6130 1360 6140
rect 1400 6130 1410 6140
rect 1420 6130 1430 6140
rect 1650 6130 1690 6140
rect 1720 6130 1770 6140
rect 1790 6130 1800 6140
rect 2420 6130 2430 6140
rect 5220 6130 5240 6140
rect 5260 6130 5270 6140
rect 5430 6130 5470 6140
rect 6630 6130 6680 6140
rect 6900 6130 6980 6140
rect 7540 6130 7580 6140
rect 8510 6130 8520 6140
rect 8550 6130 8570 6140
rect 9180 6130 9190 6140
rect 9920 6130 9930 6140
rect 9960 6130 9970 6140
rect 1110 6120 1120 6130
rect 1130 6120 1150 6130
rect 1180 6120 1190 6130
rect 1210 6120 1230 6130
rect 1240 6120 1270 6130
rect 1350 6120 1360 6130
rect 1420 6120 1430 6130
rect 1650 6120 1680 6130
rect 1730 6120 1770 6130
rect 1790 6120 1800 6130
rect 2420 6120 2430 6130
rect 5220 6120 5240 6130
rect 5250 6120 5260 6130
rect 5270 6120 5280 6130
rect 5420 6120 5450 6130
rect 5460 6120 5470 6130
rect 6660 6120 6690 6130
rect 6900 6120 6910 6130
rect 6920 6120 6990 6130
rect 7550 6120 7580 6130
rect 7690 6120 7700 6130
rect 8510 6120 8520 6130
rect 9150 6120 9160 6130
rect 9900 6120 9910 6130
rect 9920 6120 9930 6130
rect 9950 6120 9970 6130
rect 1170 6110 1180 6120
rect 1210 6110 1240 6120
rect 1250 6110 1280 6120
rect 1660 6110 1680 6120
rect 1730 6110 1760 6120
rect 1790 6110 1810 6120
rect 5210 6110 5230 6120
rect 5250 6110 5270 6120
rect 5410 6110 5450 6120
rect 6660 6110 6690 6120
rect 6920 6110 6990 6120
rect 7520 6110 7540 6120
rect 7550 6110 7560 6120
rect 7680 6110 7690 6120
rect 8510 6110 8540 6120
rect 9120 6110 9130 6120
rect 9850 6110 9860 6120
rect 9880 6110 9900 6120
rect 9950 6110 9980 6120
rect 1120 6100 1180 6110
rect 1190 6100 1200 6110
rect 1220 6100 1240 6110
rect 1250 6100 1290 6110
rect 1670 6100 1680 6110
rect 1730 6100 1750 6110
rect 1790 6100 1810 6110
rect 2430 6100 2440 6110
rect 5200 6100 5230 6110
rect 5260 6100 5270 6110
rect 5400 6100 5430 6110
rect 6670 6100 6700 6110
rect 6930 6100 6990 6110
rect 7520 6100 7550 6110
rect 7680 6100 7700 6110
rect 8510 6100 8540 6110
rect 9090 6100 9100 6110
rect 9420 6100 9450 6110
rect 9850 6100 9900 6110
rect 9950 6100 9980 6110
rect 1120 6090 1170 6100
rect 1180 6090 1210 6100
rect 1230 6090 1260 6100
rect 1270 6090 1300 6100
rect 1680 6090 1690 6100
rect 1740 6090 1750 6100
rect 1790 6090 1810 6100
rect 2470 6090 2480 6100
rect 5220 6090 5230 6100
rect 5240 6090 5250 6100
rect 5390 6090 5430 6100
rect 6670 6090 6710 6100
rect 6950 6090 6990 6100
rect 7540 6090 7550 6100
rect 9070 6090 9080 6100
rect 9380 6090 9390 6100
rect 9870 6090 9940 6100
rect 9950 6090 9980 6100
rect 1110 6080 1210 6090
rect 1230 6080 1300 6090
rect 1680 6080 1700 6090
rect 1740 6080 1750 6090
rect 1800 6080 1820 6090
rect 5210 6080 5230 6090
rect 5250 6080 5260 6090
rect 5390 6080 5410 6090
rect 6680 6080 6710 6090
rect 6950 6080 6990 6090
rect 7610 6080 7620 6090
rect 9030 6080 9060 6090
rect 9350 6080 9360 6090
rect 9880 6080 9890 6090
rect 9910 6080 9930 6090
rect 9960 6080 9970 6090
rect 1110 6070 1120 6080
rect 1140 6070 1220 6080
rect 1230 6070 1300 6080
rect 1690 6070 1760 6080
rect 1800 6070 1820 6080
rect 2440 6070 2450 6080
rect 5200 6070 5210 6080
rect 5230 6070 5250 6080
rect 5380 6070 5410 6080
rect 6680 6070 6720 6080
rect 6970 6070 7000 6080
rect 7530 6070 7540 6080
rect 9000 6070 9010 6080
rect 9020 6070 9030 6080
rect 9340 6070 9350 6080
rect 9480 6070 9490 6080
rect 9890 6070 9900 6080
rect 9950 6070 9960 6080
rect 810 6060 820 6070
rect 1010 6060 1040 6070
rect 1060 6060 1100 6070
rect 1150 6060 1300 6070
rect 1700 6060 1780 6070
rect 1800 6060 1820 6070
rect 3840 6060 3850 6070
rect 5190 6060 5200 6070
rect 5230 6060 5240 6070
rect 5380 6060 5400 6070
rect 6690 6060 6720 6070
rect 6960 6060 7000 6070
rect 8960 6060 8980 6070
rect 9010 6060 9020 6070
rect 9440 6060 9450 6070
rect 9860 6060 9870 6070
rect 9900 6060 9950 6070
rect 800 6050 840 6060
rect 850 6050 860 6060
rect 1060 6050 1290 6060
rect 1730 6050 1740 6060
rect 1790 6050 1820 6060
rect 2450 6050 2460 6060
rect 3780 6050 3790 6060
rect 4330 6050 4340 6060
rect 5180 6050 5190 6060
rect 5200 6050 5210 6060
rect 5220 6050 5240 6060
rect 5380 6050 5400 6060
rect 6700 6050 6730 6060
rect 6960 6050 6990 6060
rect 7590 6050 7600 6060
rect 8930 6050 8940 6060
rect 9250 6050 9260 6060
rect 9340 6050 9350 6060
rect 9930 6050 9940 6060
rect 780 6040 830 6050
rect 840 6040 860 6050
rect 910 6040 940 6050
rect 1040 6040 1070 6050
rect 1100 6040 1110 6050
rect 1130 6040 1200 6050
rect 1230 6040 1250 6050
rect 1260 6040 1270 6050
rect 1730 6040 1740 6050
rect 3800 6040 3810 6050
rect 5180 6040 5200 6050
rect 5210 6040 5230 6050
rect 5380 6040 5400 6050
rect 6700 6040 6730 6050
rect 6960 6040 7000 6050
rect 7510 6040 7530 6050
rect 7590 6040 7600 6050
rect 8910 6040 8930 6050
rect 9220 6040 9230 6050
rect 9440 6040 9450 6050
rect 9930 6040 9940 6050
rect 770 6030 830 6040
rect 840 6030 860 6040
rect 880 6030 1020 6040
rect 1030 6030 1060 6040
rect 1080 6030 1100 6040
rect 1120 6030 1160 6040
rect 1230 6030 1250 6040
rect 1730 6030 1750 6040
rect 4000 6030 4010 6040
rect 5200 6030 5220 6040
rect 5380 6030 5390 6040
rect 6710 6030 6740 6040
rect 6970 6030 7000 6040
rect 7500 6030 7510 6040
rect 7580 6030 7590 6040
rect 7630 6030 7640 6040
rect 8850 6030 8860 6040
rect 9920 6030 9940 6040
rect 770 6020 810 6030
rect 820 6020 840 6030
rect 890 6020 900 6030
rect 940 6020 1020 6030
rect 1060 6020 1100 6030
rect 1110 6020 1130 6030
rect 1240 6020 1260 6030
rect 1720 6020 1750 6030
rect 2470 6020 2480 6030
rect 4010 6020 4020 6030
rect 5190 6020 5200 6030
rect 5370 6020 5390 6030
rect 6720 6020 6740 6030
rect 6980 6020 7010 6030
rect 8420 6020 8440 6030
rect 8820 6020 8830 6030
rect 9910 6020 9940 6030
rect 760 6010 790 6020
rect 810 6010 830 6020
rect 940 6010 1060 6020
rect 1090 6010 1100 6020
rect 1110 6010 1130 6020
rect 1190 6010 1200 6020
rect 1720 6010 1750 6020
rect 5180 6010 5190 6020
rect 5370 6010 5390 6020
rect 6720 6010 6740 6020
rect 6980 6010 7010 6020
rect 7400 6010 7420 6020
rect 7490 6010 7500 6020
rect 8430 6010 8440 6020
rect 8790 6010 8800 6020
rect 9110 6010 9130 6020
rect 9350 6010 9360 6020
rect 9870 6010 9880 6020
rect 9900 6010 9940 6020
rect 750 6000 760 6010
rect 770 6000 780 6010
rect 790 6000 830 6010
rect 950 6000 1030 6010
rect 1070 6000 1090 6010
rect 1110 6000 1120 6010
rect 1160 6000 1170 6010
rect 1190 6000 1200 6010
rect 1720 6000 1770 6010
rect 3940 6000 3950 6010
rect 3960 6000 3970 6010
rect 4010 6000 4020 6010
rect 5370 6000 5390 6010
rect 6720 6000 6750 6010
rect 6980 6000 7010 6010
rect 7400 6000 7420 6010
rect 7490 6000 7510 6010
rect 7600 6000 7610 6010
rect 8420 6000 8430 6010
rect 8760 6000 8770 6010
rect 9100 6000 9110 6010
rect 9450 6000 9460 6010
rect 9880 6000 9900 6010
rect 9920 6000 9930 6010
rect 750 5990 760 6000
rect 770 5990 780 6000
rect 790 5990 830 6000
rect 950 5990 970 6000
rect 990 5990 1010 6000
rect 1050 5990 1090 6000
rect 1110 5990 1120 6000
rect 1190 5990 1200 6000
rect 1720 5990 1810 6000
rect 2490 5990 2500 6000
rect 3800 5990 3810 6000
rect 4010 5990 4020 6000
rect 5160 5990 5180 6000
rect 5370 5990 5380 6000
rect 6720 5990 6750 6000
rect 6980 5990 7010 6000
rect 7390 5990 7410 6000
rect 7470 5990 7510 6000
rect 7590 5990 7610 6000
rect 8730 5990 8760 6000
rect 9050 5990 9060 6000
rect 9140 5990 9150 6000
rect 9180 5990 9190 6000
rect 9450 5990 9460 6000
rect 9900 5990 9920 6000
rect 9930 5990 9940 6000
rect 740 5980 750 5990
rect 770 5980 780 5990
rect 790 5980 840 5990
rect 970 5980 990 5990
rect 1100 5980 1130 5990
rect 1180 5980 1190 5990
rect 1710 5980 1810 5990
rect 2500 5980 2510 5990
rect 3820 5980 3830 5990
rect 4010 5980 4020 5990
rect 5150 5980 5170 5990
rect 5370 5980 5380 5990
rect 6730 5980 6760 5990
rect 6990 5980 7010 5990
rect 7400 5980 7410 5990
rect 7470 5980 7490 5990
rect 7530 5980 7550 5990
rect 7590 5980 7600 5990
rect 7690 5980 7720 5990
rect 8330 5980 8350 5990
rect 8400 5980 8420 5990
rect 8700 5980 8720 5990
rect 8730 5980 8740 5990
rect 9030 5980 9040 5990
rect 9900 5980 9910 5990
rect 9960 5980 9970 5990
rect 740 5970 750 5980
rect 780 5970 840 5980
rect 870 5970 880 5980
rect 980 5970 1000 5980
rect 1090 5970 1120 5980
rect 1720 5970 1820 5980
rect 3850 5970 3860 5980
rect 3920 5970 3930 5980
rect 5150 5970 5160 5980
rect 5360 5970 5370 5980
rect 6730 5970 6760 5980
rect 6990 5970 7010 5980
rect 7450 5970 7470 5980
rect 7500 5970 7520 5980
rect 7530 5970 7550 5980
rect 7580 5970 7590 5980
rect 7660 5970 7690 5980
rect 7720 5970 7730 5980
rect 8330 5970 8350 5980
rect 8660 5970 8670 5980
rect 9230 5970 9240 5980
rect 9260 5970 9270 5980
rect 9300 5970 9310 5980
rect 9360 5970 9370 5980
rect 9420 5970 9430 5980
rect 770 5960 840 5970
rect 1050 5960 1080 5970
rect 1100 5960 1110 5970
rect 1720 5960 1780 5970
rect 1790 5960 1800 5970
rect 1810 5960 1820 5970
rect 1990 5960 2010 5970
rect 2490 5960 2510 5970
rect 3930 5960 3950 5970
rect 4500 5960 4530 5970
rect 5150 5960 5180 5970
rect 5350 5960 5370 5970
rect 6730 5960 6770 5970
rect 6990 5960 7000 5970
rect 7280 5960 7300 5970
rect 7430 5960 7460 5970
rect 7510 5960 7520 5970
rect 7530 5960 7550 5970
rect 7650 5960 7660 5970
rect 7670 5960 7680 5970
rect 7700 5960 7730 5970
rect 8330 5960 8350 5970
rect 8360 5960 8370 5970
rect 8390 5960 8410 5970
rect 8620 5960 8640 5970
rect 9100 5960 9110 5970
rect 9190 5960 9200 5970
rect 9430 5960 9440 5970
rect 9950 5960 9960 5970
rect 9980 5960 9990 5970
rect 730 5950 740 5960
rect 760 5950 840 5960
rect 910 5950 920 5960
rect 1170 5950 1180 5960
rect 1710 5950 1720 5960
rect 1730 5950 1820 5960
rect 1990 5950 2000 5960
rect 2480 5950 2530 5960
rect 3190 5950 3200 5960
rect 3860 5950 3870 5960
rect 5160 5950 5170 5960
rect 5350 5950 5360 5960
rect 6730 5950 6780 5960
rect 7530 5950 7550 5960
rect 7670 5950 7680 5960
rect 7700 5950 7710 5960
rect 8310 5950 8350 5960
rect 8360 5950 8370 5960
rect 8390 5950 8400 5960
rect 8590 5950 8610 5960
rect 8960 5950 8970 5960
rect 9090 5950 9110 5960
rect 9410 5950 9420 5960
rect 9500 5950 9510 5960
rect 9950 5950 9980 5960
rect 720 5940 730 5950
rect 760 5940 800 5950
rect 840 5940 860 5950
rect 960 5940 980 5950
rect 1170 5940 1180 5950
rect 1700 5940 1810 5950
rect 2480 5940 2540 5950
rect 3180 5940 3210 5950
rect 4340 5940 4350 5950
rect 5150 5940 5160 5950
rect 5350 5940 5360 5950
rect 6730 5940 6790 5950
rect 7000 5940 7010 5950
rect 7320 5940 7330 5950
rect 7490 5940 7550 5950
rect 8390 5940 8400 5950
rect 8560 5940 8580 5950
rect 8960 5940 8970 5950
rect 9010 5940 9020 5950
rect 9100 5940 9110 5950
rect 9280 5940 9290 5950
rect 9370 5940 9380 5950
rect 9900 5940 9910 5950
rect 700 5930 720 5940
rect 760 5930 780 5940
rect 790 5930 800 5940
rect 840 5930 850 5940
rect 1700 5930 1790 5940
rect 2470 5930 2520 5940
rect 2540 5930 2550 5940
rect 3170 5930 3210 5940
rect 3940 5930 3950 5940
rect 5350 5930 5360 5940
rect 6740 5930 6790 5940
rect 7000 5930 7010 5940
rect 7310 5930 7350 5940
rect 8120 5930 8130 5940
rect 8370 5930 8390 5940
rect 8850 5930 8860 5940
rect 9370 5930 9380 5940
rect 9960 5930 9970 5940
rect 700 5920 710 5930
rect 750 5920 760 5930
rect 790 5920 810 5930
rect 1720 5920 1780 5930
rect 2460 5920 2540 5930
rect 2550 5920 2570 5930
rect 3160 5920 3210 5930
rect 3840 5920 3860 5930
rect 5340 5920 5360 5930
rect 6740 5920 6800 5930
rect 7000 5920 7010 5930
rect 7310 5920 7320 5930
rect 7340 5920 7360 5930
rect 8090 5920 8100 5930
rect 8370 5920 8380 5930
rect 8510 5920 8520 5930
rect 8830 5920 8840 5930
rect 8920 5920 8930 5930
rect 8970 5920 8980 5930
rect 9020 5920 9030 5930
rect 9150 5920 9160 5930
rect 9200 5920 9210 5930
rect 9960 5920 9970 5930
rect 680 5910 700 5920
rect 750 5910 760 5920
rect 770 5910 830 5920
rect 1740 5910 1760 5920
rect 2390 5910 2410 5920
rect 2450 5910 2560 5920
rect 3150 5910 3220 5920
rect 3760 5910 3770 5920
rect 3840 5910 3860 5920
rect 5340 5910 5360 5920
rect 6750 5910 6800 5920
rect 7000 5910 7010 5920
rect 8370 5910 8380 5920
rect 8470 5910 8480 5920
rect 8930 5910 8940 5920
rect 9020 5910 9030 5920
rect 9150 5910 9160 5920
rect 9200 5910 9210 5920
rect 670 5900 700 5910
rect 740 5900 750 5910
rect 770 5900 810 5910
rect 820 5900 830 5910
rect 920 5900 950 5910
rect 1740 5900 1760 5910
rect 1830 5900 1860 5910
rect 2360 5900 2560 5910
rect 3150 5900 3220 5910
rect 3760 5900 3770 5910
rect 3860 5900 3870 5910
rect 3920 5900 3930 5910
rect 4010 5900 4020 5910
rect 4210 5900 4220 5910
rect 5120 5900 5130 5910
rect 5340 5900 5350 5910
rect 6760 5900 6800 5910
rect 7000 5900 7010 5910
rect 7300 5900 7320 5910
rect 8250 5900 8260 5910
rect 8350 5900 8360 5910
rect 8440 5900 8450 5910
rect 9070 5900 9080 5910
rect 9320 5900 9330 5910
rect 9380 5900 9390 5910
rect 650 5890 690 5900
rect 740 5890 790 5900
rect 820 5890 830 5900
rect 920 5890 950 5900
rect 1010 5890 1020 5900
rect 1740 5890 1860 5900
rect 2350 5890 2570 5900
rect 3140 5890 3220 5900
rect 3770 5890 3780 5900
rect 4010 5890 4020 5900
rect 4230 5890 4240 5900
rect 4280 5890 4290 5900
rect 5340 5890 5350 5900
rect 6760 5890 6800 5900
rect 7000 5890 7020 5900
rect 7290 5890 7330 5900
rect 7360 5890 7390 5900
rect 8150 5890 8160 5900
rect 8350 5890 8360 5900
rect 8410 5890 8420 5900
rect 8720 5890 8730 5900
rect 8800 5890 8810 5900
rect 8940 5890 8950 5900
rect 8980 5890 8990 5900
rect 9280 5890 9290 5900
rect 640 5880 710 5890
rect 800 5880 820 5890
rect 930 5880 940 5890
rect 1770 5880 1780 5890
rect 1790 5880 1830 5890
rect 1850 5880 1870 5890
rect 2340 5880 2590 5890
rect 3110 5880 3230 5890
rect 3750 5880 3760 5890
rect 3880 5880 3890 5890
rect 4010 5880 4030 5890
rect 5340 5880 5350 5890
rect 6760 5880 6800 5890
rect 7010 5880 7020 5890
rect 7300 5880 7330 5890
rect 7350 5880 7370 5890
rect 7380 5880 7390 5890
rect 8030 5880 8040 5890
rect 8150 5880 8160 5890
rect 8370 5880 8390 5890
rect 8690 5880 8700 5890
rect 8900 5880 8910 5890
rect 9080 5880 9090 5890
rect 9210 5880 9220 5890
rect 390 5870 400 5880
rect 640 5870 690 5880
rect 790 5870 800 5880
rect 870 5870 880 5880
rect 940 5870 980 5880
rect 1850 5870 1870 5880
rect 2330 5870 2600 5880
rect 3100 5870 3230 5880
rect 3890 5870 3900 5880
rect 4020 5870 4030 5880
rect 5110 5870 5120 5880
rect 5330 5870 5350 5880
rect 6760 5870 6800 5880
rect 6990 5870 7000 5880
rect 7010 5870 7020 5880
rect 7330 5870 7340 5880
rect 7350 5870 7360 5880
rect 7380 5870 7390 5880
rect 7930 5870 7950 5880
rect 8030 5870 8040 5880
rect 8150 5870 8160 5880
rect 8340 5870 8350 5880
rect 8660 5870 8670 5880
rect 8750 5870 8760 5880
rect 8900 5870 8910 5880
rect 9090 5870 9100 5880
rect 9210 5870 9220 5880
rect 370 5860 380 5870
rect 590 5860 600 5870
rect 650 5860 670 5870
rect 770 5860 870 5870
rect 890 5860 900 5870
rect 960 5860 1000 5870
rect 1850 5860 1870 5870
rect 2300 5860 2590 5870
rect 3080 5860 3240 5870
rect 3770 5860 3780 5870
rect 3820 5860 3860 5870
rect 3880 5860 3890 5870
rect 5110 5860 5120 5870
rect 5330 5860 5350 5870
rect 6770 5860 6780 5870
rect 6990 5860 7020 5870
rect 7370 5860 7400 5870
rect 7960 5860 7980 5870
rect 7990 5860 8010 5870
rect 8150 5860 8160 5870
rect 8310 5860 8320 5870
rect 8730 5860 8740 5870
rect 8990 5860 9000 5870
rect 9160 5860 9170 5870
rect 9210 5860 9220 5870
rect 9300 5860 9310 5870
rect 9920 5860 9930 5870
rect 340 5850 380 5860
rect 590 5850 610 5860
rect 630 5850 650 5860
rect 770 5850 790 5860
rect 880 5850 890 5860
rect 960 5850 970 5860
rect 1850 5850 1870 5860
rect 2290 5850 2600 5860
rect 3060 5850 3230 5860
rect 3760 5850 3770 5860
rect 3800 5850 3810 5860
rect 3820 5850 3840 5860
rect 3860 5850 3880 5860
rect 5330 5850 5350 5860
rect 6770 5850 6780 5860
rect 6990 5850 7020 5860
rect 7880 5850 7890 5860
rect 7960 5850 7970 5860
rect 8000 5850 8010 5860
rect 8150 5850 8160 5860
rect 8260 5850 8280 5860
rect 8710 5850 8720 5860
rect 8910 5850 8920 5860
rect 8950 5850 8960 5860
rect 9100 5850 9110 5860
rect 9160 5850 9170 5860
rect 9220 5850 9230 5860
rect 9920 5850 9930 5860
rect 580 5840 630 5850
rect 770 5840 780 5850
rect 890 5840 930 5850
rect 1860 5840 1880 5850
rect 2280 5840 2310 5850
rect 2360 5840 2610 5850
rect 3050 5840 3230 5850
rect 3860 5840 3870 5850
rect 5100 5840 5110 5850
rect 5330 5840 5350 5850
rect 6770 5840 6790 5850
rect 7000 5840 7020 5850
rect 7870 5840 7880 5850
rect 7960 5840 7970 5850
rect 8090 5840 8100 5850
rect 8140 5840 8160 5850
rect 8240 5840 8250 5850
rect 8710 5840 8720 5850
rect 8910 5840 8920 5850
rect 9000 5840 9010 5850
rect 9970 5840 9990 5850
rect 580 5830 600 5840
rect 760 5830 780 5840
rect 1850 5830 1880 5840
rect 2270 5830 2300 5840
rect 2360 5830 2460 5840
rect 2490 5830 2620 5840
rect 3030 5830 3230 5840
rect 3740 5830 3770 5840
rect 3790 5830 3800 5840
rect 3830 5830 3860 5840
rect 3940 5830 3950 5840
rect 4590 5830 4610 5840
rect 5100 5830 5110 5840
rect 5330 5830 5350 5840
rect 6780 5830 6800 5840
rect 6990 5830 7000 5840
rect 7010 5830 7020 5840
rect 7880 5830 7890 5840
rect 7970 5830 7980 5840
rect 8090 5830 8100 5840
rect 8110 5830 8130 5840
rect 8220 5830 8230 5840
rect 8630 5830 8640 5840
rect 8670 5830 8680 5840
rect 8800 5830 8810 5840
rect 9000 5830 9010 5840
rect 9160 5830 9170 5840
rect 9920 5830 9930 5840
rect 9960 5830 9990 5840
rect 570 5820 590 5830
rect 750 5820 790 5830
rect 1850 5820 1880 5830
rect 2270 5820 2300 5830
rect 2360 5820 2430 5830
rect 2490 5820 2620 5830
rect 3020 5820 3150 5830
rect 3170 5820 3230 5830
rect 3740 5820 3750 5830
rect 3940 5820 3950 5830
rect 3960 5820 3970 5830
rect 4570 5820 4610 5830
rect 5330 5820 5350 5830
rect 6780 5820 6800 5830
rect 6990 5820 7000 5830
rect 7980 5820 8000 5830
rect 8100 5820 8110 5830
rect 9120 5820 9130 5830
rect 9960 5820 9970 5830
rect 560 5810 580 5820
rect 630 5810 650 5820
rect 740 5810 750 5820
rect 1850 5810 1890 5820
rect 2250 5810 2290 5820
rect 2350 5810 2420 5820
rect 2490 5810 2620 5820
rect 3000 5810 3130 5820
rect 3170 5810 3230 5820
rect 3750 5810 3760 5820
rect 3800 5810 3830 5820
rect 3860 5810 3870 5820
rect 3940 5810 3950 5820
rect 4570 5810 4620 5820
rect 5330 5810 5350 5820
rect 6790 5810 6800 5820
rect 7860 5810 7870 5820
rect 7880 5810 7890 5820
rect 8160 5810 8170 5820
rect 8920 5810 8930 5820
rect 9010 5810 9020 5820
rect 9060 5810 9070 5820
rect 9950 5810 9960 5820
rect 550 5800 570 5810
rect 610 5800 630 5810
rect 800 5800 810 5810
rect 840 5800 850 5810
rect 1850 5800 1890 5810
rect 2250 5800 2270 5810
rect 2350 5800 2420 5810
rect 2490 5800 2610 5810
rect 3000 5800 3110 5810
rect 3160 5800 3230 5810
rect 3750 5800 3770 5810
rect 3780 5800 3790 5810
rect 3810 5800 3820 5810
rect 3840 5800 3850 5810
rect 3900 5800 3910 5810
rect 3950 5800 3960 5810
rect 4580 5800 4620 5810
rect 5090 5800 5100 5810
rect 5330 5800 5350 5810
rect 6790 5800 6800 5810
rect 7000 5800 7010 5810
rect 7830 5800 7850 5810
rect 7870 5800 7890 5810
rect 8010 5800 8020 5810
rect 8120 5800 8140 5810
rect 8680 5800 8690 5810
rect 8720 5800 8730 5810
rect 550 5790 560 5800
rect 610 5790 650 5800
rect 720 5790 740 5800
rect 1870 5790 1890 5800
rect 1900 5790 1930 5800
rect 2240 5790 2260 5800
rect 2350 5790 2410 5800
rect 2480 5790 2610 5800
rect 2970 5790 3080 5800
rect 3160 5790 3240 5800
rect 3840 5790 3860 5800
rect 3890 5790 3920 5800
rect 4050 5790 4060 5800
rect 4580 5790 4620 5800
rect 5090 5790 5100 5800
rect 5330 5790 5340 5800
rect 6790 5790 6810 5800
rect 7000 5790 7010 5800
rect 7750 5790 7790 5800
rect 7870 5790 7900 5800
rect 7910 5790 7920 5800
rect 7990 5790 8000 5800
rect 8100 5790 8110 5800
rect 8810 5790 8820 5800
rect 8910 5790 8920 5800
rect 610 5780 650 5790
rect 700 5780 720 5790
rect 880 5780 910 5790
rect 1870 5780 1950 5790
rect 2230 5780 2250 5790
rect 2340 5780 2390 5790
rect 2470 5780 2480 5790
rect 2490 5780 2600 5790
rect 2960 5780 3110 5790
rect 3170 5780 3240 5790
rect 3840 5780 3860 5790
rect 3880 5780 3890 5790
rect 3900 5780 3920 5790
rect 3970 5780 3980 5790
rect 4060 5780 4070 5790
rect 4480 5780 4490 5790
rect 4560 5780 4620 5790
rect 5330 5780 5340 5790
rect 6800 5780 6810 5790
rect 6990 5780 7010 5790
rect 7780 5780 7790 5790
rect 8050 5780 8070 5790
rect 8900 5780 8910 5790
rect 8950 5780 8960 5790
rect 550 5770 570 5780
rect 600 5770 610 5780
rect 630 5770 650 5780
rect 690 5770 720 5780
rect 820 5770 830 5780
rect 840 5770 870 5780
rect 1880 5770 1950 5780
rect 2220 5770 2230 5780
rect 2330 5770 2350 5780
rect 2370 5770 2400 5780
rect 2470 5770 2600 5780
rect 2960 5770 3120 5780
rect 3180 5770 3240 5780
rect 3870 5770 3880 5780
rect 3960 5770 3970 5780
rect 4070 5770 4080 5780
rect 4560 5770 4610 5780
rect 4680 5770 4720 5780
rect 4740 5770 4750 5780
rect 5320 5770 5340 5780
rect 6800 5770 6810 5780
rect 6990 5770 7010 5780
rect 7750 5770 7770 5780
rect 8010 5770 8030 5780
rect 8380 5770 8390 5780
rect 540 5760 580 5770
rect 640 5760 660 5770
rect 680 5760 710 5770
rect 770 5760 780 5770
rect 820 5760 830 5770
rect 840 5760 860 5770
rect 1880 5760 1960 5770
rect 2210 5760 2240 5770
rect 2320 5760 2350 5770
rect 2370 5760 2390 5770
rect 2400 5760 2410 5770
rect 2450 5760 2590 5770
rect 2960 5760 3050 5770
rect 3100 5760 3120 5770
rect 3180 5760 3240 5770
rect 3950 5760 3960 5770
rect 4090 5760 4100 5770
rect 4510 5760 4520 5770
rect 4540 5760 4600 5770
rect 4680 5760 4710 5770
rect 4740 5760 4750 5770
rect 5320 5760 5340 5770
rect 6790 5760 6820 5770
rect 6990 5760 7010 5770
rect 7980 5760 7990 5770
rect 8380 5760 8390 5770
rect 8690 5760 8700 5770
rect 540 5750 580 5760
rect 640 5750 710 5760
rect 770 5750 790 5760
rect 810 5750 820 5760
rect 850 5750 870 5760
rect 1880 5750 1960 5760
rect 2210 5750 2220 5760
rect 2320 5750 2340 5760
rect 2350 5750 2560 5760
rect 2570 5750 2580 5760
rect 2970 5750 3040 5760
rect 3180 5750 3230 5760
rect 3970 5750 3980 5760
rect 4500 5750 4520 5760
rect 4550 5750 4560 5760
rect 4580 5750 4600 5760
rect 4640 5750 4650 5760
rect 4670 5750 4680 5760
rect 4750 5750 4770 5760
rect 5080 5750 5090 5760
rect 5310 5750 5330 5760
rect 6790 5750 6810 5760
rect 6990 5750 7000 5760
rect 7920 5750 7970 5760
rect 8420 5750 8430 5760
rect 8730 5750 8740 5760
rect 8840 5750 8850 5760
rect 8920 5750 8930 5760
rect 530 5740 540 5750
rect 610 5740 630 5750
rect 700 5740 750 5750
rect 780 5740 800 5750
rect 820 5740 830 5750
rect 860 5740 870 5750
rect 1890 5740 1960 5750
rect 2200 5740 2220 5750
rect 2310 5740 2320 5750
rect 2340 5740 2550 5750
rect 2960 5740 3030 5750
rect 3180 5740 3230 5750
rect 3760 5740 3770 5750
rect 3950 5740 4000 5750
rect 4350 5740 4370 5750
rect 4500 5740 4560 5750
rect 4590 5740 4600 5750
rect 4750 5740 4770 5750
rect 5310 5740 5330 5750
rect 6800 5740 6820 5750
rect 6980 5740 7000 5750
rect 7920 5740 7930 5750
rect 8270 5740 8280 5750
rect 8860 5740 8880 5750
rect 8890 5740 8910 5750
rect 590 5730 610 5740
rect 1900 5730 1960 5740
rect 2200 5730 2220 5740
rect 2300 5730 2330 5740
rect 2340 5730 2530 5740
rect 2960 5730 3010 5740
rect 3180 5730 3230 5740
rect 3750 5730 3800 5740
rect 4000 5730 4010 5740
rect 4350 5730 4360 5740
rect 4520 5730 4530 5740
rect 4580 5730 4600 5740
rect 5300 5730 5320 5740
rect 6810 5730 6820 5740
rect 6980 5730 6990 5740
rect 7850 5730 7870 5740
rect 7890 5730 7910 5740
rect 8240 5730 8250 5740
rect 560 5720 700 5730
rect 730 5720 760 5730
rect 1910 5720 1960 5730
rect 2200 5720 2210 5730
rect 2290 5720 2330 5730
rect 2350 5720 2530 5730
rect 2830 5720 2840 5730
rect 2950 5720 3000 5730
rect 3030 5720 3050 5730
rect 3180 5720 3230 5730
rect 3770 5720 3780 5730
rect 3810 5720 3820 5730
rect 4290 5720 4300 5730
rect 4340 5720 4350 5730
rect 4380 5720 4390 5730
rect 4400 5720 4410 5730
rect 4520 5720 4530 5730
rect 4590 5720 4610 5730
rect 5300 5720 5320 5730
rect 6810 5720 6820 5730
rect 6980 5720 6990 5730
rect 7790 5720 7800 5730
rect 7820 5720 7890 5730
rect 8180 5720 8190 5730
rect 8240 5720 8250 5730
rect 8390 5720 8400 5730
rect 8740 5720 8750 5730
rect 490 5710 550 5720
rect 630 5710 670 5720
rect 1910 5710 1950 5720
rect 2190 5710 2210 5720
rect 2280 5710 2310 5720
rect 2350 5710 2530 5720
rect 2820 5710 2930 5720
rect 2940 5710 3010 5720
rect 3020 5710 3040 5720
rect 3190 5710 3230 5720
rect 3790 5710 3800 5720
rect 3820 5710 3840 5720
rect 4280 5710 4310 5720
rect 4400 5710 4410 5720
rect 4560 5710 4660 5720
rect 4760 5710 4770 5720
rect 5070 5710 5080 5720
rect 5300 5710 5320 5720
rect 6820 5710 6830 5720
rect 6920 5710 6930 5720
rect 6980 5710 6990 5720
rect 7610 5710 7640 5720
rect 7750 5710 7770 5720
rect 7790 5710 7840 5720
rect 7860 5710 7890 5720
rect 8280 5710 8290 5720
rect 8430 5710 8440 5720
rect 8700 5710 8710 5720
rect 460 5700 510 5710
rect 630 5700 670 5710
rect 790 5700 800 5710
rect 1180 5700 1210 5710
rect 1930 5700 1960 5710
rect 2190 5700 2210 5710
rect 2280 5700 2300 5710
rect 2330 5700 2510 5710
rect 2810 5700 3030 5710
rect 3180 5700 3230 5710
rect 3820 5700 3840 5710
rect 4040 5700 4060 5710
rect 4230 5700 4250 5710
rect 4290 5700 4300 5710
rect 4320 5700 4340 5710
rect 4550 5700 4580 5710
rect 4600 5700 4630 5710
rect 4640 5700 4660 5710
rect 4710 5700 4730 5710
rect 4760 5700 4790 5710
rect 5300 5700 5310 5710
rect 6820 5700 6840 5710
rect 6960 5700 6990 5710
rect 7730 5700 7740 5710
rect 7750 5700 7800 5710
rect 8140 5700 8150 5710
rect 550 5690 560 5700
rect 630 5690 670 5700
rect 800 5690 810 5700
rect 1130 5690 1180 5700
rect 1940 5690 1960 5700
rect 1970 5690 1980 5700
rect 2190 5690 2200 5700
rect 2270 5690 2290 5700
rect 2330 5690 2480 5700
rect 2800 5690 2840 5700
rect 2880 5690 2900 5700
rect 2920 5690 3020 5700
rect 3180 5690 3240 5700
rect 4000 5690 4010 5700
rect 4270 5690 4280 5700
rect 4320 5690 4340 5700
rect 4550 5690 4570 5700
rect 4600 5690 4630 5700
rect 4680 5690 4760 5700
rect 4770 5690 4800 5700
rect 5290 5690 5310 5700
rect 6820 5690 6840 5700
rect 6980 5690 6990 5700
rect 7700 5690 7750 5700
rect 8110 5690 8120 5700
rect 8180 5690 8190 5700
rect 550 5680 560 5690
rect 620 5680 650 5690
rect 790 5680 810 5690
rect 1080 5680 1090 5690
rect 1100 5680 1140 5690
rect 1930 5680 1990 5690
rect 2180 5680 2210 5690
rect 2270 5680 2290 5690
rect 2320 5680 2470 5690
rect 2800 5680 2840 5690
rect 2920 5680 3020 5690
rect 3180 5680 3210 5690
rect 3220 5680 3240 5690
rect 4190 5680 4200 5690
rect 4250 5680 4270 5690
rect 4300 5680 4310 5690
rect 4570 5680 4640 5690
rect 4710 5680 4760 5690
rect 4790 5680 4800 5690
rect 6820 5680 6840 5690
rect 6980 5680 7000 5690
rect 7670 5680 7710 5690
rect 7720 5680 7740 5690
rect 7880 5680 7900 5690
rect 8040 5680 8050 5690
rect 8110 5680 8120 5690
rect 8180 5680 8190 5690
rect 8220 5680 8230 5690
rect 8400 5680 8410 5690
rect 540 5670 550 5680
rect 630 5670 650 5680
rect 790 5670 800 5680
rect 810 5670 830 5680
rect 1930 5670 1980 5680
rect 2180 5670 2200 5680
rect 2270 5670 2280 5680
rect 2300 5670 2380 5680
rect 2390 5670 2470 5680
rect 2800 5670 2820 5680
rect 2910 5670 2950 5680
rect 2960 5670 3010 5680
rect 3150 5670 3170 5680
rect 3180 5670 3210 5680
rect 3220 5670 3250 5680
rect 3900 5670 3910 5680
rect 4180 5670 4200 5680
rect 4290 5670 4310 5680
rect 4360 5670 4370 5680
rect 4410 5670 4420 5680
rect 4580 5670 4600 5680
rect 4610 5670 4630 5680
rect 4710 5670 4720 5680
rect 4740 5670 4770 5680
rect 5100 5670 5110 5680
rect 5290 5670 5300 5680
rect 6830 5670 6850 5680
rect 6970 5670 6990 5680
rect 7650 5670 7660 5680
rect 7690 5670 7710 5680
rect 7880 5670 7900 5680
rect 8110 5670 8120 5680
rect 8150 5670 8160 5680
rect 8250 5670 8260 5680
rect 8400 5670 8410 5680
rect 8440 5670 8450 5680
rect 620 5660 650 5670
rect 780 5660 800 5670
rect 1940 5660 1980 5670
rect 2170 5660 2190 5670
rect 2260 5660 2280 5670
rect 2300 5660 2380 5670
rect 2390 5660 2470 5670
rect 2800 5660 2820 5670
rect 2910 5660 2960 5670
rect 2970 5660 3010 5670
rect 3150 5660 3190 5670
rect 3200 5660 3250 5670
rect 3730 5660 3740 5670
rect 3890 5660 3900 5670
rect 4280 5660 4320 5670
rect 4350 5660 4360 5670
rect 4390 5660 4400 5670
rect 4410 5660 4420 5670
rect 4580 5660 4600 5670
rect 4750 5660 4780 5670
rect 5100 5660 5130 5670
rect 5290 5660 5300 5670
rect 6830 5660 6850 5670
rect 6940 5660 6990 5670
rect 7660 5660 7690 5670
rect 7890 5660 7900 5670
rect 8020 5660 8030 5670
rect 8060 5660 8070 5670
rect 8290 5660 8300 5670
rect 610 5650 660 5660
rect 760 5650 780 5660
rect 1960 5650 1980 5660
rect 2170 5650 2190 5660
rect 2260 5650 2270 5660
rect 2290 5650 2360 5660
rect 2420 5650 2480 5660
rect 2800 5650 2820 5660
rect 2970 5650 3010 5660
rect 3160 5650 3250 5660
rect 3710 5650 3720 5660
rect 3750 5650 3760 5660
rect 3810 5650 3820 5660
rect 3900 5650 3910 5660
rect 4210 5650 4220 5660
rect 4280 5650 4300 5660
rect 4330 5650 4340 5660
rect 4400 5650 4410 5660
rect 4580 5650 4600 5660
rect 4720 5650 4780 5660
rect 5290 5650 5300 5660
rect 5710 5650 5730 5660
rect 6830 5650 6850 5660
rect 6950 5650 6960 5660
rect 6980 5650 7000 5660
rect 7580 5650 7600 5660
rect 7630 5650 7650 5660
rect 7890 5650 7900 5660
rect 8290 5650 8300 5660
rect 8470 5650 8480 5660
rect 9990 5650 9990 5660
rect 530 5640 570 5650
rect 610 5640 660 5650
rect 1960 5640 1970 5650
rect 2160 5640 2180 5650
rect 2250 5640 2270 5650
rect 2290 5640 2350 5650
rect 2400 5640 2470 5650
rect 2730 5640 2760 5650
rect 2810 5640 2820 5650
rect 2980 5640 3010 5650
rect 3170 5640 3250 5650
rect 3740 5640 3750 5650
rect 3800 5640 3810 5650
rect 3870 5640 3880 5650
rect 3900 5640 3910 5650
rect 4210 5640 4240 5650
rect 4270 5640 4280 5650
rect 4330 5640 4340 5650
rect 4730 5640 4750 5650
rect 5070 5640 5100 5650
rect 5120 5640 5130 5650
rect 5280 5640 5290 5650
rect 5600 5640 5770 5650
rect 6840 5640 6850 5650
rect 6970 5640 6980 5650
rect 7570 5640 7620 5650
rect 8160 5640 8170 5650
rect 520 5630 620 5640
rect 630 5630 660 5640
rect 1940 5630 1950 5640
rect 1960 5630 1970 5640
rect 2110 5630 2140 5640
rect 2150 5630 2180 5640
rect 2250 5630 2260 5640
rect 2290 5630 2350 5640
rect 2440 5630 2470 5640
rect 2730 5630 2790 5640
rect 2810 5630 2830 5640
rect 3170 5630 3250 5640
rect 3710 5630 3720 5640
rect 3900 5630 3910 5640
rect 4090 5630 4100 5640
rect 4200 5630 4230 5640
rect 4260 5630 4290 5640
rect 5080 5630 5100 5640
rect 5280 5630 5290 5640
rect 5550 5630 5720 5640
rect 5760 5630 5790 5640
rect 5840 5630 5860 5640
rect 6840 5630 6860 5640
rect 6970 5630 6990 5640
rect 7510 5630 7580 5640
rect 8120 5630 8130 5640
rect 8160 5630 8170 5640
rect 8190 5630 8200 5640
rect 8230 5630 8240 5640
rect 520 5620 620 5630
rect 630 5620 660 5630
rect 730 5620 740 5630
rect 1940 5620 1950 5630
rect 1960 5620 2000 5630
rect 2030 5620 2050 5630
rect 2090 5620 2180 5630
rect 2250 5620 2260 5630
rect 2280 5620 2350 5630
rect 2420 5620 2470 5630
rect 2720 5620 2800 5630
rect 2820 5620 2850 5630
rect 3170 5620 3250 5630
rect 3810 5620 3820 5630
rect 3840 5620 3860 5630
rect 3900 5620 3910 5630
rect 4090 5620 4100 5630
rect 4220 5620 4230 5630
rect 4260 5620 4290 5630
rect 5110 5620 5120 5630
rect 5280 5620 5290 5630
rect 5540 5620 5600 5630
rect 5780 5620 5870 5630
rect 5940 5620 5950 5630
rect 6850 5620 6860 5630
rect 6960 5620 6990 5630
rect 7460 5620 7480 5630
rect 7490 5620 7530 5630
rect 7840 5620 7900 5630
rect 8030 5620 8040 5630
rect 8100 5620 8120 5630
rect 8230 5620 8240 5630
rect 8260 5620 8270 5630
rect 8410 5620 8420 5630
rect 520 5610 670 5620
rect 1950 5610 2010 5620
rect 2020 5610 2060 5620
rect 2110 5610 2180 5620
rect 2250 5610 2260 5620
rect 2270 5610 2350 5620
rect 2420 5610 2460 5620
rect 2720 5610 2810 5620
rect 2840 5610 2880 5620
rect 3160 5610 3240 5620
rect 3700 5610 3720 5620
rect 4120 5610 4130 5620
rect 4190 5610 4220 5620
rect 5070 5610 5090 5620
rect 5280 5610 5290 5620
rect 5510 5610 5580 5620
rect 5820 5610 5880 5620
rect 5890 5610 5960 5620
rect 5990 5610 6060 5620
rect 6200 5610 6270 5620
rect 6280 5610 6290 5620
rect 6320 5610 6430 5620
rect 6440 5610 6450 5620
rect 6850 5610 6870 5620
rect 6960 5610 6980 5620
rect 7440 5610 7480 5620
rect 7490 5610 7500 5620
rect 7810 5610 7820 5620
rect 7900 5610 7910 5620
rect 8030 5610 8040 5620
rect 8070 5610 8080 5620
rect 8300 5610 8310 5620
rect 8350 5610 8360 5620
rect 8460 5610 8470 5620
rect 9990 5610 9990 5620
rect 510 5600 670 5610
rect 700 5600 710 5610
rect 1950 5600 2030 5610
rect 2040 5600 2050 5610
rect 2110 5600 2180 5610
rect 2240 5600 2350 5610
rect 2410 5600 2450 5610
rect 2720 5600 2820 5610
rect 2870 5600 2890 5610
rect 2910 5600 2940 5610
rect 3170 5600 3250 5610
rect 3680 5600 3690 5610
rect 4190 5600 4210 5610
rect 4260 5600 4290 5610
rect 5280 5600 5290 5610
rect 5480 5600 5490 5610
rect 5500 5600 5560 5610
rect 5840 5600 6070 5610
rect 6170 5600 6530 5610
rect 6860 5600 6880 5610
rect 6970 5600 6980 5610
rect 7430 5600 7450 5610
rect 7910 5600 7920 5610
rect 8030 5600 8040 5610
rect 8320 5600 8330 5610
rect 9010 5600 9050 5610
rect 9990 5600 9990 5610
rect 510 5590 560 5600
rect 570 5590 620 5600
rect 630 5590 680 5600
rect 690 5590 700 5600
rect 1950 5590 2050 5600
rect 2080 5590 2090 5600
rect 2110 5590 2180 5600
rect 2240 5590 2350 5600
rect 2380 5590 2390 5600
rect 2400 5590 2440 5600
rect 2660 5590 2680 5600
rect 2710 5590 2840 5600
rect 2880 5590 2940 5600
rect 3160 5590 3250 5600
rect 3420 5590 3430 5600
rect 4100 5590 4110 5600
rect 4150 5590 4170 5600
rect 4180 5590 4190 5600
rect 4310 5590 4330 5600
rect 5270 5590 5280 5600
rect 5470 5590 5520 5600
rect 5870 5590 6090 5600
rect 6150 5590 6320 5600
rect 6420 5590 6610 5600
rect 6860 5590 6880 5600
rect 6960 5590 6980 5600
rect 7300 5590 7320 5600
rect 7420 5590 7430 5600
rect 8170 5590 8180 5600
rect 8200 5590 8210 5600
rect 8240 5590 8250 5600
rect 8270 5590 8280 5600
rect 9990 5590 9990 5600
rect 510 5580 600 5590
rect 610 5580 620 5590
rect 630 5580 670 5590
rect 1950 5580 2090 5590
rect 2100 5580 2180 5590
rect 2240 5580 2340 5590
rect 2380 5580 2430 5590
rect 2690 5580 2850 5590
rect 2900 5580 2950 5590
rect 3160 5580 3250 5590
rect 3430 5580 3450 5590
rect 3770 5580 3780 5590
rect 3820 5580 3830 5590
rect 4110 5580 4130 5590
rect 4150 5580 4160 5590
rect 4240 5580 4250 5590
rect 4290 5580 4320 5590
rect 5090 5580 5100 5590
rect 5270 5580 5280 5590
rect 5460 5580 5490 5590
rect 5880 5580 6090 5590
rect 6110 5580 6120 5590
rect 6130 5580 6300 5590
rect 6460 5580 6620 5590
rect 6870 5580 6880 5590
rect 6960 5580 6980 5590
rect 7300 5580 7310 5590
rect 7400 5580 7410 5590
rect 7720 5580 7730 5590
rect 7750 5580 7760 5590
rect 7840 5580 7880 5590
rect 7920 5580 7930 5590
rect 8270 5580 8280 5590
rect 510 5570 600 5580
rect 630 5570 660 5580
rect 1950 5570 2100 5580
rect 2110 5570 2170 5580
rect 2240 5570 2340 5580
rect 2380 5570 2420 5580
rect 2690 5570 2860 5580
rect 2920 5570 2960 5580
rect 3160 5570 3240 5580
rect 3680 5570 3690 5580
rect 3810 5570 3820 5580
rect 3860 5570 3870 5580
rect 4100 5570 4120 5580
rect 4160 5570 4170 5580
rect 4240 5570 4280 5580
rect 5090 5570 5100 5580
rect 5270 5570 5280 5580
rect 5460 5570 5490 5580
rect 5900 5570 6240 5580
rect 6250 5570 6270 5580
rect 6530 5570 6540 5580
rect 6550 5570 6620 5580
rect 6870 5570 6880 5580
rect 6970 5570 6980 5580
rect 7290 5570 7320 5580
rect 7360 5570 7370 5580
rect 7680 5570 7690 5580
rect 7920 5570 7930 5580
rect 8040 5570 8050 5580
rect 8080 5570 8090 5580
rect 8330 5570 8340 5580
rect 8960 5570 8970 5580
rect 510 5560 580 5570
rect 1960 5560 2170 5570
rect 2240 5560 2340 5570
rect 2360 5560 2400 5570
rect 2680 5560 2690 5570
rect 2700 5560 2870 5570
rect 2930 5560 2980 5570
rect 3170 5560 3240 5570
rect 3460 5560 3470 5570
rect 3840 5560 3850 5570
rect 4110 5560 4120 5570
rect 4160 5560 4170 5570
rect 4190 5560 4200 5570
rect 4210 5560 4300 5570
rect 4490 5560 4500 5570
rect 5270 5560 5280 5570
rect 5450 5560 5510 5570
rect 5940 5560 6220 5570
rect 6580 5560 6670 5570
rect 6960 5560 6970 5570
rect 7300 5560 7310 5570
rect 7360 5560 7370 5570
rect 7660 5560 7670 5570
rect 7880 5560 7890 5570
rect 8040 5560 8050 5570
rect 8080 5560 8090 5570
rect 8870 5560 8890 5570
rect 500 5550 580 5560
rect 600 5550 610 5560
rect 650 5550 660 5560
rect 1970 5550 2100 5560
rect 2110 5550 2170 5560
rect 2240 5550 2350 5560
rect 2370 5550 2400 5560
rect 2700 5550 2870 5560
rect 2950 5550 2990 5560
rect 3170 5550 3230 5560
rect 3660 5550 3680 5560
rect 3740 5550 3750 5560
rect 3790 5550 3800 5560
rect 3830 5550 3840 5560
rect 3910 5550 3920 5560
rect 4110 5550 4150 5560
rect 4160 5550 4170 5560
rect 4190 5550 4200 5560
rect 4210 5550 4270 5560
rect 4280 5550 4300 5560
rect 4330 5550 4350 5560
rect 4370 5550 4380 5560
rect 4480 5550 4500 5560
rect 5090 5550 5100 5560
rect 5260 5550 5270 5560
rect 5450 5550 5500 5560
rect 5940 5550 6200 5560
rect 6590 5550 6670 5560
rect 6880 5550 6890 5560
rect 6960 5550 6970 5560
rect 7260 5550 7300 5560
rect 7320 5550 7330 5560
rect 7650 5550 7660 5560
rect 7790 5550 7800 5560
rect 7830 5550 7840 5560
rect 7880 5550 7890 5560
rect 8210 5550 8220 5560
rect 8240 5550 8250 5560
rect 8950 5550 8960 5560
rect 510 5540 570 5550
rect 600 5540 610 5550
rect 620 5540 630 5550
rect 1960 5540 2160 5550
rect 2240 5540 2410 5550
rect 2690 5540 2870 5550
rect 2960 5540 2990 5550
rect 3160 5540 3230 5550
rect 3810 5540 3820 5550
rect 4110 5540 4140 5550
rect 4150 5540 4160 5550
rect 4230 5540 4250 5550
rect 4280 5540 4300 5550
rect 4330 5540 4340 5550
rect 4350 5540 4370 5550
rect 5090 5540 5120 5550
rect 5260 5540 5270 5550
rect 5430 5540 5490 5550
rect 5550 5540 5600 5550
rect 5950 5540 6080 5550
rect 6090 5540 6180 5550
rect 6600 5540 6670 5550
rect 6880 5540 6890 5550
rect 7260 5540 7280 5550
rect 7300 5540 7310 5550
rect 7710 5540 7720 5550
rect 7830 5540 7840 5550
rect 7880 5540 7890 5550
rect 7930 5540 7940 5550
rect 8140 5540 8150 5550
rect 8860 5540 8870 5550
rect 8900 5540 8910 5550
rect 500 5530 520 5540
rect 540 5530 560 5540
rect 600 5530 620 5540
rect 640 5530 650 5540
rect 1970 5530 2160 5540
rect 2240 5530 2390 5540
rect 2690 5530 2850 5540
rect 2860 5530 2870 5540
rect 2900 5530 2920 5540
rect 2970 5530 3030 5540
rect 3160 5530 3220 5540
rect 3770 5530 3780 5540
rect 4110 5530 4160 5540
rect 4180 5530 4190 5540
rect 4260 5530 4270 5540
rect 4290 5530 4310 5540
rect 4350 5530 4360 5540
rect 5090 5530 5110 5540
rect 5260 5530 5270 5540
rect 5420 5530 5480 5540
rect 5510 5530 5610 5540
rect 5970 5530 6170 5540
rect 6600 5530 6610 5540
rect 6620 5530 6680 5540
rect 6880 5530 6890 5540
rect 6970 5530 6980 5540
rect 7290 5530 7300 5540
rect 7330 5530 7340 5540
rect 7550 5530 7560 5540
rect 7600 5530 7610 5540
rect 7650 5530 7660 5540
rect 7880 5530 7890 5540
rect 7930 5530 7940 5540
rect 8050 5530 8060 5540
rect 8090 5530 8100 5540
rect 8780 5530 8800 5540
rect 8860 5530 8870 5540
rect 500 5520 510 5530
rect 530 5520 550 5530
rect 610 5520 620 5530
rect 640 5520 650 5530
rect 930 5520 940 5530
rect 1970 5520 2160 5530
rect 2240 5520 2390 5530
rect 2700 5520 2840 5530
rect 2900 5520 2940 5530
rect 2980 5520 3050 5530
rect 3160 5520 3200 5530
rect 3210 5520 3220 5530
rect 3660 5520 3670 5530
rect 3730 5520 3740 5530
rect 3750 5520 3760 5530
rect 3790 5520 3800 5530
rect 4130 5520 4160 5530
rect 4200 5520 4220 5530
rect 4250 5520 4280 5530
rect 4350 5520 4370 5530
rect 5260 5520 5270 5530
rect 5410 5520 5470 5530
rect 5480 5520 5630 5530
rect 5960 5520 6050 5530
rect 6100 5520 6160 5530
rect 6600 5520 6710 5530
rect 6880 5520 6890 5530
rect 7290 5520 7310 5530
rect 7330 5520 7340 5530
rect 7370 5520 7380 5530
rect 7520 5520 7530 5530
rect 7650 5520 7660 5530
rect 7880 5520 7890 5530
rect 7930 5520 7940 5530
rect 8050 5520 8060 5530
rect 8090 5520 8100 5530
rect 8760 5520 8770 5530
rect 460 5510 480 5520
rect 490 5510 500 5520
rect 610 5510 620 5520
rect 940 5510 950 5520
rect 1970 5510 2160 5520
rect 2240 5510 2270 5520
rect 2280 5510 2370 5520
rect 2620 5510 2630 5520
rect 2640 5510 2650 5520
rect 2700 5510 2840 5520
rect 2910 5510 2940 5520
rect 2990 5510 3060 5520
rect 3160 5510 3200 5520
rect 3210 5510 3220 5520
rect 3780 5510 3790 5520
rect 4130 5510 4150 5520
rect 4190 5510 4260 5520
rect 4300 5510 4330 5520
rect 4360 5510 4370 5520
rect 5110 5510 5120 5520
rect 5410 5510 5670 5520
rect 5960 5510 6050 5520
rect 6110 5510 6160 5520
rect 6600 5510 6730 5520
rect 6960 5510 6970 5520
rect 7250 5510 7270 5520
rect 7630 5510 7640 5520
rect 7650 5510 7660 5520
rect 7800 5510 7810 5520
rect 7880 5510 7900 5520
rect 7930 5510 7940 5520
rect 8090 5510 8100 5520
rect 8950 5510 8960 5520
rect 8990 5510 9000 5520
rect 350 5500 430 5510
rect 590 5500 600 5510
rect 1970 5500 2160 5510
rect 2240 5500 2280 5510
rect 2290 5500 2370 5510
rect 2610 5500 2660 5510
rect 2690 5500 2790 5510
rect 2910 5500 2940 5510
rect 3000 5500 3060 5510
rect 3150 5500 3200 5510
rect 3210 5500 3220 5510
rect 3660 5500 3670 5510
rect 3720 5500 3730 5510
rect 3740 5500 3750 5510
rect 4090 5500 4120 5510
rect 4140 5500 4150 5510
rect 4200 5500 4210 5510
rect 4230 5500 4240 5510
rect 4300 5500 4330 5510
rect 4360 5500 4390 5510
rect 4430 5500 4460 5510
rect 5100 5500 5120 5510
rect 5250 5500 5260 5510
rect 5410 5500 5680 5510
rect 5960 5500 6040 5510
rect 6120 5500 6160 5510
rect 6590 5500 6730 5510
rect 6890 5500 6900 5510
rect 6960 5500 6970 5510
rect 7230 5500 7280 5510
rect 7500 5500 7510 5510
rect 7630 5500 7640 5510
rect 7720 5500 7730 5510
rect 7740 5500 7750 5510
rect 7800 5500 7810 5510
rect 7840 5500 7850 5510
rect 7890 5500 7900 5510
rect 8720 5500 8730 5510
rect 8910 5500 8920 5510
rect 8950 5500 8960 5510
rect 9110 5500 9120 5510
rect 370 5490 400 5500
rect 1980 5490 2160 5500
rect 2240 5490 2290 5500
rect 2300 5490 2370 5500
rect 2600 5490 2670 5500
rect 2690 5490 2730 5500
rect 2740 5490 2750 5500
rect 2920 5490 2940 5500
rect 3010 5490 3070 5500
rect 3140 5490 3200 5500
rect 3680 5490 3690 5500
rect 3710 5490 3730 5500
rect 4090 5490 4100 5500
rect 4120 5490 4150 5500
rect 4190 5490 4200 5500
rect 4220 5490 4250 5500
rect 4360 5490 4380 5500
rect 4430 5490 4460 5500
rect 5100 5490 5110 5500
rect 5250 5490 5260 5500
rect 5410 5490 5520 5500
rect 5540 5490 5670 5500
rect 5960 5490 6020 5500
rect 6120 5490 6160 5500
rect 6540 5490 6730 5500
rect 6950 5490 6960 5500
rect 7220 5490 7260 5500
rect 7270 5490 7280 5500
rect 7300 5490 7310 5500
rect 7330 5490 7340 5500
rect 7380 5490 7390 5500
rect 7500 5490 7510 5500
rect 7630 5490 7640 5500
rect 8760 5490 8770 5500
rect 8870 5490 8880 5500
rect 9040 5490 9050 5500
rect 400 5480 420 5490
rect 560 5480 570 5490
rect 590 5480 600 5490
rect 960 5480 970 5490
rect 1980 5480 2160 5490
rect 2240 5480 2340 5490
rect 2590 5480 2680 5490
rect 2690 5480 2730 5490
rect 3020 5480 3080 5490
rect 3130 5480 3200 5490
rect 3650 5480 3660 5490
rect 4000 5480 4010 5490
rect 4080 5480 4090 5490
rect 4130 5480 4140 5490
rect 4180 5480 4190 5490
rect 4430 5480 4470 5490
rect 4500 5480 4510 5490
rect 5250 5480 5260 5490
rect 5410 5480 5520 5490
rect 5960 5480 6000 5490
rect 6010 5480 6020 5490
rect 6120 5480 6150 5490
rect 6530 5480 6730 5490
rect 6960 5480 6970 5490
rect 7230 5480 7300 5490
rect 7310 5480 7320 5490
rect 7380 5480 7390 5490
rect 7590 5480 7600 5490
rect 7880 5480 7890 5490
rect 7930 5480 7940 5490
rect 8870 5480 8880 5490
rect 430 5470 440 5480
rect 550 5470 570 5480
rect 1980 5470 2160 5480
rect 2240 5470 2340 5480
rect 2600 5470 2730 5480
rect 3040 5470 3080 5480
rect 3110 5470 3190 5480
rect 3580 5470 3620 5480
rect 3650 5470 3660 5480
rect 4050 5470 4070 5480
rect 4080 5470 4090 5480
rect 4160 5470 4170 5480
rect 4250 5470 4260 5480
rect 4270 5470 4320 5480
rect 4440 5470 4470 5480
rect 4610 5470 4620 5480
rect 5400 5470 5500 5480
rect 5960 5470 6000 5480
rect 6120 5470 6150 5480
rect 6530 5470 6730 5480
rect 6950 5470 6970 5480
rect 7230 5470 7240 5480
rect 7250 5470 7260 5480
rect 7280 5470 7300 5480
rect 7380 5470 7390 5480
rect 7580 5470 7590 5480
rect 7660 5470 7670 5480
rect 7870 5470 7880 5480
rect 8690 5470 8700 5480
rect 8960 5470 8970 5480
rect 9000 5470 9010 5480
rect 440 5460 450 5470
rect 1990 5460 2160 5470
rect 2240 5460 2350 5470
rect 2600 5460 2740 5470
rect 3040 5460 3170 5470
rect 3590 5460 3600 5470
rect 4080 5460 4110 5470
rect 4150 5460 4160 5470
rect 4180 5460 4190 5470
rect 4270 5460 4380 5470
rect 4450 5460 4460 5470
rect 4490 5460 4520 5470
rect 4530 5460 4550 5470
rect 4570 5460 4590 5470
rect 4620 5460 4630 5470
rect 4700 5460 4720 5470
rect 5080 5460 5100 5470
rect 5400 5460 5490 5470
rect 5960 5460 5990 5470
rect 6130 5460 6160 5470
rect 6530 5460 6740 5470
rect 6900 5460 6910 5470
rect 6930 5460 6960 5470
rect 7230 5460 7250 5470
rect 7280 5460 7290 5470
rect 7370 5460 7380 5470
rect 7620 5460 7630 5470
rect 7710 5460 7720 5470
rect 7810 5460 7820 5470
rect 7920 5460 7930 5470
rect 8690 5460 8700 5470
rect 8730 5460 8740 5470
rect 8880 5460 8890 5470
rect 8920 5460 8930 5470
rect 8960 5460 8970 5470
rect 2010 5450 2160 5460
rect 2240 5450 2360 5460
rect 2630 5450 2760 5460
rect 3010 5450 3160 5460
rect 3590 5450 3600 5460
rect 4080 5450 4100 5460
rect 4120 5450 4150 5460
rect 4270 5450 4290 5460
rect 4300 5450 4340 5460
rect 4350 5450 4380 5460
rect 4480 5450 4520 5460
rect 4580 5450 4590 5460
rect 4660 5450 4750 5460
rect 5100 5450 5110 5460
rect 5240 5450 5250 5460
rect 5400 5450 5470 5460
rect 5600 5450 5650 5460
rect 5960 5450 5990 5460
rect 6130 5450 6160 5460
rect 6520 5450 6730 5460
rect 6940 5450 6960 5460
rect 7200 5450 7210 5460
rect 7220 5450 7250 5460
rect 7340 5450 7350 5460
rect 7360 5450 7370 5460
rect 7510 5450 7520 5460
rect 7610 5450 7620 5460
rect 7810 5450 7820 5460
rect 7910 5450 7920 5460
rect 8770 5450 8780 5460
rect 8810 5450 8830 5460
rect 8870 5450 8890 5460
rect 440 5440 450 5450
rect 2010 5440 2160 5450
rect 2240 5440 2360 5450
rect 2630 5440 2780 5450
rect 3020 5440 3160 5450
rect 4070 5440 4080 5450
rect 4110 5440 4120 5450
rect 4270 5440 4310 5450
rect 4320 5440 4340 5450
rect 4350 5440 4360 5450
rect 4370 5440 4420 5450
rect 4470 5440 4520 5450
rect 4550 5440 4590 5450
rect 4620 5440 4630 5450
rect 4650 5440 4660 5450
rect 4670 5440 4700 5450
rect 4710 5440 4730 5450
rect 5100 5440 5110 5450
rect 5240 5440 5250 5450
rect 5400 5440 5450 5450
rect 5580 5440 5650 5450
rect 5950 5440 5990 5450
rect 6130 5440 6160 5450
rect 6530 5440 6730 5450
rect 6940 5440 6950 5450
rect 7190 5440 7200 5450
rect 7220 5440 7240 5450
rect 7600 5440 7610 5450
rect 7710 5440 7720 5450
rect 8620 5440 8630 5450
rect 8660 5440 8670 5450
rect 8770 5440 8780 5450
rect 8880 5440 8890 5450
rect 9060 5440 9070 5450
rect 9110 5440 9120 5450
rect 440 5430 450 5440
rect 570 5430 580 5440
rect 2020 5430 2160 5440
rect 2240 5430 2360 5440
rect 2680 5430 2730 5440
rect 2740 5430 2760 5440
rect 2770 5430 2790 5440
rect 2820 5430 2830 5440
rect 3030 5430 3050 5440
rect 3060 5430 3150 5440
rect 4330 5430 4340 5440
rect 4400 5430 4410 5440
rect 4460 5430 4470 5440
rect 4480 5430 4520 5440
rect 4550 5430 4580 5440
rect 4600 5430 4630 5440
rect 4700 5430 4720 5440
rect 4740 5430 4760 5440
rect 5080 5430 5110 5440
rect 5400 5430 5450 5440
rect 5570 5430 5580 5440
rect 5950 5430 5980 5440
rect 6130 5430 6150 5440
rect 6600 5430 6730 5440
rect 6900 5430 6910 5440
rect 7180 5430 7190 5440
rect 7210 5430 7250 5440
rect 7670 5430 7680 5440
rect 7710 5430 7720 5440
rect 7740 5430 7750 5440
rect 7870 5430 7880 5440
rect 8740 5430 8750 5440
rect 8930 5430 8940 5440
rect 8970 5430 8980 5440
rect 440 5420 450 5430
rect 2020 5420 2050 5430
rect 2060 5420 2160 5430
rect 2240 5420 2370 5430
rect 2700 5420 2720 5430
rect 2740 5420 2770 5430
rect 2820 5420 2830 5430
rect 3040 5420 3070 5430
rect 4340 5420 4350 5430
rect 4470 5420 4480 5430
rect 4490 5420 4550 5430
rect 4570 5420 4590 5430
rect 4610 5420 4630 5430
rect 4670 5420 4710 5430
rect 4730 5420 4780 5430
rect 5110 5420 5120 5430
rect 5420 5420 5440 5430
rect 5950 5420 5980 5430
rect 6130 5420 6160 5430
rect 6610 5420 6730 5430
rect 6900 5420 6910 5430
rect 6950 5420 6960 5430
rect 7180 5420 7210 5430
rect 7230 5420 7260 5430
rect 7300 5420 7310 5430
rect 7670 5420 7680 5430
rect 8400 5420 8410 5430
rect 8460 5420 8470 5430
rect 8700 5420 8710 5430
rect 8820 5420 8830 5430
rect 8930 5420 8940 5430
rect 8980 5420 8990 5430
rect 9550 5420 9560 5430
rect 560 5410 570 5420
rect 2020 5410 2040 5420
rect 2050 5410 2160 5420
rect 2240 5410 2360 5420
rect 2810 5410 2830 5420
rect 3050 5410 3070 5420
rect 4090 5410 4100 5420
rect 4310 5410 4340 5420
rect 4400 5410 4410 5420
rect 4460 5410 4470 5420
rect 4480 5410 4520 5420
rect 4570 5410 4600 5420
rect 4630 5410 4660 5420
rect 4680 5410 4770 5420
rect 5080 5410 5090 5420
rect 5100 5410 5110 5420
rect 5410 5410 5440 5420
rect 5940 5410 5970 5420
rect 6130 5410 6160 5420
rect 6630 5410 6720 5420
rect 6900 5410 6910 5420
rect 6960 5410 6970 5420
rect 7180 5410 7200 5420
rect 7240 5410 7260 5420
rect 7280 5410 7290 5420
rect 7560 5410 7570 5420
rect 8370 5410 8380 5420
rect 8700 5410 8710 5420
rect 8780 5410 8790 5420
rect 9080 5410 9090 5420
rect 410 5400 430 5410
rect 560 5400 570 5410
rect 760 5400 770 5410
rect 2020 5400 2040 5410
rect 2060 5400 2170 5410
rect 2240 5400 2360 5410
rect 2800 5400 2820 5410
rect 3580 5400 3590 5410
rect 4090 5400 4100 5410
rect 4230 5400 4240 5410
rect 4460 5400 4470 5410
rect 4520 5400 4540 5410
rect 4560 5400 4580 5410
rect 4590 5400 4610 5410
rect 4620 5400 4750 5410
rect 5090 5400 5100 5410
rect 5400 5400 5430 5410
rect 5940 5400 5970 5410
rect 6130 5400 6160 5410
rect 6660 5400 6720 5410
rect 6900 5400 6910 5410
rect 6930 5400 6970 5410
rect 7190 5400 7200 5410
rect 7240 5400 7290 5410
rect 7520 5400 7530 5410
rect 7560 5400 7580 5410
rect 7770 5400 7780 5410
rect 8350 5400 8360 5410
rect 8480 5400 8490 5410
rect 8520 5400 8530 5410
rect 8670 5400 8680 5410
rect 9060 5400 9070 5410
rect 400 5390 410 5400
rect 510 5390 520 5400
rect 560 5390 570 5400
rect 2040 5390 2050 5400
rect 2060 5390 2170 5400
rect 2240 5390 2360 5400
rect 4220 5390 4240 5400
rect 4410 5390 4440 5400
rect 4450 5390 4460 5400
rect 4510 5390 4520 5400
rect 4560 5390 4590 5400
rect 4600 5390 4630 5400
rect 4650 5390 4750 5400
rect 5080 5390 5090 5400
rect 5380 5390 5400 5400
rect 5940 5390 5970 5400
rect 6130 5390 6160 5400
rect 6670 5390 6720 5400
rect 6900 5390 6910 5400
rect 7190 5390 7210 5400
rect 7240 5390 7250 5400
rect 7260 5390 7290 5400
rect 7520 5390 7530 5400
rect 7560 5390 7570 5400
rect 7580 5390 7590 5400
rect 7640 5390 7650 5400
rect 7680 5390 7690 5400
rect 7730 5390 7740 5400
rect 8420 5390 8440 5400
rect 8750 5390 8760 5400
rect 8940 5390 8950 5400
rect 9480 5390 9490 5400
rect 9520 5390 9530 5400
rect 380 5380 390 5390
rect 480 5380 500 5390
rect 540 5380 560 5390
rect 2030 5380 2080 5390
rect 2090 5380 2160 5390
rect 2240 5380 2370 5390
rect 3800 5380 3810 5390
rect 4080 5380 4100 5390
rect 4470 5380 4480 5390
rect 4490 5380 4510 5390
rect 4560 5380 4620 5390
rect 4640 5380 4650 5390
rect 4680 5380 4710 5390
rect 5370 5380 5380 5390
rect 5940 5380 5970 5390
rect 6130 5380 6160 5390
rect 6690 5380 6730 5390
rect 6930 5380 6940 5390
rect 7200 5380 7210 5390
rect 7240 5380 7260 5390
rect 7280 5380 7300 5390
rect 7590 5380 7600 5390
rect 7700 5380 7710 5390
rect 8390 5380 8400 5390
rect 8710 5380 8720 5390
rect 8790 5380 8800 5390
rect 8940 5380 8950 5390
rect 9530 5380 9550 5390
rect 360 5370 370 5380
rect 490 5370 500 5380
rect 530 5370 560 5380
rect 2020 5370 2080 5380
rect 2110 5370 2170 5380
rect 2250 5370 2360 5380
rect 3570 5370 3580 5380
rect 3800 5370 3820 5380
rect 4080 5370 4100 5380
rect 4180 5370 4190 5380
rect 4460 5370 4490 5380
rect 4560 5370 4590 5380
rect 4620 5370 4630 5380
rect 4660 5370 4700 5380
rect 5080 5370 5090 5380
rect 5230 5370 5240 5380
rect 5380 5370 5390 5380
rect 5400 5370 5410 5380
rect 5940 5370 5970 5380
rect 6130 5370 6160 5380
rect 6700 5370 6740 5380
rect 6920 5370 6950 5380
rect 7220 5370 7260 5380
rect 7290 5370 7300 5380
rect 7310 5370 7330 5380
rect 7600 5370 7610 5380
rect 8450 5370 8460 5380
rect 8570 5370 8590 5380
rect 8640 5370 8650 5380
rect 8710 5370 8720 5380
rect 8890 5370 8900 5380
rect 330 5360 340 5370
rect 450 5360 530 5370
rect 2020 5360 2030 5370
rect 2040 5360 2080 5370
rect 2110 5360 2170 5370
rect 2250 5360 2360 5370
rect 4170 5360 4190 5370
rect 4440 5360 4460 5370
rect 4520 5360 4540 5370
rect 4650 5360 4700 5370
rect 5080 5360 5090 5370
rect 5230 5360 5240 5370
rect 5380 5360 5420 5370
rect 5930 5360 5970 5370
rect 6140 5360 6160 5370
rect 6720 5360 6760 5370
rect 6930 5360 6950 5370
rect 7220 5360 7280 5370
rect 7290 5360 7320 5370
rect 7630 5360 7640 5370
rect 8350 5360 8360 5370
rect 8390 5360 8400 5370
rect 8570 5360 8580 5370
rect 8680 5360 8690 5370
rect 9440 5360 9450 5370
rect 300 5350 330 5360
rect 450 5350 540 5360
rect 2050 5350 2060 5360
rect 2080 5350 2110 5360
rect 2120 5350 2170 5360
rect 2250 5350 2360 5360
rect 3880 5350 3890 5360
rect 4100 5350 4120 5360
rect 4160 5350 4190 5360
rect 4470 5350 4490 5360
rect 4510 5350 4520 5360
rect 4640 5350 4690 5360
rect 4720 5350 4730 5360
rect 5370 5350 5390 5360
rect 5520 5350 5530 5360
rect 5930 5350 5970 5360
rect 6140 5350 6160 5360
rect 6720 5350 6760 5360
rect 6930 5350 6950 5360
rect 7250 5350 7270 5360
rect 7290 5350 7330 5360
rect 8280 5350 8290 5360
rect 8430 5350 8440 5360
rect 8530 5350 8540 5360
rect 8600 5350 8610 5360
rect 8720 5350 8730 5360
rect 8760 5350 8770 5360
rect 9280 5350 9290 5360
rect 9360 5350 9370 5360
rect 9410 5350 9420 5360
rect 260 5340 270 5350
rect 410 5340 540 5350
rect 2090 5340 2120 5350
rect 2130 5340 2170 5350
rect 2250 5340 2370 5350
rect 3560 5340 3570 5350
rect 4080 5340 4110 5350
rect 4120 5340 4140 5350
rect 4490 5340 4510 5350
rect 4570 5340 4580 5350
rect 4620 5340 4700 5350
rect 4720 5340 4730 5350
rect 5080 5340 5090 5350
rect 5360 5340 5370 5350
rect 5440 5340 5520 5350
rect 5570 5340 5580 5350
rect 5930 5340 5960 5350
rect 6150 5340 6170 5350
rect 6730 5340 6750 5350
rect 6910 5340 6940 5350
rect 7260 5340 7270 5350
rect 7280 5340 7310 5350
rect 7320 5340 7340 5350
rect 8160 5340 8170 5350
rect 8400 5340 8410 5350
rect 8610 5340 8620 5350
rect 8720 5340 8730 5350
rect 8800 5340 8810 5350
rect 8830 5340 8840 5350
rect 9270 5340 9280 5350
rect 250 5330 260 5340
rect 350 5330 560 5340
rect 2090 5330 2110 5340
rect 2130 5330 2170 5340
rect 2250 5330 2360 5340
rect 4100 5330 4140 5340
rect 4450 5330 4460 5340
rect 4490 5330 4510 5340
rect 4560 5330 4690 5340
rect 4720 5330 4730 5340
rect 4750 5330 4780 5340
rect 5080 5330 5090 5340
rect 5350 5330 5410 5340
rect 5460 5330 5510 5340
rect 5600 5330 5610 5340
rect 5870 5330 5900 5340
rect 5920 5330 5940 5340
rect 6150 5330 6170 5340
rect 6740 5330 6760 5340
rect 6910 5330 6940 5340
rect 7280 5330 7290 5340
rect 8290 5330 8300 5340
rect 9320 5330 9330 5340
rect 9340 5330 9350 5340
rect 310 5320 570 5330
rect 2060 5320 2080 5330
rect 2090 5320 2110 5330
rect 2130 5320 2170 5330
rect 2250 5320 2370 5330
rect 4110 5320 4140 5330
rect 4500 5320 4520 5330
rect 4580 5320 4600 5330
rect 4630 5320 4650 5330
rect 4710 5320 4730 5330
rect 4750 5320 4760 5330
rect 5090 5320 5130 5330
rect 5460 5320 5500 5330
rect 5640 5320 5660 5330
rect 5870 5320 5940 5330
rect 6150 5320 6170 5330
rect 6750 5320 6780 5330
rect 6910 5320 6950 5330
rect 7270 5320 7280 5330
rect 7310 5320 7320 5330
rect 8100 5320 8110 5330
rect 8540 5320 8550 5330
rect 9260 5320 9270 5330
rect 9420 5320 9430 5330
rect 9450 5320 9460 5330
rect 300 5310 570 5320
rect 2070 5310 2100 5320
rect 2130 5310 2170 5320
rect 2250 5310 2370 5320
rect 4110 5310 4130 5320
rect 4570 5310 4590 5320
rect 4600 5310 4610 5320
rect 4640 5310 4650 5320
rect 4720 5310 4730 5320
rect 4760 5310 4770 5320
rect 5080 5310 5130 5320
rect 5150 5310 5160 5320
rect 5220 5310 5230 5320
rect 5670 5310 5700 5320
rect 5860 5310 5930 5320
rect 6150 5310 6170 5320
rect 6790 5310 6800 5320
rect 6920 5310 6940 5320
rect 7260 5310 7270 5320
rect 8110 5310 8120 5320
rect 8580 5310 8590 5320
rect 8690 5310 8700 5320
rect 9130 5310 9150 5320
rect 210 5300 220 5310
rect 260 5300 560 5310
rect 2080 5300 2090 5310
rect 2140 5300 2180 5310
rect 2250 5300 2370 5310
rect 4600 5300 4620 5310
rect 4660 5300 4680 5310
rect 4700 5300 4720 5310
rect 5090 5300 5110 5310
rect 5120 5300 5130 5310
rect 5220 5300 5230 5310
rect 5680 5300 5700 5310
rect 5840 5300 5930 5310
rect 6160 5300 6180 5310
rect 6570 5300 6640 5310
rect 6790 5300 6810 5310
rect 6910 5300 6930 5310
rect 7230 5300 7240 5310
rect 7260 5300 7270 5310
rect 8000 5300 8010 5310
rect 8030 5300 8040 5310
rect 8420 5300 8430 5310
rect 8470 5300 8480 5310
rect 9120 5300 9130 5310
rect 9150 5300 9160 5310
rect 9260 5300 9270 5310
rect 9340 5300 9350 5310
rect 9520 5300 9530 5310
rect 9560 5300 9570 5310
rect 200 5290 210 5300
rect 240 5290 300 5300
rect 320 5290 590 5300
rect 2080 5290 2090 5300
rect 2150 5290 2180 5300
rect 2250 5290 2370 5300
rect 2490 5290 2520 5300
rect 2680 5290 2700 5300
rect 4690 5290 4710 5300
rect 4740 5290 4750 5300
rect 5080 5290 5100 5300
rect 5120 5290 5140 5300
rect 5220 5290 5230 5300
rect 5590 5290 5650 5300
rect 5660 5290 5700 5300
rect 5850 5290 5920 5300
rect 6160 5290 6180 5300
rect 6520 5290 6550 5300
rect 6590 5290 6640 5300
rect 6670 5290 6680 5300
rect 6780 5290 6800 5300
rect 7250 5290 7260 5300
rect 8120 5290 8140 5300
rect 8170 5290 8180 5300
rect 8310 5290 8320 5300
rect 8370 5290 8380 5300
rect 8430 5290 8440 5300
rect 8660 5290 8670 5300
rect 9120 5290 9130 5300
rect 9520 5290 9530 5300
rect 190 5280 200 5290
rect 220 5280 310 5290
rect 330 5280 600 5290
rect 2080 5280 2090 5290
rect 2150 5280 2190 5290
rect 2250 5280 2370 5290
rect 2480 5280 2530 5290
rect 2680 5280 2700 5290
rect 4660 5280 4670 5290
rect 4710 5280 4750 5290
rect 5070 5280 5080 5290
rect 5120 5280 5140 5290
rect 5220 5280 5230 5290
rect 5580 5280 5690 5290
rect 5850 5280 5920 5290
rect 6170 5280 6190 5290
rect 6460 5280 6500 5290
rect 6590 5280 6630 5290
rect 6670 5280 6730 5290
rect 6780 5280 6790 5290
rect 6910 5280 6920 5290
rect 7240 5280 7250 5290
rect 8040 5280 8050 5290
rect 8130 5280 8140 5290
rect 8260 5280 8270 5290
rect 8370 5280 8380 5290
rect 8410 5280 8420 5290
rect 9040 5280 9050 5290
rect 9270 5280 9280 5290
rect 9970 5280 9980 5290
rect 180 5270 190 5280
rect 200 5270 300 5280
rect 340 5270 610 5280
rect 2160 5270 2190 5280
rect 2250 5270 2370 5280
rect 2480 5270 2560 5280
rect 2680 5270 2700 5280
rect 4710 5270 4780 5280
rect 5160 5270 5170 5280
rect 5490 5270 5500 5280
rect 5570 5270 5630 5280
rect 5660 5270 5680 5280
rect 5860 5270 5910 5280
rect 6170 5270 6190 5280
rect 6430 5270 6470 5280
rect 6580 5270 6620 5280
rect 6660 5270 6680 5280
rect 6750 5270 6760 5280
rect 6780 5270 6800 5280
rect 6910 5270 6930 5280
rect 7230 5270 7260 5280
rect 8000 5270 8010 5280
rect 8130 5270 8140 5280
rect 8280 5270 8290 5280
rect 8450 5270 8460 5280
rect 9330 5270 9340 5280
rect 9350 5270 9360 5280
rect 9860 5270 9870 5280
rect 180 5260 320 5270
rect 350 5260 610 5270
rect 2160 5260 2180 5270
rect 2240 5260 2380 5270
rect 2470 5260 2570 5270
rect 2650 5260 2700 5270
rect 3520 5260 3530 5270
rect 4710 5260 4720 5270
rect 4740 5260 4760 5270
rect 5480 5260 5630 5270
rect 5840 5260 5880 5270
rect 6170 5260 6200 5270
rect 6430 5260 6470 5270
rect 6500 5260 6560 5270
rect 6570 5260 6590 5270
rect 6620 5260 6640 5270
rect 6780 5260 6800 5270
rect 6910 5260 6930 5270
rect 7260 5260 7270 5270
rect 8260 5260 8270 5270
rect 8950 5260 8960 5270
rect 9130 5260 9140 5270
rect 9360 5260 9370 5270
rect 9880 5260 9890 5270
rect 170 5250 340 5260
rect 370 5250 610 5260
rect 2170 5250 2180 5260
rect 2250 5250 2380 5260
rect 2470 5250 2590 5260
rect 2650 5250 2700 5260
rect 2750 5250 2790 5260
rect 4710 5250 4720 5260
rect 4740 5250 4760 5260
rect 5520 5250 5550 5260
rect 5600 5250 5630 5260
rect 5810 5250 5850 5260
rect 6180 5250 6210 5260
rect 6230 5250 6240 5260
rect 6450 5250 6530 5260
rect 6600 5250 6620 5260
rect 7230 5250 7240 5260
rect 7260 5250 7270 5260
rect 8050 5250 8060 5260
rect 8260 5250 8270 5260
rect 8280 5250 8290 5260
rect 9040 5250 9050 5260
rect 9100 5250 9110 5260
rect 9360 5250 9370 5260
rect 9390 5250 9400 5260
rect 9890 5250 9900 5260
rect 9950 5250 9960 5260
rect 9980 5250 9990 5260
rect 150 5240 370 5250
rect 380 5240 600 5250
rect 2160 5240 2180 5250
rect 2250 5240 2380 5250
rect 2470 5240 2610 5250
rect 2650 5240 2690 5250
rect 2740 5240 2790 5250
rect 4710 5240 4740 5250
rect 5060 5240 5070 5250
rect 5120 5240 5140 5250
rect 5220 5240 5230 5250
rect 5560 5240 5590 5250
rect 5780 5240 5820 5250
rect 6180 5240 6240 5250
rect 6250 5240 6270 5250
rect 6580 5240 6630 5250
rect 7260 5240 7270 5250
rect 8010 5240 8020 5250
rect 8340 5240 8350 5250
rect 8380 5240 8390 5250
rect 8490 5240 8500 5250
rect 9170 5240 9180 5250
rect 9390 5240 9400 5250
rect 9750 5240 9760 5250
rect 9980 5240 9990 5250
rect 140 5230 430 5240
rect 440 5230 620 5240
rect 2160 5230 2190 5240
rect 2250 5230 2380 5240
rect 2470 5230 2630 5240
rect 2660 5230 2690 5240
rect 2730 5230 2790 5240
rect 2840 5230 2870 5240
rect 4670 5230 4680 5240
rect 4720 5230 4740 5240
rect 5210 5230 5230 5240
rect 5600 5230 5620 5240
rect 5730 5230 5790 5240
rect 6180 5230 6300 5240
rect 6310 5230 6330 5240
rect 6600 5230 6610 5240
rect 7270 5230 7280 5240
rect 8100 5230 8110 5240
rect 8840 5230 8860 5240
rect 8980 5230 8990 5240
rect 9320 5230 9330 5240
rect 9960 5230 9970 5240
rect 120 5220 430 5230
rect 450 5220 620 5230
rect 2110 5220 2120 5230
rect 2160 5220 2190 5230
rect 2250 5220 2380 5230
rect 2470 5220 2650 5230
rect 2660 5220 2690 5230
rect 2730 5220 2790 5230
rect 2830 5220 2880 5230
rect 3500 5220 3510 5230
rect 4740 5220 4780 5230
rect 5210 5220 5230 5230
rect 5670 5220 5720 5230
rect 6180 5220 6340 5230
rect 6590 5220 6600 5230
rect 7270 5220 7290 5230
rect 7300 5220 7310 5230
rect 8220 5220 8230 5230
rect 8300 5220 8310 5230
rect 8410 5220 8420 5230
rect 8830 5220 8840 5230
rect 9050 5220 9060 5230
rect 9090 5220 9100 5230
rect 9140 5220 9150 5230
rect 9930 5220 9940 5230
rect 100 5210 620 5220
rect 2100 5210 2120 5220
rect 2180 5210 2210 5220
rect 2250 5210 2380 5220
rect 2460 5210 2570 5220
rect 2610 5210 2670 5220
rect 2730 5210 2800 5220
rect 2820 5210 2890 5220
rect 4770 5210 4780 5220
rect 5200 5210 5230 5220
rect 6180 5210 6270 5220
rect 6330 5210 6360 5220
rect 6560 5210 6580 5220
rect 7190 5210 7260 5220
rect 7290 5210 7330 5220
rect 8020 5210 8030 5220
rect 8220 5210 8230 5220
rect 8270 5210 8280 5220
rect 8310 5210 8320 5220
rect 8830 5210 8840 5220
rect 8990 5210 9000 5220
rect 9100 5210 9110 5220
rect 9710 5210 9720 5220
rect 9790 5210 9800 5220
rect 9860 5210 9870 5220
rect 9900 5210 9910 5220
rect 9940 5210 9950 5220
rect 9980 5210 9990 5220
rect 90 5200 620 5210
rect 650 5200 680 5210
rect 2090 5200 2120 5210
rect 2190 5200 2210 5210
rect 2250 5200 2380 5210
rect 2460 5200 2570 5210
rect 2620 5200 2650 5210
rect 2660 5200 2670 5210
rect 2730 5200 2790 5210
rect 2810 5200 2890 5210
rect 3490 5200 3500 5210
rect 5200 5200 5230 5210
rect 6190 5200 6270 5210
rect 6350 5200 6440 5210
rect 6460 5200 6510 5210
rect 6520 5200 6560 5210
rect 7140 5200 7160 5210
rect 7180 5200 7230 5210
rect 7280 5200 7290 5210
rect 7320 5200 7330 5210
rect 8180 5200 8190 5210
rect 8220 5200 8230 5210
rect 8340 5200 8350 5210
rect 8750 5200 8760 5210
rect 9090 5200 9100 5210
rect 9180 5200 9190 5210
rect 9330 5200 9340 5210
rect 9920 5200 9930 5210
rect 9950 5200 9980 5210
rect 70 5190 620 5200
rect 660 5190 680 5200
rect 2090 5190 2130 5200
rect 2250 5190 2390 5200
rect 2460 5190 2560 5200
rect 2660 5190 2670 5200
rect 2740 5190 2790 5200
rect 2810 5190 2890 5200
rect 5060 5190 5070 5200
rect 5190 5190 5230 5200
rect 6190 5190 6270 5200
rect 6360 5190 6400 5200
rect 7220 5190 7260 5200
rect 7280 5190 7290 5200
rect 8120 5190 8130 5200
rect 8180 5190 8190 5200
rect 8220 5190 8230 5200
rect 8700 5190 8710 5200
rect 8780 5190 8790 5200
rect 8840 5190 8850 5200
rect 9060 5190 9070 5200
rect 9090 5190 9100 5200
rect 9740 5190 9750 5200
rect 9830 5190 9840 5200
rect 9870 5190 9880 5200
rect 9890 5190 9900 5200
rect 60 5180 620 5190
rect 640 5180 660 5190
rect 2100 5180 2110 5190
rect 2120 5180 2130 5190
rect 2250 5180 2380 5190
rect 2460 5180 2510 5190
rect 2520 5180 2560 5190
rect 2670 5180 2680 5190
rect 2750 5180 2780 5190
rect 2810 5180 2880 5190
rect 3480 5180 3490 5190
rect 5200 5180 5220 5190
rect 6220 5180 6270 5190
rect 7260 5180 7290 5190
rect 8030 5180 8040 5190
rect 8090 5180 8100 5190
rect 8670 5180 8680 5190
rect 8720 5180 8730 5190
rect 8750 5180 8760 5190
rect 8780 5180 8790 5190
rect 8870 5180 8880 5190
rect 9010 5180 9020 5190
rect 9140 5180 9150 5190
rect 9530 5180 9540 5190
rect 9950 5180 9960 5190
rect 40 5170 620 5180
rect 660 5170 680 5180
rect 2100 5170 2110 5180
rect 2190 5170 2210 5180
rect 2250 5170 2390 5180
rect 2460 5170 2550 5180
rect 2680 5170 2690 5180
rect 2790 5170 2860 5180
rect 5200 5170 5220 5180
rect 6230 5170 6280 5180
rect 7280 5170 7290 5180
rect 8090 5170 8100 5180
rect 8130 5170 8140 5180
rect 8630 5170 8640 5180
rect 8720 5170 8730 5180
rect 8930 5170 8940 5180
rect 8960 5170 8970 5180
rect 8980 5170 8990 5180
rect 9510 5170 9520 5180
rect 9710 5170 9720 5180
rect 9810 5170 9820 5180
rect 9960 5170 9970 5180
rect 30 5160 130 5170
rect 140 5160 610 5170
rect 2180 5160 2230 5170
rect 2260 5160 2390 5170
rect 2420 5160 2430 5170
rect 2460 5160 2550 5170
rect 2670 5160 2700 5170
rect 2800 5160 2850 5170
rect 3470 5160 3480 5170
rect 5200 5160 5220 5170
rect 8090 5160 8100 5170
rect 8610 5160 8620 5170
rect 8700 5160 8710 5170
rect 8810 5160 8820 5170
rect 8930 5160 8940 5170
rect 8960 5160 8970 5170
rect 8980 5160 8990 5170
rect 9100 5160 9110 5170
rect 9560 5160 9570 5170
rect 9880 5160 9890 5170
rect 20 5150 130 5160
rect 140 5150 580 5160
rect 590 5150 610 5160
rect 2190 5150 2230 5160
rect 2260 5150 2400 5160
rect 2410 5150 2430 5160
rect 2460 5150 2530 5160
rect 2660 5150 2710 5160
rect 2800 5150 2810 5160
rect 2820 5150 2850 5160
rect 5200 5150 5230 5160
rect 7290 5150 7310 5160
rect 8040 5150 8050 5160
rect 8150 5150 8160 5160
rect 8760 5150 8770 5160
rect 8880 5150 8890 5160
rect 8930 5150 8940 5160
rect 9030 5150 9040 5160
rect 9100 5150 9110 5160
rect 9750 5150 9760 5160
rect 9910 5150 9920 5160
rect 0 5140 130 5150
rect 140 5140 570 5150
rect 2200 5140 2220 5150
rect 2260 5140 2430 5150
rect 2460 5140 2530 5150
rect 2650 5140 2680 5150
rect 2690 5140 2730 5150
rect 2820 5140 2850 5150
rect 3470 5140 3490 5150
rect 5090 5140 5100 5150
rect 5200 5140 5220 5150
rect 7300 5140 7310 5150
rect 8620 5140 8640 5150
rect 8760 5140 8770 5150
rect 8840 5140 8860 5150
rect 8880 5140 8890 5150
rect 8930 5140 8940 5150
rect 9080 5140 9100 5150
rect 9380 5140 9400 5150
rect 9590 5140 9600 5150
rect 9620 5140 9630 5150
rect 0 5130 130 5140
rect 140 5130 530 5140
rect 540 5130 570 5140
rect 2110 5130 2120 5140
rect 2200 5130 2220 5140
rect 2260 5130 2420 5140
rect 2460 5130 2540 5140
rect 2660 5130 2750 5140
rect 3450 5130 3460 5140
rect 3480 5130 3490 5140
rect 5210 5130 5220 5140
rect 7300 5130 7310 5140
rect 8050 5130 8060 5140
rect 8080 5130 8090 5140
rect 8480 5130 8490 5140
rect 8660 5130 8670 5140
rect 8930 5130 8940 5140
rect 8980 5130 8990 5140
rect 9510 5130 9520 5140
rect 0 5120 130 5130
rect 150 5120 520 5130
rect 560 5120 570 5130
rect 2110 5120 2130 5130
rect 2200 5120 2230 5130
rect 2260 5120 2420 5130
rect 2460 5120 2550 5130
rect 2660 5120 2750 5130
rect 3460 5120 3490 5130
rect 5110 5120 5120 5130
rect 5210 5120 5220 5130
rect 7300 5120 7310 5130
rect 8690 5120 8700 5130
rect 8960 5120 8970 5130
rect 9300 5120 9310 5130
rect 9410 5120 9420 5130
rect 9810 5120 9820 5130
rect 0 5110 130 5120
rect 150 5110 520 5120
rect 2130 5110 2140 5120
rect 2200 5110 2230 5120
rect 2260 5110 2410 5120
rect 2420 5110 2430 5120
rect 2470 5110 2560 5120
rect 2610 5110 2770 5120
rect 3450 5110 3460 5120
rect 5140 5110 5150 5120
rect 5210 5110 5220 5120
rect 7300 5110 7310 5120
rect 8770 5110 8780 5120
rect 9400 5110 9410 5120
rect 9600 5110 9610 5120
rect 9730 5110 9740 5120
rect 9800 5110 9810 5120
rect 0 5100 140 5110
rect 150 5100 520 5110
rect 2140 5100 2150 5110
rect 2200 5100 2230 5110
rect 2260 5100 2410 5110
rect 2460 5100 2580 5110
rect 2590 5100 2650 5110
rect 2660 5100 2730 5110
rect 2750 5100 2780 5110
rect 3430 5100 3440 5110
rect 3470 5100 3500 5110
rect 5140 5100 5150 5110
rect 5210 5100 5220 5110
rect 7290 5100 7300 5110
rect 8860 5100 8870 5110
rect 8890 5100 8900 5110
rect 9370 5100 9380 5110
rect 0 5090 140 5100
rect 160 5090 470 5100
rect 2140 5090 2150 5100
rect 2220 5090 2230 5100
rect 2270 5090 2410 5100
rect 2420 5090 2430 5100
rect 2470 5090 2720 5100
rect 2750 5090 2790 5100
rect 3450 5090 3470 5100
rect 5210 5090 5220 5100
rect 7290 5090 7300 5100
rect 8420 5090 8430 5100
rect 8670 5090 8680 5100
rect 8890 5090 8900 5100
rect 9430 5090 9440 5100
rect 9820 5090 9830 5100
rect 0 5080 140 5090
rect 160 5080 480 5090
rect 500 5080 520 5090
rect 2220 5080 2230 5090
rect 2270 5080 2430 5090
rect 2460 5080 2710 5090
rect 2720 5080 2790 5090
rect 3450 5080 3460 5090
rect 3500 5080 3510 5090
rect 5150 5080 5160 5090
rect 5210 5080 5220 5090
rect 7290 5080 7300 5090
rect 8380 5080 8390 5090
rect 8700 5080 8710 5090
rect 9150 5080 9160 5090
rect 9260 5080 9270 5090
rect 9550 5080 9560 5090
rect 0 5070 140 5080
rect 170 5070 450 5080
rect 480 5070 540 5080
rect 2280 5070 2430 5080
rect 2480 5070 2680 5080
rect 2710 5070 2790 5080
rect 3410 5070 3420 5080
rect 3510 5070 3520 5080
rect 5220 5070 5230 5080
rect 7240 5070 7250 5080
rect 7290 5070 7300 5080
rect 8490 5070 8500 5080
rect 8510 5070 8520 5080
rect 9110 5070 9120 5080
rect 9380 5070 9390 5080
rect 9460 5070 9470 5080
rect 0 5060 40 5070
rect 70 5060 150 5070
rect 170 5060 370 5070
rect 2230 5060 2240 5070
rect 2280 5060 2420 5070
rect 2500 5060 2670 5070
rect 2700 5060 2740 5070
rect 3400 5060 3420 5070
rect 3520 5060 3530 5070
rect 5220 5060 5230 5070
rect 6300 5060 6320 5070
rect 7290 5060 7300 5070
rect 8280 5060 8290 5070
rect 8350 5060 8360 5070
rect 8430 5060 8440 5070
rect 8790 5060 8810 5070
rect 9430 5060 9440 5070
rect 9530 5060 9540 5070
rect 9630 5060 9640 5070
rect 0 5050 30 5060
rect 50 5050 160 5060
rect 170 5050 310 5060
rect 320 5050 360 5060
rect 2230 5050 2240 5060
rect 2270 5050 2430 5060
rect 2520 5050 2650 5060
rect 2700 5050 2720 5060
rect 3400 5050 3410 5060
rect 5150 5050 5160 5060
rect 5220 5050 5230 5060
rect 6300 5050 6320 5060
rect 7300 5050 7320 5060
rect 8180 5050 8190 5060
rect 9040 5050 9050 5060
rect 9310 5050 9320 5060
rect 9570 5050 9580 5060
rect 0 5040 40 5050
rect 50 5040 300 5050
rect 320 5040 360 5050
rect 2270 5040 2430 5050
rect 2520 5040 2600 5050
rect 2630 5040 2640 5050
rect 5150 5040 5160 5050
rect 5220 5040 5230 5050
rect 5710 5040 5800 5050
rect 6310 5040 6330 5050
rect 7210 5040 7230 5050
rect 7290 5040 7300 5050
rect 7310 5040 7360 5050
rect 8680 5040 8690 5050
rect 9060 5040 9070 5050
rect 9170 5040 9180 5050
rect 9280 5040 9290 5050
rect 9390 5040 9400 5050
rect 0 5030 170 5040
rect 180 5030 340 5040
rect 2280 5030 2440 5040
rect 2520 5030 2650 5040
rect 3410 5030 3420 5040
rect 5150 5030 5160 5040
rect 5200 5030 5210 5040
rect 5680 5030 5800 5040
rect 6300 5030 6350 5040
rect 7210 5030 7230 5040
rect 7300 5030 7310 5040
rect 8360 5030 8370 5040
rect 8990 5030 9000 5040
rect 9540 5030 9550 5040
rect 9580 5030 9590 5040
rect 0 5020 170 5030
rect 200 5020 350 5030
rect 2280 5020 2440 5030
rect 2540 5020 2580 5030
rect 2620 5020 2650 5030
rect 3400 5020 3420 5030
rect 3510 5020 3520 5030
rect 5660 5020 5800 5030
rect 6310 5020 6370 5030
rect 7300 5020 7310 5030
rect 8090 5020 8110 5030
rect 8320 5020 8330 5030
rect 8340 5020 8350 5030
rect 8390 5020 8400 5030
rect 8440 5020 8450 5030
rect 9140 5020 9150 5030
rect 9450 5020 9460 5030
rect 0 5010 170 5020
rect 200 5010 380 5020
rect 2300 5010 2450 5020
rect 2500 5010 2510 5020
rect 2550 5010 2570 5020
rect 3400 5010 3410 5020
rect 3510 5010 3520 5020
rect 4160 5010 4170 5020
rect 5200 5010 5230 5020
rect 5630 5010 5740 5020
rect 5780 5010 5800 5020
rect 6310 5010 6390 5020
rect 6400 5010 6410 5020
rect 7210 5010 7230 5020
rect 7300 5010 7310 5020
rect 8080 5010 8090 5020
rect 8110 5010 8120 5020
rect 8260 5010 8270 5020
rect 8290 5010 8300 5020
rect 8380 5010 8390 5020
rect 8500 5010 8510 5020
rect 8540 5010 8550 5020
rect 8890 5010 8910 5020
rect 8960 5010 8970 5020
rect 9000 5010 9010 5020
rect 9320 5010 9330 5020
rect 0 5000 180 5010
rect 220 5000 370 5010
rect 2300 5000 2450 5010
rect 3510 5000 3520 5010
rect 4120 5000 4130 5010
rect 5160 5000 5170 5010
rect 5200 5000 5230 5010
rect 5620 5000 5710 5010
rect 5780 5000 5790 5010
rect 6320 5000 6330 5010
rect 6340 5000 6350 5010
rect 6360 5000 6420 5010
rect 7210 5000 7230 5010
rect 7300 5000 7310 5010
rect 8000 5000 8010 5010
rect 8180 5000 8190 5010
rect 8370 5000 8380 5010
rect 8880 5000 8890 5010
rect 8920 5000 8930 5010
rect 8960 5000 8970 5010
rect 9180 5000 9190 5010
rect 0 4990 200 5000
rect 230 4990 370 5000
rect 2310 4990 2440 5000
rect 2590 4990 2600 5000
rect 3400 4990 3410 5000
rect 3510 4990 3530 5000
rect 4020 4990 4030 5000
rect 4200 4990 4220 5000
rect 4270 4990 4300 5000
rect 5170 4990 5180 5000
rect 5190 4990 5230 5000
rect 5600 4990 5700 5000
rect 5780 4990 5790 5000
rect 6330 4990 6340 5000
rect 6370 4990 6470 5000
rect 7300 4990 7310 5000
rect 8040 4990 8050 5000
rect 8230 4990 8240 5000
rect 8380 4990 8390 5000
rect 8880 4990 8890 5000
rect 9040 4990 9050 5000
rect 9150 4990 9160 5000
rect 9300 4990 9310 5000
rect 9410 4990 9440 5000
rect 0 4980 210 4990
rect 240 4980 370 4990
rect 2310 4980 2450 4990
rect 3390 4980 3400 4990
rect 3510 4980 3520 4990
rect 4010 4980 4030 4990
rect 4220 4980 4230 4990
rect 4280 4980 4290 4990
rect 4330 4980 4340 4990
rect 4560 4980 4570 4990
rect 5220 4980 5230 4990
rect 5570 4980 5660 4990
rect 5670 4980 5690 4990
rect 5770 4980 5780 4990
rect 6330 4980 6340 4990
rect 6390 4980 6480 4990
rect 8070 4980 8080 4990
rect 8230 4980 8240 4990
rect 8330 4980 8340 4990
rect 8820 4980 8830 4990
rect 8880 4980 8890 4990
rect 9300 4980 9310 4990
rect 0 4970 220 4980
rect 260 4970 370 4980
rect 2320 4970 2460 4980
rect 3390 4970 3400 4980
rect 3510 4970 3520 4980
rect 4000 4970 4010 4980
rect 4080 4970 4090 4980
rect 4200 4970 4210 4980
rect 4280 4970 4290 4980
rect 4360 4970 4370 4980
rect 4390 4970 4410 4980
rect 4510 4970 4520 4980
rect 5510 4970 5640 4980
rect 5770 4970 5780 4980
rect 6120 4970 6150 4980
rect 6330 4970 6340 4980
rect 6400 4970 6500 4980
rect 7310 4970 7320 4980
rect 8000 4970 8010 4980
rect 8050 4970 8060 4980
rect 8070 4970 8080 4980
rect 8120 4970 8130 4980
rect 8150 4970 8160 4980
rect 9010 4970 9020 4980
rect 9670 4970 9680 4980
rect 0 4960 240 4970
rect 280 4960 380 4970
rect 2330 4960 2460 4970
rect 3500 4960 3520 4970
rect 4080 4960 4090 4970
rect 4190 4960 4200 4970
rect 4380 4960 4390 4970
rect 4400 4960 4420 4970
rect 4620 4960 4690 4970
rect 5230 4960 5240 4970
rect 5510 4960 5620 4970
rect 5770 4960 5790 4970
rect 5810 4960 5820 4970
rect 5830 4960 5880 4970
rect 5920 4960 5980 4970
rect 6040 4960 6200 4970
rect 6320 4960 6340 4970
rect 6410 4960 6540 4970
rect 7310 4960 7320 4970
rect 7860 4960 7870 4970
rect 7910 4960 7920 4970
rect 8000 4960 8010 4970
rect 8190 4960 8200 4970
rect 8270 4960 8280 4970
rect 8370 4960 8380 4970
rect 8740 4960 8750 4970
rect 9050 4960 9060 4970
rect 9160 4960 9170 4970
rect 0 4950 260 4960
rect 300 4950 390 4960
rect 2340 4950 2460 4960
rect 3380 4950 3390 4960
rect 3500 4950 3520 4960
rect 4000 4950 4010 4960
rect 4390 4950 4420 4960
rect 4450 4950 4490 4960
rect 4590 4950 4600 4960
rect 4610 4950 4620 4960
rect 4650 4950 4710 4960
rect 5190 4950 5200 4960
rect 5230 4950 5240 4960
rect 5500 4950 5610 4960
rect 5760 4950 5980 4960
rect 6010 4950 6230 4960
rect 6240 4950 6340 4960
rect 6430 4950 6610 4960
rect 8000 4950 8010 4960
rect 8190 4950 8200 4960
rect 8270 4950 8280 4960
rect 8390 4950 8400 4960
rect 8650 4950 8670 4960
rect 8770 4950 8780 4960
rect 8850 4950 8860 4960
rect 8890 4950 8900 4960
rect 9690 4950 9700 4960
rect 0 4940 180 4950
rect 190 4940 220 4950
rect 250 4940 260 4950
rect 2340 4940 2460 4950
rect 3510 4940 3520 4950
rect 4090 4940 4100 4950
rect 4180 4940 4190 4950
rect 4430 4940 4440 4950
rect 4480 4940 4490 4950
rect 4520 4940 4530 4950
rect 4640 4940 4660 4950
rect 4710 4940 4720 4950
rect 4740 4940 4750 4950
rect 4760 4940 4780 4950
rect 5190 4940 5200 4950
rect 5490 4940 5600 4950
rect 5750 4940 6140 4950
rect 6190 4940 6340 4950
rect 6440 4940 6580 4950
rect 6590 4940 6640 4950
rect 6670 4940 6680 4950
rect 7930 4940 7940 4950
rect 8230 4940 8240 4950
rect 8270 4940 8280 4950
rect 8310 4940 8320 4950
rect 8630 4940 8640 4950
rect 8740 4940 8750 4950
rect 8770 4940 8780 4950
rect 8980 4940 8990 4950
rect 9240 4940 9250 4950
rect 9550 4940 9560 4950
rect 0 4930 110 4940
rect 2340 4930 2470 4940
rect 3370 4930 3380 4940
rect 3510 4930 3520 4940
rect 3990 4930 4000 4940
rect 4180 4930 4190 4940
rect 4550 4930 4560 4940
rect 4710 4930 4740 4940
rect 4760 4930 4790 4940
rect 5190 4930 5210 4940
rect 5470 4930 5590 4940
rect 5740 4930 5790 4940
rect 5900 4930 5930 4940
rect 5940 4930 6140 4940
rect 6200 4930 6230 4940
rect 6300 4930 6330 4940
rect 6450 4930 6680 4940
rect 7230 4930 7240 4940
rect 7320 4930 7330 4940
rect 7870 4930 7880 4940
rect 8210 4930 8220 4940
rect 9260 4930 9270 4940
rect 9540 4930 9550 4940
rect 0 4920 80 4930
rect 2350 4920 2470 4930
rect 3370 4920 3380 4930
rect 3480 4920 3500 4930
rect 3510 4920 3520 4930
rect 4140 4920 4150 4930
rect 4170 4920 4190 4930
rect 4360 4920 4380 4930
rect 4480 4920 4490 4930
rect 4540 4920 4550 4930
rect 4600 4920 4610 4930
rect 4740 4920 4770 4930
rect 4810 4920 4820 4930
rect 5040 4920 5050 4930
rect 5060 4920 5090 4930
rect 5190 4920 5210 4930
rect 5450 4920 5580 4930
rect 5740 4920 5790 4930
rect 5930 4920 5960 4930
rect 5970 4920 6130 4930
rect 6450 4920 6690 4930
rect 7320 4920 7330 4930
rect 7760 4920 7770 4930
rect 7790 4920 7800 4930
rect 7860 4920 7870 4930
rect 7900 4920 7910 4930
rect 8130 4920 8140 4930
rect 8600 4920 8610 4930
rect 8660 4920 8670 4930
rect 8850 4920 8860 4930
rect 8900 4920 8910 4930
rect 8940 4920 8950 4930
rect 9020 4920 9030 4930
rect 9060 4920 9070 4930
rect 9090 4920 9100 4930
rect 0 4910 60 4920
rect 2370 4910 2480 4920
rect 2490 4910 2500 4920
rect 3360 4910 3380 4920
rect 3480 4910 3500 4920
rect 4000 4910 4010 4920
rect 4150 4910 4160 4920
rect 4170 4910 4180 4920
rect 4500 4910 4530 4920
rect 4570 4910 4580 4920
rect 4660 4910 4680 4920
rect 4790 4910 4830 4920
rect 5030 4910 5040 4920
rect 5060 4910 5080 4920
rect 5190 4910 5210 4920
rect 5240 4910 5250 4920
rect 5420 4910 5570 4920
rect 5740 4910 5790 4920
rect 5980 4910 6060 4920
rect 6080 4910 6090 4920
rect 6470 4910 6690 4920
rect 7760 4910 7770 4920
rect 7900 4910 7910 4920
rect 8010 4910 8020 4920
rect 8520 4910 8530 4920
rect 8540 4910 8550 4920
rect 8780 4910 8800 4920
rect 9090 4910 9100 4920
rect 9120 4910 9130 4920
rect 9480 4910 9490 4920
rect 9690 4910 9710 4920
rect 0 4900 40 4910
rect 2370 4900 2510 4910
rect 3340 4900 3350 4910
rect 3370 4900 3410 4910
rect 3470 4900 3480 4910
rect 3910 4900 3940 4910
rect 3950 4900 3970 4910
rect 4070 4900 4080 4910
rect 4160 4900 4180 4910
rect 4570 4900 4580 4910
rect 4600 4900 4620 4910
rect 4720 4900 4730 4910
rect 4830 4900 4840 4910
rect 4850 4900 4870 4910
rect 5050 4900 5070 4910
rect 5180 4900 5210 4910
rect 5240 4900 5250 4910
rect 5380 4900 5550 4910
rect 5730 4900 5790 4910
rect 6470 4900 6700 4910
rect 7230 4900 7240 4910
rect 7320 4900 7330 4910
rect 7720 4900 7730 4910
rect 7860 4900 7870 4910
rect 7940 4900 7950 4910
rect 8010 4900 8020 4910
rect 8060 4900 8070 4910
rect 8090 4900 8100 4910
rect 8200 4900 8220 4910
rect 8480 4900 8490 4910
rect 8560 4900 8570 4910
rect 8960 4900 8970 4910
rect 9080 4900 9090 4910
rect 9110 4900 9120 4910
rect 9450 4900 9460 4910
rect 9580 4900 9590 4910
rect 9620 4900 9630 4910
rect 0 4890 30 4900
rect 2380 4890 2520 4900
rect 2580 4890 2590 4900
rect 3330 4890 3350 4900
rect 3370 4890 3410 4900
rect 3460 4890 3480 4900
rect 3750 4890 3760 4900
rect 3860 4890 3870 4900
rect 3890 4890 3900 4900
rect 3940 4890 3960 4900
rect 4050 4890 4060 4900
rect 4170 4890 4190 4900
rect 4780 4890 4790 4900
rect 4820 4890 4830 4900
rect 4840 4890 4880 4900
rect 5030 4890 5060 4900
rect 5100 4890 5110 4900
rect 5180 4890 5210 4900
rect 5240 4890 5250 4900
rect 5380 4890 5540 4900
rect 5730 4890 5790 4900
rect 6480 4890 6700 4900
rect 7230 4890 7240 4900
rect 7320 4890 7330 4900
rect 7730 4890 7740 4900
rect 8070 4890 8090 4900
rect 8470 4890 8480 4900
rect 8570 4890 8580 4900
rect 8640 4890 8650 4900
rect 8670 4890 8680 4900
rect 8830 4890 8840 4900
rect 9100 4890 9110 4900
rect 9300 4890 9310 4900
rect 9410 4890 9420 4900
rect 0 4880 10 4890
rect 2370 4880 2520 4890
rect 3330 4880 3340 4890
rect 3370 4880 3430 4890
rect 3470 4880 3480 4890
rect 3710 4880 3730 4890
rect 3750 4880 3760 4890
rect 3840 4880 3850 4890
rect 3870 4880 3890 4890
rect 3910 4880 3920 4890
rect 3950 4880 3960 4890
rect 4030 4880 4040 4890
rect 4800 4880 4810 4890
rect 4830 4880 4870 4890
rect 4880 4880 4910 4890
rect 5180 4880 5210 4890
rect 5220 4880 5250 4890
rect 5380 4880 5520 4890
rect 5740 4880 5800 4890
rect 6500 4880 6710 4890
rect 7190 4880 7210 4890
rect 7230 4880 7240 4890
rect 7320 4880 7330 4890
rect 7740 4880 7750 4890
rect 7770 4880 7780 4890
rect 7800 4880 7810 4890
rect 8110 4880 8120 4890
rect 8130 4880 8140 4890
rect 8510 4880 8520 4890
rect 8540 4880 8550 4890
rect 8610 4880 8620 4890
rect 8700 4880 8710 4890
rect 8800 4880 8810 4890
rect 8840 4880 8850 4890
rect 8910 4880 8920 4890
rect 8940 4880 8950 4890
rect 9330 4880 9340 4890
rect 9530 4880 9540 4890
rect 9680 4880 9690 4890
rect 2370 4870 2530 4880
rect 2540 4870 2550 4880
rect 3350 4870 3360 4880
rect 3370 4870 3430 4880
rect 3740 4870 3750 4880
rect 3790 4870 3800 4880
rect 3910 4870 3920 4880
rect 3990 4870 4000 4880
rect 4840 4870 4850 4880
rect 4880 4870 4930 4880
rect 5180 4870 5210 4880
rect 5220 4870 5230 4880
rect 5240 4870 5250 4880
rect 5380 4870 5510 4880
rect 5750 4870 5800 4880
rect 6510 4870 6710 4880
rect 7210 4870 7220 4880
rect 7240 4870 7250 4880
rect 7750 4870 7760 4880
rect 7770 4870 7780 4880
rect 7830 4870 7840 4880
rect 7910 4870 7920 4880
rect 8020 4870 8030 4880
rect 8500 4870 8510 4880
rect 8810 4870 8820 4880
rect 8850 4870 8860 4880
rect 9090 4870 9100 4880
rect 9460 4870 9470 4880
rect 9530 4870 9540 4880
rect 9560 4870 9570 4880
rect 2370 4860 2570 4870
rect 2580 4860 2610 4870
rect 3350 4860 3370 4870
rect 3380 4860 3420 4870
rect 3730 4860 3790 4870
rect 3830 4860 3840 4870
rect 3980 4860 3990 4870
rect 4000 4860 4010 4870
rect 4870 4860 4880 4870
rect 4940 4860 4950 4870
rect 5180 4860 5240 4870
rect 5370 4860 5500 4870
rect 5750 4860 5810 4870
rect 6520 4860 6700 4870
rect 7760 4860 7770 4870
rect 7910 4860 7920 4870
rect 8470 4860 8480 4870
rect 9390 4860 9400 4870
rect 9420 4860 9430 4870
rect 9560 4860 9570 4870
rect 9590 4860 9600 4870
rect 9630 4860 9640 4870
rect 2380 4850 2610 4860
rect 3330 4850 3340 4860
rect 3360 4850 3370 4860
rect 3380 4850 3410 4860
rect 3670 4850 3680 4860
rect 3720 4850 3750 4860
rect 3770 4850 3820 4860
rect 3850 4850 3860 4860
rect 3980 4850 3990 4860
rect 4900 4850 4910 4860
rect 5190 4850 5240 4860
rect 5370 4850 5480 4860
rect 5740 4850 5830 4860
rect 6530 4850 6710 4860
rect 7870 4850 7880 4860
rect 8040 4850 8050 4860
rect 8300 4850 8310 4860
rect 8620 4850 8630 4860
rect 9420 4850 9430 4860
rect 9490 4850 9510 4860
rect 9550 4850 9560 4860
rect 2380 4840 2630 4850
rect 3360 4840 3370 4850
rect 3380 4840 3410 4850
rect 3720 4840 3730 4850
rect 3770 4840 3800 4850
rect 3850 4840 3860 4850
rect 3960 4840 3980 4850
rect 4940 4840 4950 4850
rect 5180 4840 5190 4850
rect 5200 4840 5240 4850
rect 5370 4840 5470 4850
rect 5740 4840 5840 4850
rect 6530 4840 6710 4850
rect 7330 4840 7340 4850
rect 7700 4840 7710 4850
rect 7730 4840 7750 4850
rect 7810 4840 7820 4850
rect 8280 4840 8290 4850
rect 8510 4840 8530 4850
rect 8570 4840 8580 4850
rect 9320 4840 9330 4850
rect 9670 4840 9680 4850
rect 9750 4840 9760 4850
rect 2390 4830 2630 4840
rect 3370 4830 3380 4840
rect 3390 4830 3400 4840
rect 3570 4830 3590 4840
rect 3960 4830 3970 4840
rect 4980 4830 4990 4840
rect 5180 4830 5190 4840
rect 5220 4830 5240 4840
rect 5370 4830 5460 4840
rect 5730 4830 5850 4840
rect 6530 4830 6720 4840
rect 7270 4830 7280 4840
rect 7750 4830 7760 4840
rect 7840 4830 7850 4840
rect 8210 4830 8220 4840
rect 8270 4830 8280 4840
rect 8650 4830 8660 4840
rect 8700 4830 8710 4840
rect 8770 4830 8780 4840
rect 9470 4830 9480 4840
rect 2390 4820 2650 4830
rect 2670 4820 2680 4830
rect 3370 4820 3380 4830
rect 3560 4820 3570 4830
rect 3580 4820 3590 4830
rect 3640 4820 3650 4830
rect 3940 4820 3960 4830
rect 5170 4820 5190 4830
rect 5370 4820 5450 4830
rect 5730 4820 5870 4830
rect 6550 4820 6720 4830
rect 7240 4820 7250 4830
rect 8480 4820 8490 4830
rect 8550 4820 8560 4830
rect 8660 4820 8670 4830
rect 9060 4820 9070 4830
rect 9400 4820 9410 4830
rect 9430 4820 9440 4830
rect 9570 4820 9580 4830
rect 9600 4820 9610 4830
rect 9640 4820 9650 4830
rect 2390 4810 2420 4820
rect 2430 4810 2670 4820
rect 3260 4810 3270 4820
rect 3380 4810 3390 4820
rect 3550 4810 3560 4820
rect 3570 4810 3580 4820
rect 3630 4810 3640 4820
rect 3920 4810 3940 4820
rect 5010 4810 5030 4820
rect 5360 4810 5460 4820
rect 5700 4810 5890 4820
rect 6580 4810 6720 4820
rect 7340 4810 7350 4820
rect 7770 4810 7780 4820
rect 7870 4810 7900 4820
rect 8300 4810 8310 4820
rect 9690 4810 9700 4820
rect 2390 4800 2430 4810
rect 2450 4800 2670 4810
rect 3250 4800 3260 4810
rect 3560 4800 3570 4810
rect 3620 4800 3630 4810
rect 5020 4800 5040 4810
rect 5170 4800 5180 4810
rect 5360 4800 5430 4810
rect 5700 4800 5910 4810
rect 5920 4800 5940 4810
rect 6580 4800 6730 4810
rect 7710 4800 7720 4810
rect 7740 4800 7750 4810
rect 8150 4800 8160 4810
rect 8700 4800 8710 4810
rect 9010 4800 9020 4810
rect 9050 4800 9060 4810
rect 2420 4790 2430 4800
rect 2440 4790 2680 4800
rect 3370 4790 3380 4800
rect 3540 4790 3550 4800
rect 3610 4790 3620 4800
rect 5030 4790 5050 4800
rect 5180 4790 5190 4800
rect 5350 4790 5420 4800
rect 5690 4790 5950 4800
rect 6580 4790 6720 4800
rect 7710 4790 7720 4800
rect 7800 4790 7810 4800
rect 8160 4790 8170 4800
rect 8200 4790 8210 4800
rect 8490 4790 8500 4800
rect 8520 4790 8530 4800
rect 8640 4790 8670 4800
rect 9480 4790 9490 4800
rect 9580 4790 9590 4800
rect 9600 4790 9610 4800
rect 2420 4780 2430 4790
rect 2440 4780 2690 4790
rect 3350 4780 3370 4790
rect 3550 4780 3560 4790
rect 3600 4780 3610 4790
rect 3880 4780 3890 4790
rect 5200 4780 5210 4790
rect 5340 4780 5410 4790
rect 5690 4780 5780 4790
rect 5840 4780 5960 4790
rect 6590 4780 6720 4790
rect 7340 4780 7350 4790
rect 7740 4780 7750 4790
rect 8020 4780 8030 4790
rect 8080 4780 8090 4790
rect 8170 4780 8180 4790
rect 8920 4780 8930 4790
rect 9030 4780 9050 4790
rect 9410 4780 9420 4790
rect 2450 4770 2690 4780
rect 3250 4770 3270 4780
rect 3350 4770 3360 4780
rect 5050 4770 5060 4780
rect 5230 4770 5240 4780
rect 5340 4770 5410 4780
rect 5670 4770 5780 4780
rect 5880 4770 5970 4780
rect 6620 4770 6630 4780
rect 6640 4770 6720 4780
rect 7340 4770 7350 4780
rect 8000 4770 8010 4780
rect 8090 4770 8100 4780
rect 8120 4770 8130 4780
rect 8180 4770 8190 4780
rect 8240 4770 8250 4780
rect 8290 4770 8300 4780
rect 8940 4770 8950 4780
rect 9300 4770 9310 4780
rect 2460 4760 2500 4770
rect 2510 4760 2720 4770
rect 3110 4760 3120 4770
rect 3250 4760 3260 4770
rect 3280 4760 3290 4770
rect 3350 4760 3360 4770
rect 3520 4760 3530 4770
rect 3540 4760 3560 4770
rect 3580 4760 3590 4770
rect 5080 4760 5090 4770
rect 5340 4760 5410 4770
rect 5670 4760 5760 4770
rect 5900 4760 5970 4770
rect 6640 4760 6720 4770
rect 8390 4760 8400 4770
rect 8910 4760 8920 4770
rect 8950 4760 8960 4770
rect 9310 4760 9320 4770
rect 9340 4760 9350 4770
rect 2480 4750 2490 4760
rect 2510 4750 2730 4760
rect 3250 4750 3260 4760
rect 3280 4750 3290 4760
rect 3350 4750 3370 4760
rect 3550 4750 3560 4760
rect 3570 4750 3580 4760
rect 3850 4750 3860 4760
rect 5090 4750 5100 4760
rect 5340 4750 5410 4760
rect 5660 4750 5760 4760
rect 5910 4750 5980 4760
rect 6640 4750 6730 4760
rect 7310 4750 7320 4760
rect 8040 4750 8070 4760
rect 8100 4750 8110 4760
rect 8200 4750 8220 4760
rect 8360 4750 8370 4760
rect 8390 4750 8400 4760
rect 8960 4750 8970 4760
rect 9440 4750 9450 4760
rect 2510 4740 2720 4750
rect 3280 4740 3290 4750
rect 3360 4740 3370 4750
rect 3510 4740 3520 4750
rect 3550 4740 3580 4750
rect 5100 4740 5110 4750
rect 5340 4740 5400 4750
rect 5650 4740 5750 4750
rect 5920 4740 5990 4750
rect 6640 4740 6720 4750
rect 6730 4740 6740 4750
rect 7300 4740 7310 4750
rect 8060 4740 8070 4750
rect 8100 4740 8110 4750
rect 8310 4740 8320 4750
rect 8920 4740 8930 4750
rect 9880 4740 9890 4750
rect 2550 4730 2710 4740
rect 3350 4730 3360 4740
rect 3540 4730 3560 4740
rect 5330 4730 5400 4740
rect 5640 4730 5740 4740
rect 5920 4730 6020 4740
rect 6310 4730 6320 4740
rect 6640 4730 6750 4740
rect 7360 4730 7370 4740
rect 7950 4730 7960 4740
rect 8020 4730 8030 4740
rect 8060 4730 8070 4740
rect 8130 4730 8140 4740
rect 8180 4730 8190 4740
rect 8250 4730 8260 4740
rect 8380 4730 8390 4740
rect 8830 4730 8840 4740
rect 8920 4730 8930 4740
rect 9010 4730 9020 4740
rect 9860 4730 9870 4740
rect 2550 4720 2710 4730
rect 3350 4720 3360 4730
rect 3500 4720 3510 4730
rect 3540 4720 3550 4730
rect 5130 4720 5140 4730
rect 5330 4720 5400 4730
rect 5640 4720 5740 4730
rect 5940 4720 6030 4730
rect 6240 4720 6250 4730
rect 6270 4720 6300 4730
rect 6640 4720 6760 4730
rect 7290 4720 7310 4730
rect 7360 4720 7370 4730
rect 9010 4720 9020 4730
rect 9330 4720 9340 4730
rect 2560 4710 2620 4720
rect 2650 4710 2710 4720
rect 3360 4710 3370 4720
rect 5100 4710 5110 4720
rect 5140 4710 5150 4720
rect 5200 4710 5210 4720
rect 5330 4710 5400 4720
rect 5650 4710 5770 4720
rect 5930 4710 6030 4720
rect 6070 4710 6080 4720
rect 6230 4710 6320 4720
rect 6640 4710 6760 4720
rect 7750 4710 7760 4720
rect 7800 4710 7810 4720
rect 7890 4710 7900 4720
rect 8070 4710 8080 4720
rect 8170 4710 8180 4720
rect 8650 4710 8660 4720
rect 8780 4710 8790 4720
rect 8890 4710 8900 4720
rect 9280 4710 9290 4720
rect 2580 4700 2640 4710
rect 3360 4700 3370 4710
rect 5150 4700 5160 4710
rect 5190 4700 5200 4710
rect 5220 4700 5230 4710
rect 5320 4700 5400 4710
rect 5650 4700 5780 4710
rect 5930 4700 6040 4710
rect 6050 4700 6100 4710
rect 6200 4700 6320 4710
rect 6650 4700 6750 4710
rect 7360 4700 7370 4710
rect 7730 4700 7740 4710
rect 7850 4700 7860 4710
rect 7990 4700 8000 4710
rect 8140 4700 8150 4710
rect 8610 4700 8630 4710
rect 8810 4700 8820 4710
rect 8860 4700 8870 4710
rect 9830 4700 9840 4710
rect 3360 4690 3370 4700
rect 3500 4690 3510 4700
rect 5110 4690 5120 4700
rect 5160 4690 5170 4700
rect 5310 4690 5390 4700
rect 5660 4690 5800 4700
rect 5820 4690 5830 4700
rect 5920 4690 6140 4700
rect 6180 4690 6320 4700
rect 6640 4690 6700 4700
rect 6710 4690 6760 4700
rect 7720 4690 7730 4700
rect 7890 4690 7900 4700
rect 7920 4690 7940 4700
rect 8110 4690 8120 4700
rect 8930 4690 8940 4700
rect 8960 4690 8970 4700
rect 3160 4680 3180 4690
rect 3370 4680 3390 4690
rect 3480 4680 3490 4690
rect 5170 4680 5180 4690
rect 5240 4680 5250 4690
rect 5310 4680 5390 4690
rect 5680 4680 6320 4690
rect 6640 4680 6700 4690
rect 6710 4680 6750 4690
rect 7370 4680 7380 4690
rect 7650 4680 7660 4690
rect 7720 4680 7730 4690
rect 7760 4680 7770 4690
rect 8110 4680 8120 4690
rect 8640 4680 8650 4690
rect 3280 4670 3290 4680
rect 3350 4670 3390 4680
rect 5300 4670 5390 4680
rect 5780 4670 6330 4680
rect 6640 4670 6750 4680
rect 7300 4670 7330 4680
rect 7380 4670 7390 4680
rect 7610 4670 7620 4680
rect 8030 4670 8040 4680
rect 8070 4670 8080 4680
rect 8110 4670 8120 4680
rect 8520 4670 8530 4680
rect 8820 4670 8830 4680
rect 8870 4670 8880 4680
rect 8900 4670 8910 4680
rect 3140 4660 3150 4670
rect 3160 4660 3170 4670
rect 3270 4660 3280 4670
rect 3350 4660 3380 4670
rect 3400 4660 3410 4670
rect 5130 4660 5140 4670
rect 5220 4660 5230 4670
rect 5300 4660 5390 4670
rect 5790 4660 5940 4670
rect 5990 4660 6080 4670
rect 6190 4660 6230 4670
rect 6250 4660 6300 4670
rect 6640 4660 6690 4670
rect 6700 4660 6750 4670
rect 7310 4660 7320 4670
rect 7380 4660 7390 4670
rect 7600 4660 7610 4670
rect 7760 4660 7770 4670
rect 7880 4660 7890 4670
rect 7970 4660 7980 4670
rect 8040 4660 8060 4670
rect 8110 4660 8120 4670
rect 8500 4660 8510 4670
rect 8790 4660 8800 4670
rect 8900 4660 8910 4670
rect 8990 4660 9000 4670
rect 9260 4660 9270 4670
rect 3150 4650 3160 4660
rect 3340 4650 3370 4660
rect 3400 4650 3420 4660
rect 3470 4650 3480 4660
rect 5150 4650 5160 4660
rect 5190 4650 5200 4660
rect 5300 4650 5390 4660
rect 6260 4650 6300 4660
rect 6640 4650 6690 4660
rect 6700 4650 6750 4660
rect 7240 4650 7260 4660
rect 7650 4650 7660 4660
rect 7780 4650 7790 4660
rect 8970 4650 8980 4660
rect 3340 4640 3370 4650
rect 3390 4640 3410 4650
rect 3460 4640 3470 4650
rect 5200 4640 5210 4650
rect 5300 4640 5400 4650
rect 6630 4640 6650 4650
rect 6660 4640 6750 4650
rect 7600 4640 7610 4650
rect 7730 4640 7740 4650
rect 7940 4640 7950 4650
rect 8610 4640 8620 4650
rect 9250 4640 9260 4650
rect 3360 4630 3410 4640
rect 5290 4630 5400 4640
rect 6630 4630 6750 4640
rect 7930 4630 7940 4640
rect 7970 4630 7980 4640
rect 8030 4630 8070 4640
rect 8320 4630 8330 4640
rect 8340 4630 8350 4640
rect 8950 4630 8960 4640
rect 8970 4630 8990 4640
rect 3350 4620 3370 4630
rect 3390 4620 3410 4630
rect 3420 4620 3460 4630
rect 5210 4620 5220 4630
rect 5280 4620 5380 4630
rect 6620 4620 6750 4630
rect 7530 4620 7540 4630
rect 7580 4620 7590 4630
rect 7640 4620 7650 4630
rect 7690 4620 7700 4630
rect 3300 4610 3310 4620
rect 3340 4610 3350 4620
rect 3400 4610 3430 4620
rect 5210 4610 5220 4620
rect 5280 4610 5380 4620
rect 6590 4610 6600 4620
rect 6610 4610 6740 4620
rect 7380 4610 7390 4620
rect 7510 4610 7520 4620
rect 7580 4610 7590 4620
rect 7690 4610 7700 4620
rect 7770 4610 7780 4620
rect 7820 4610 7830 4620
rect 8560 4610 8570 4620
rect 9240 4610 9250 4620
rect 3290 4600 3300 4610
rect 3390 4600 3420 4610
rect 5280 4600 5390 4610
rect 5800 4600 5820 4610
rect 6580 4600 6740 4610
rect 7310 4600 7330 4610
rect 7580 4600 7590 4610
rect 7680 4600 7690 4610
rect 7740 4600 7750 4610
rect 7770 4600 7790 4610
rect 7830 4600 7840 4610
rect 7940 4600 7950 4610
rect 8320 4600 8330 4610
rect 8340 4600 8350 4610
rect 8380 4600 8390 4610
rect 8530 4600 8540 4610
rect 8620 4600 8630 4610
rect 8650 4600 8660 4610
rect 8840 4600 8860 4610
rect 8970 4600 8980 4610
rect 3290 4590 3300 4600
rect 3340 4590 3350 4600
rect 5230 4590 5240 4600
rect 5280 4590 5390 4600
rect 5790 4590 5830 4600
rect 5870 4590 5890 4600
rect 5910 4590 6010 4600
rect 6580 4590 6740 4600
rect 7320 4590 7340 4600
rect 7380 4590 7390 4600
rect 7480 4590 7490 4600
rect 7540 4590 7550 4600
rect 7650 4590 7660 4600
rect 7740 4590 7750 4600
rect 8310 4590 8320 4600
rect 8350 4590 8360 4600
rect 8490 4590 8500 4600
rect 3330 4580 3340 4590
rect 3370 4580 3380 4590
rect 5280 4580 5390 4590
rect 5790 4580 5810 4590
rect 5820 4580 5840 4590
rect 5860 4580 5960 4590
rect 5980 4580 6030 4590
rect 6070 4580 6080 4590
rect 6100 4580 6110 4590
rect 6580 4580 6740 4590
rect 7320 4580 7330 4590
rect 7340 4580 7350 4590
rect 7520 4580 7530 4590
rect 8240 4580 8250 4590
rect 8350 4580 8360 4590
rect 8490 4580 8500 4590
rect 8520 4580 8530 4590
rect 9990 4580 9990 4590
rect 3330 4570 3340 4580
rect 3440 4570 3450 4580
rect 5280 4570 5290 4580
rect 5300 4570 5410 4580
rect 5430 4570 5450 4580
rect 5610 4570 5630 4580
rect 5790 4570 5800 4580
rect 5810 4570 6130 4580
rect 6570 4570 6740 4580
rect 7320 4570 7330 4580
rect 7380 4570 7390 4580
rect 8100 4570 8110 4580
rect 8210 4570 8220 4580
rect 8490 4570 8500 4580
rect 8520 4570 8550 4580
rect 8960 4570 8970 4580
rect 9980 4570 9990 4580
rect 3140 4560 3150 4570
rect 3260 4560 3270 4570
rect 3350 4560 3360 4570
rect 5240 4560 5250 4570
rect 5300 4560 5410 4570
rect 5430 4560 5460 4570
rect 5610 4560 5640 4570
rect 5650 4560 5660 4570
rect 5830 4560 5870 4570
rect 5900 4560 5950 4570
rect 6000 4560 6140 4570
rect 6560 4560 6730 4570
rect 7320 4560 7360 4570
rect 7670 4560 7680 4570
rect 7770 4560 7780 4570
rect 8320 4560 8340 4570
rect 8630 4560 8640 4570
rect 9230 4560 9240 4570
rect 9980 4560 9990 4570
rect 3250 4550 3260 4560
rect 3270 4550 3280 4560
rect 3320 4550 3330 4560
rect 5290 4550 5470 4560
rect 5610 4550 5670 4560
rect 5800 4550 5810 4560
rect 5830 4550 5870 4560
rect 5910 4550 5930 4560
rect 6010 4550 6090 4560
rect 6110 4550 6130 4560
rect 6240 4550 6270 4560
rect 6550 4550 6730 4560
rect 7320 4550 7330 4560
rect 7370 4550 7380 4560
rect 7490 4550 7500 4560
rect 7530 4550 7540 4560
rect 8020 4550 8030 4560
rect 8190 4550 8200 4560
rect 8650 4550 8660 4560
rect 9690 4550 9700 4560
rect 9980 4550 9990 4560
rect 3260 4540 3280 4550
rect 3320 4540 3340 4550
rect 3420 4540 3430 4550
rect 5250 4540 5260 4550
rect 5290 4540 5300 4550
rect 5310 4540 5460 4550
rect 5610 4540 5670 4550
rect 5800 4540 5810 4550
rect 5840 4540 5870 4550
rect 6020 4540 6060 4550
rect 6120 4540 6140 4550
rect 6160 4540 6200 4550
rect 6230 4540 6270 4550
rect 6550 4540 6720 4550
rect 7330 4540 7360 4550
rect 7370 4540 7380 4550
rect 7490 4540 7500 4550
rect 7620 4540 7630 4550
rect 7700 4540 7710 4550
rect 8060 4540 8070 4550
rect 8130 4540 8140 4550
rect 8220 4540 8230 4550
rect 8240 4540 8250 4550
rect 8290 4540 8300 4550
rect 8530 4540 8540 4550
rect 8570 4540 8580 4550
rect 9960 4540 9990 4550
rect 3250 4530 3270 4540
rect 3310 4530 3320 4540
rect 3340 4530 3350 4540
rect 3420 4530 3430 4540
rect 5290 4530 5300 4540
rect 5320 4530 5400 4540
rect 5410 4530 5450 4540
rect 5620 4530 5680 4540
rect 5810 4530 5820 4540
rect 5840 4530 5870 4540
rect 6020 4530 6040 4540
rect 6130 4530 6140 4540
rect 6150 4530 6160 4540
rect 6170 4530 6200 4540
rect 6230 4530 6260 4540
rect 6540 4530 6720 4540
rect 7330 4530 7340 4540
rect 7380 4530 7390 4540
rect 7670 4530 7680 4540
rect 7920 4530 7930 4540
rect 7960 4530 7970 4540
rect 8040 4530 8050 4540
rect 8090 4530 8100 4540
rect 8130 4530 8140 4540
rect 8160 4530 8170 4540
rect 8290 4530 8300 4540
rect 8370 4530 8380 4540
rect 9950 4530 9990 4540
rect 3250 4520 3270 4530
rect 3300 4520 3330 4530
rect 5290 4520 5300 4530
rect 5320 4520 5460 4530
rect 5620 4520 5690 4530
rect 5810 4520 5830 4530
rect 5850 4520 5870 4530
rect 6130 4520 6150 4530
rect 6180 4520 6260 4530
rect 6540 4520 6720 4530
rect 7350 4520 7360 4530
rect 7390 4520 7400 4530
rect 7530 4520 7540 4530
rect 8010 4520 8020 4530
rect 8130 4520 8140 4530
rect 8940 4520 8950 4530
rect 9940 4520 9980 4530
rect 3000 4510 3010 4520
rect 3240 4510 3260 4520
rect 3300 4510 3330 4520
rect 5270 4510 5280 4520
rect 5340 4510 5460 4520
rect 5610 4510 5690 4520
rect 5820 4510 5830 4520
rect 5840 4510 5850 4520
rect 6190 4510 6250 4520
rect 6530 4510 6710 4520
rect 7330 4510 7360 4520
rect 7890 4510 7900 4520
rect 8050 4510 8060 4520
rect 8330 4510 8340 4520
rect 9940 4510 9970 4520
rect 3250 4500 3260 4510
rect 3300 4500 3310 4510
rect 5300 4500 5310 4510
rect 5350 4500 5470 4510
rect 5610 4500 5700 4510
rect 6170 4500 6250 4510
rect 6530 4500 6710 4510
rect 7360 4500 7380 4510
rect 7400 4500 7410 4510
rect 7500 4500 7510 4510
rect 7810 4500 7820 4510
rect 7850 4500 7860 4510
rect 7940 4500 7950 4510
rect 8200 4500 8210 4510
rect 8330 4500 8340 4510
rect 9930 4500 9960 4510
rect 3260 4490 3270 4500
rect 5360 4490 5390 4500
rect 5420 4490 5480 4500
rect 5600 4490 5710 4500
rect 5820 4490 5830 4500
rect 5870 4490 5880 4500
rect 6170 4490 6240 4500
rect 6530 4490 6710 4500
rect 7330 4490 7340 4500
rect 7360 4490 7370 4500
rect 7770 4490 7780 4500
rect 7920 4490 7930 4500
rect 7990 4490 8000 4500
rect 8020 4490 8030 4500
rect 8170 4490 8180 4500
rect 9930 4490 9950 4500
rect 3000 4480 3030 4490
rect 3270 4480 3280 4490
rect 5360 4480 5400 4490
rect 5420 4480 5490 4490
rect 5590 4480 5720 4490
rect 5810 4480 5840 4490
rect 5860 4480 5900 4490
rect 6160 4480 6190 4490
rect 6210 4480 6230 4490
rect 6530 4480 6710 4490
rect 7360 4480 7370 4490
rect 7850 4480 7860 4490
rect 7880 4480 7890 4490
rect 8250 4480 8270 4490
rect 8300 4480 8310 4490
rect 9910 4480 9940 4490
rect 3080 4470 3090 4480
rect 5310 4470 5320 4480
rect 5350 4470 5400 4480
rect 5430 4470 5500 4480
rect 5590 4470 5730 4480
rect 5800 4470 5840 4480
rect 5860 4470 5890 4480
rect 6140 4470 6180 4480
rect 6210 4470 6220 4480
rect 6530 4470 6710 4480
rect 7360 4470 7370 4480
rect 8080 4470 8090 4480
rect 9210 4470 9220 4480
rect 9890 4470 9930 4480
rect 3000 4460 3010 4470
rect 3080 4460 3090 4470
rect 5290 4460 5310 4470
rect 5350 4460 5410 4470
rect 5430 4460 5500 4470
rect 5590 4460 5740 4470
rect 5790 4460 5830 4470
rect 5850 4460 5890 4470
rect 5920 4460 5930 4470
rect 6130 4460 6180 4470
rect 6520 4460 6710 4470
rect 7340 4460 7360 4470
rect 7410 4460 7420 4470
rect 7770 4460 7800 4470
rect 7960 4460 7970 4470
rect 8080 4460 8090 4470
rect 9880 4460 9920 4470
rect 3020 4450 3040 4460
rect 3290 4450 3300 4460
rect 5290 4450 5300 4460
rect 5320 4450 5330 4460
rect 5360 4450 5420 4460
rect 5430 4450 5500 4460
rect 5600 4450 5750 4460
rect 5790 4450 5830 4460
rect 5850 4450 5890 4460
rect 5930 4450 5960 4460
rect 6120 4450 6140 4460
rect 6530 4450 6710 4460
rect 7340 4450 7350 4460
rect 7830 4450 7840 4460
rect 7920 4450 7930 4460
rect 8000 4450 8010 4460
rect 8080 4450 8090 4460
rect 8180 4450 8190 4460
rect 8260 4450 8270 4460
rect 9870 4450 9910 4460
rect 2840 4440 2850 4450
rect 3000 4440 3030 4450
rect 3170 4440 3180 4450
rect 3290 4440 3300 4450
rect 5300 4440 5320 4450
rect 5330 4440 5340 4450
rect 5370 4440 5420 4450
rect 5430 4440 5500 4450
rect 5600 4440 5760 4450
rect 5790 4440 5820 4450
rect 5850 4440 5900 4450
rect 5920 4440 5940 4450
rect 5980 4440 6010 4450
rect 6030 4440 6070 4450
rect 6100 4440 6120 4450
rect 6520 4440 6700 4450
rect 7920 4440 7930 4450
rect 8080 4440 8090 4450
rect 8100 4440 8110 4450
rect 8140 4440 8150 4450
rect 8210 4440 8220 4450
rect 9870 4440 9890 4450
rect 2820 4430 2830 4440
rect 2840 4430 2850 4440
rect 3040 4430 3050 4440
rect 3180 4430 3190 4440
rect 5370 4430 5410 4440
rect 5430 4430 5510 4440
rect 5600 4430 5780 4440
rect 5800 4430 5820 4440
rect 5840 4430 5940 4440
rect 6180 4430 6190 4440
rect 6530 4430 6690 4440
rect 7340 4430 7370 4440
rect 7800 4430 7810 4440
rect 7890 4430 7900 4440
rect 8040 4430 8050 4440
rect 8860 4430 8870 4440
rect 9840 4430 9880 4440
rect 2990 4420 3020 4430
rect 3270 4420 3280 4430
rect 3370 4420 3380 4430
rect 5320 4420 5330 4430
rect 5340 4420 5350 4430
rect 5380 4420 5410 4430
rect 5440 4420 5510 4430
rect 5600 4420 5790 4430
rect 5840 4420 5960 4430
rect 5970 4420 6010 4430
rect 6170 4420 6200 4430
rect 6520 4420 6680 4430
rect 7240 4420 7250 4430
rect 7270 4420 7280 4430
rect 7340 4420 7350 4430
rect 7370 4420 7380 4430
rect 7410 4420 7420 4430
rect 9830 4420 9860 4430
rect 2980 4410 2990 4420
rect 3240 4410 3270 4420
rect 5310 4410 5320 4420
rect 5380 4410 5410 4420
rect 5450 4410 5520 4420
rect 5590 4410 5810 4420
rect 5860 4410 6010 4420
rect 6060 4410 6070 4420
rect 6110 4410 6130 4420
rect 6520 4410 6680 4420
rect 7240 4410 7250 4420
rect 7260 4410 7300 4420
rect 7340 4410 7370 4420
rect 7960 4410 7970 4420
rect 8000 4410 8010 4420
rect 8890 4410 8900 4420
rect 9840 4410 9850 4420
rect 2970 4400 3000 4410
rect 3010 4400 3020 4410
rect 3260 4400 3290 4410
rect 3360 4400 3370 4410
rect 5390 4400 5400 4410
rect 5460 4400 5520 4410
rect 5570 4400 5810 4410
rect 5820 4400 5840 4410
rect 5910 4400 5950 4410
rect 5970 4400 6020 4410
rect 6050 4400 6070 4410
rect 6100 4400 6140 4410
rect 6520 4400 6680 4410
rect 7240 4400 7250 4410
rect 7290 4400 7300 4410
rect 7340 4400 7370 4410
rect 7900 4400 7910 4410
rect 8850 4400 8860 4410
rect 9840 4400 9860 4410
rect 2810 4390 2820 4400
rect 2840 4390 2850 4400
rect 2970 4390 3010 4400
rect 3270 4390 3280 4400
rect 4650 4390 4680 4400
rect 5360 4390 5370 4400
rect 5390 4390 5440 4400
rect 5460 4390 5520 4400
rect 5570 4390 5800 4400
rect 5840 4390 5860 4400
rect 5970 4390 6010 4400
rect 6040 4390 6080 4400
rect 6110 4390 6130 4400
rect 6510 4390 6680 4400
rect 7240 4390 7250 4400
rect 7270 4390 7280 4400
rect 7340 4390 7370 4400
rect 7420 4390 7430 4400
rect 8850 4390 8860 4400
rect 8880 4390 8890 4400
rect 9190 4390 9200 4400
rect 9530 4390 9540 4400
rect 9850 4390 9860 4400
rect 2970 4380 3010 4390
rect 3040 4380 3050 4390
rect 3060 4380 3070 4390
rect 3240 4380 3250 4390
rect 3260 4380 3280 4390
rect 4630 4380 4700 4390
rect 5330 4380 5340 4390
rect 5400 4380 5420 4390
rect 5460 4380 5520 4390
rect 5570 4380 5800 4390
rect 5880 4380 5890 4390
rect 5980 4380 6000 4390
rect 6050 4380 6070 4390
rect 6500 4380 6680 4390
rect 7240 4380 7250 4390
rect 7270 4380 7280 4390
rect 7300 4380 7310 4390
rect 7330 4380 7370 4390
rect 7420 4380 7430 4390
rect 7810 4380 7820 4390
rect 7970 4380 7980 4390
rect 9520 4380 9530 4390
rect 9850 4380 9860 4390
rect 2860 4370 2870 4380
rect 2980 4370 3010 4380
rect 3070 4370 3080 4380
rect 3240 4370 3260 4380
rect 3270 4370 3280 4380
rect 4610 4370 4720 4380
rect 5340 4370 5350 4380
rect 5370 4370 5380 4380
rect 5410 4370 5430 4380
rect 5470 4370 5520 4380
rect 5560 4370 5800 4380
rect 5900 4370 5930 4380
rect 6500 4370 6680 4380
rect 7250 4370 7290 4380
rect 7340 4370 7370 4380
rect 8690 4370 8710 4380
rect 9840 4370 9850 4380
rect 2820 4360 2830 4370
rect 2960 4360 2970 4370
rect 2980 4360 3000 4370
rect 3060 4360 3070 4370
rect 3240 4360 3260 4370
rect 3270 4360 3290 4370
rect 4610 4360 4750 4370
rect 5340 4360 5350 4370
rect 5410 4360 5420 4370
rect 5470 4360 5540 4370
rect 5560 4360 5810 4370
rect 5940 4360 5950 4370
rect 6500 4360 6670 4370
rect 7250 4360 7260 4370
rect 7270 4360 7280 4370
rect 7330 4360 7360 4370
rect 7370 4360 7380 4370
rect 7410 4360 7420 4370
rect 8650 4360 8660 4370
rect 9180 4360 9190 4370
rect 9830 4360 9850 4370
rect 9990 4360 9990 4370
rect 2960 4350 2970 4360
rect 2980 4350 3000 4360
rect 3030 4350 3060 4360
rect 3280 4350 3300 4360
rect 4600 4350 4780 4360
rect 4800 4350 4810 4360
rect 5340 4350 5350 4360
rect 5470 4350 5820 4360
rect 5950 4350 6000 4360
rect 6490 4350 6670 4360
rect 7380 4350 7420 4360
rect 7840 4350 7850 4360
rect 8860 4350 8870 4360
rect 9820 4350 9840 4360
rect 2930 4340 2940 4350
rect 2970 4340 2980 4350
rect 2990 4340 3000 4350
rect 3020 4340 3040 4350
rect 3260 4340 3270 4350
rect 4590 4340 4830 4350
rect 5390 4340 5400 4350
rect 5430 4340 5450 4350
rect 5470 4340 5860 4350
rect 5950 4340 6060 4350
rect 6480 4340 6670 4350
rect 7240 4340 7260 4350
rect 7280 4340 7290 4350
rect 7380 4340 7420 4350
rect 8490 4340 8510 4350
rect 8610 4340 8620 4350
rect 9800 4340 9830 4350
rect 9950 4340 9960 4350
rect 9980 4340 9990 4350
rect 2930 4330 2940 4340
rect 2980 4330 3000 4340
rect 3020 4330 3030 4340
rect 3260 4330 3270 4340
rect 4590 4330 4840 4340
rect 5400 4330 5410 4340
rect 5480 4330 5880 4340
rect 5940 4330 6190 4340
rect 6200 4330 6220 4340
rect 6480 4330 6670 4340
rect 7350 4330 7360 4340
rect 8440 4330 8450 4340
rect 8550 4330 8560 4340
rect 8660 4330 8670 4340
rect 9800 4330 9820 4340
rect 9890 4330 9900 4340
rect 9960 4330 9980 4340
rect 2920 4320 2960 4330
rect 2970 4320 3010 4330
rect 3160 4320 3170 4330
rect 3280 4320 3300 4330
rect 4590 4320 4860 4330
rect 5490 4320 5900 4330
rect 5910 4320 6180 4330
rect 6470 4320 6580 4330
rect 6590 4320 6660 4330
rect 7340 4320 7350 4330
rect 8460 4320 8470 4330
rect 8560 4320 8570 4330
rect 9790 4320 9820 4330
rect 9840 4320 9860 4330
rect 9940 4320 9970 4330
rect 2920 4310 3000 4320
rect 3170 4310 3180 4320
rect 3280 4310 3300 4320
rect 4580 4310 4680 4320
rect 4780 4310 4880 4320
rect 5350 4310 5360 4320
rect 5410 4310 5420 4320
rect 5500 4310 5940 4320
rect 5950 4310 5970 4320
rect 5980 4310 5990 4320
rect 6010 4310 6140 4320
rect 6460 4310 6570 4320
rect 6590 4310 6660 4320
rect 7190 4310 7200 4320
rect 7310 4310 7320 4320
rect 8490 4310 8500 4320
rect 8570 4310 8580 4320
rect 9780 4310 9810 4320
rect 9890 4310 9900 4320
rect 9970 4310 9980 4320
rect 2950 4300 2960 4310
rect 3160 4300 3170 4310
rect 3220 4300 3230 4310
rect 4570 4300 4650 4310
rect 4810 4300 4890 4310
rect 5500 4300 5920 4310
rect 6450 4300 6550 4310
rect 6580 4300 6660 4310
rect 7250 4300 7260 4310
rect 8710 4300 8720 4310
rect 8860 4300 8870 4310
rect 9770 4300 9800 4310
rect 9880 4300 9900 4310
rect 9910 4300 9930 4310
rect 2920 4290 2940 4300
rect 2950 4290 2970 4300
rect 3170 4290 3180 4300
rect 3210 4290 3220 4300
rect 4570 4290 4650 4300
rect 4820 4290 4890 4300
rect 5510 4290 5930 4300
rect 6450 4290 6550 4300
rect 6580 4290 6650 4300
rect 7200 4290 7220 4300
rect 8440 4290 8450 4300
rect 8580 4290 8590 4300
rect 9760 4290 9800 4300
rect 9880 4290 9900 4300
rect 9910 4290 9920 4300
rect 9950 4290 9960 4300
rect 2920 4280 2940 4290
rect 2960 4280 2980 4290
rect 3060 4280 3080 4290
rect 3290 4280 3300 4290
rect 4570 4280 4610 4290
rect 4620 4280 4630 4290
rect 4820 4280 4910 4290
rect 5430 4280 5440 4290
rect 5510 4280 5940 4290
rect 6440 4280 6540 4290
rect 6570 4280 6650 4290
rect 8680 4280 8710 4290
rect 9750 4280 9770 4290
rect 9790 4280 9800 4290
rect 9830 4280 9840 4290
rect 9860 4280 9870 4290
rect 9880 4280 9900 4290
rect 9910 4280 9920 4290
rect 2960 4270 2970 4280
rect 3040 4270 3090 4280
rect 3230 4270 3240 4280
rect 4210 4270 4230 4280
rect 4560 4270 4610 4280
rect 4820 4270 4910 4280
rect 5390 4270 5410 4280
rect 5510 4270 5950 4280
rect 6430 4270 6540 4280
rect 6570 4270 6650 4280
rect 8850 4270 8860 4280
rect 9740 4270 9760 4280
rect 9830 4270 9850 4280
rect 9880 4270 9890 4280
rect 2820 4260 2830 4270
rect 2950 4260 2960 4270
rect 3040 4260 3050 4270
rect 3060 4260 3090 4270
rect 4200 4260 4290 4270
rect 4560 4260 4610 4270
rect 4840 4260 4910 4270
rect 5390 4260 5410 4270
rect 5430 4260 5450 4270
rect 5520 4260 5650 4270
rect 5660 4260 5950 4270
rect 6380 4260 6400 4270
rect 6420 4260 6530 4270
rect 6560 4260 6650 4270
rect 7050 4260 7070 4270
rect 7080 4260 7090 4270
rect 8470 4260 8480 4270
rect 9740 4260 9760 4270
rect 9820 4260 9860 4270
rect 9880 4260 9890 4270
rect 2940 4250 2950 4260
rect 3140 4250 3150 4260
rect 3170 4250 3180 4260
rect 4200 4250 4300 4260
rect 4550 4250 4610 4260
rect 4840 4250 4910 4260
rect 5520 4250 5660 4260
rect 5670 4250 5980 4260
rect 6370 4250 6520 4260
rect 6560 4250 6660 4260
rect 7040 4250 7050 4260
rect 7160 4250 7170 4260
rect 7390 4250 7410 4260
rect 8470 4250 8480 4260
rect 9730 4250 9750 4260
rect 9810 4250 9820 4260
rect 9830 4250 9850 4260
rect 9900 4250 9920 4260
rect 2920 4240 2930 4250
rect 3140 4240 3150 4250
rect 4190 4240 4330 4250
rect 4530 4240 4600 4250
rect 4850 4240 4910 4250
rect 5530 4240 5650 4250
rect 5690 4240 5990 4250
rect 6300 4240 6310 4250
rect 6370 4240 6520 4250
rect 6560 4240 6660 4250
rect 7050 4240 7080 4250
rect 7150 4240 7170 4250
rect 7360 4240 7370 4250
rect 8450 4240 8460 4250
rect 8470 4240 8480 4250
rect 8840 4240 8850 4250
rect 9730 4240 9740 4250
rect 2870 4230 2880 4240
rect 3190 4230 3200 4240
rect 4170 4230 4330 4240
rect 4530 4230 4600 4240
rect 4830 4230 4910 4240
rect 5540 4230 5650 4240
rect 5720 4230 5990 4240
rect 6070 4230 6080 4240
rect 6270 4230 6330 4240
rect 6360 4230 6520 4240
rect 6570 4230 6660 4240
rect 7090 4230 7120 4240
rect 7270 4230 7330 4240
rect 9720 4230 9730 4240
rect 9810 4230 9820 4240
rect 9870 4230 9880 4240
rect 9940 4230 9950 4240
rect 2910 4220 2920 4230
rect 3080 4220 3090 4230
rect 3140 4220 3150 4230
rect 4170 4220 4330 4230
rect 4520 4220 4600 4230
rect 4770 4220 4920 4230
rect 5480 4220 5490 4230
rect 5550 4220 5650 4230
rect 5720 4220 6110 4230
rect 6260 4220 6510 4230
rect 6580 4220 6670 4230
rect 7240 4220 7300 4230
rect 7390 4220 7450 4230
rect 9370 4220 9380 4230
rect 9710 4220 9720 4230
rect 9870 4220 9880 4230
rect 9930 4220 9940 4230
rect 3040 4210 3050 4220
rect 3070 4210 3100 4220
rect 3120 4210 3150 4220
rect 3180 4210 3190 4220
rect 3240 4210 3250 4220
rect 4160 4210 4270 4220
rect 4280 4210 4330 4220
rect 4510 4210 4590 4220
rect 4710 4210 4950 4220
rect 5550 4210 5650 4220
rect 5750 4210 5840 4220
rect 5910 4210 6120 4220
rect 6250 4210 6320 4220
rect 6330 4210 6500 4220
rect 6580 4210 6670 4220
rect 7150 4210 7170 4220
rect 7180 4210 7210 4220
rect 7230 4210 7280 4220
rect 7350 4210 7380 4220
rect 8830 4210 8840 4220
rect 9330 4210 9340 4220
rect 9680 4210 9710 4220
rect 9730 4210 9740 4220
rect 9870 4210 9880 4220
rect 9920 4210 9930 4220
rect 9950 4210 9960 4220
rect 3180 4200 3200 4210
rect 3240 4200 3250 4210
rect 4150 4200 4230 4210
rect 4300 4200 4350 4210
rect 4480 4200 4970 4210
rect 5560 4200 5660 4210
rect 5810 4200 5830 4210
rect 5920 4200 6150 4210
rect 6160 4200 6180 4210
rect 6210 4200 6240 4210
rect 6250 4200 6270 4210
rect 6290 4200 6490 4210
rect 6580 4200 6660 4210
rect 7230 4200 7340 4210
rect 7460 4200 7470 4210
rect 9310 4200 9320 4210
rect 9670 4200 9710 4210
rect 9720 4200 9750 4210
rect 9930 4200 9950 4210
rect 9960 4200 9970 4210
rect 3150 4190 3170 4200
rect 3180 4190 3210 4200
rect 3230 4190 3240 4200
rect 4150 4190 4220 4200
rect 4300 4190 4370 4200
rect 4480 4190 4980 4200
rect 5420 4190 5430 4200
rect 5570 4190 5660 4200
rect 5920 4190 6180 4200
rect 6190 4190 6280 4200
rect 6290 4190 6480 4200
rect 6560 4190 6670 4200
rect 7220 4190 7230 4200
rect 7270 4190 7290 4200
rect 9220 4190 9240 4200
rect 9270 4190 9280 4200
rect 9670 4190 9690 4200
rect 9720 4190 9780 4200
rect 9860 4190 9870 4200
rect 9900 4190 9910 4200
rect 9980 4190 9990 4200
rect 3110 4180 3130 4190
rect 3160 4180 3170 4190
rect 3190 4180 3200 4190
rect 4140 4180 4200 4190
rect 4330 4180 4370 4190
rect 4460 4180 4680 4190
rect 4690 4180 4800 4190
rect 4820 4180 4960 4190
rect 4970 4180 4990 4190
rect 5400 4180 5420 4190
rect 5570 4180 5670 4190
rect 5930 4180 6260 4190
rect 6280 4180 6290 4190
rect 6300 4180 6480 4190
rect 6580 4180 6670 4190
rect 7230 4180 7240 4190
rect 7310 4180 7320 4190
rect 9190 4180 9200 4190
rect 9320 4180 9340 4190
rect 9670 4180 9690 4190
rect 9710 4180 9760 4190
rect 9790 4180 9800 4190
rect 9850 4180 9880 4190
rect 3110 4170 3130 4180
rect 4120 4170 4190 4180
rect 4340 4170 4380 4180
rect 4460 4170 4670 4180
rect 4710 4170 5000 4180
rect 5400 4170 5420 4180
rect 5590 4170 5670 4180
rect 5920 4170 6170 4180
rect 6180 4170 6470 4180
rect 6580 4170 6670 4180
rect 7250 4170 7260 4180
rect 7330 4170 7340 4180
rect 8820 4170 8830 4180
rect 9280 4170 9290 4180
rect 9320 4170 9340 4180
rect 9660 4170 9700 4180
rect 9800 4170 9810 4180
rect 9870 4170 9890 4180
rect 3110 4160 3120 4170
rect 4110 4160 4210 4170
rect 4340 4160 4400 4170
rect 4420 4160 4640 4170
rect 4710 4160 5010 4170
rect 5420 4160 5440 4170
rect 5600 4160 5680 4170
rect 5920 4160 6460 4170
rect 6540 4160 6560 4170
rect 6580 4160 6670 4170
rect 7250 4160 7260 4170
rect 9210 4160 9230 4170
rect 9660 4160 9690 4170
rect 9790 4160 9820 4170
rect 9880 4160 9890 4170
rect 3180 4150 3200 4160
rect 3270 4150 3280 4160
rect 4110 4150 4180 4160
rect 4340 4150 4610 4160
rect 4720 4150 5010 4160
rect 5440 4150 5450 4160
rect 5610 4150 5690 4160
rect 5940 4150 6440 4160
rect 6540 4150 6560 4160
rect 6580 4150 6670 4160
rect 7360 4150 7370 4160
rect 7410 4150 7470 4160
rect 9260 4150 9280 4160
rect 9310 4150 9320 4160
rect 9650 4150 9680 4160
rect 9780 4150 9820 4160
rect 9890 4150 9900 4160
rect 9990 4150 9990 4160
rect 4100 4140 4190 4150
rect 4350 4140 4590 4150
rect 4720 4140 4770 4150
rect 4900 4140 5010 4150
rect 5450 4140 5460 4150
rect 5620 4140 5690 4150
rect 5950 4140 6430 4150
rect 6520 4140 6670 4150
rect 7390 4140 7470 4150
rect 9280 4140 9300 4150
rect 9630 4140 9660 4150
rect 9800 4140 9810 4150
rect 9820 4140 9860 4150
rect 9910 4140 9920 4150
rect 9940 4140 9950 4150
rect 3130 4130 3140 4140
rect 3270 4130 3280 4140
rect 4090 4130 4180 4140
rect 4350 4130 4580 4140
rect 4950 4130 4980 4140
rect 5450 4130 5460 4140
rect 5630 4130 5700 4140
rect 5950 4130 6420 4140
rect 6520 4130 6670 4140
rect 7430 4130 7450 4140
rect 8810 4130 8820 4140
rect 9630 4130 9650 4140
rect 9820 4130 9860 4140
rect 9990 4130 9990 4140
rect 3030 4120 3040 4130
rect 3250 4120 3260 4130
rect 3270 4120 3280 4130
rect 4090 4120 4170 4130
rect 4390 4120 4400 4130
rect 4410 4120 4560 4130
rect 5450 4120 5460 4130
rect 5490 4120 5500 4130
rect 5640 4120 5710 4130
rect 5950 4120 6410 4130
rect 6480 4120 6500 4130
rect 6520 4120 6670 4130
rect 9630 4120 9660 4130
rect 9840 4120 9870 4130
rect 9970 4120 9990 4130
rect 3140 4110 3170 4120
rect 3220 4110 3240 4120
rect 3260 4110 3280 4120
rect 4090 4110 4170 4120
rect 4420 4110 4550 4120
rect 5460 4110 5470 4120
rect 5490 4110 5500 4120
rect 5650 4110 5710 4120
rect 5950 4110 6400 4120
rect 6470 4110 6480 4120
rect 6490 4110 6500 4120
rect 6520 4110 6660 4120
rect 9630 4110 9650 4120
rect 9770 4110 9780 4120
rect 9800 4110 9820 4120
rect 9980 4110 9990 4120
rect 3200 4100 3220 4110
rect 3240 4100 3250 4110
rect 3270 4100 3280 4110
rect 4080 4100 4160 4110
rect 4440 4100 4550 4110
rect 5030 4100 5050 4110
rect 5490 4100 5500 4110
rect 5660 4100 5720 4110
rect 5730 4100 5780 4110
rect 5950 4100 6390 4110
rect 6460 4100 6470 4110
rect 6490 4100 6500 4110
rect 6510 4100 6660 4110
rect 9620 4100 9640 4110
rect 9760 4100 9790 4110
rect 3190 4090 3210 4100
rect 3260 4090 3270 4100
rect 4080 4090 4160 4100
rect 4440 4090 4540 4100
rect 4920 4090 5020 4100
rect 5030 4090 5060 4100
rect 5460 4090 5470 4100
rect 5680 4090 5800 4100
rect 5960 4090 6370 4100
rect 6440 4090 6460 4100
rect 6490 4090 6500 4100
rect 6510 4090 6650 4100
rect 7490 4090 7500 4100
rect 8800 4090 8810 4100
rect 9210 4090 9220 4100
rect 9610 4090 9620 4100
rect 9630 4090 9650 4100
rect 9710 4090 9870 4100
rect 9900 4090 9920 4100
rect 3080 4080 3130 4090
rect 3170 4080 3220 4090
rect 3240 4080 3270 4090
rect 4070 4080 4120 4090
rect 4140 4080 4160 4090
rect 4440 4080 4540 4090
rect 4880 4080 4930 4090
rect 5030 4080 5070 4090
rect 5440 4080 5450 4090
rect 5460 4080 5470 4090
rect 5490 4080 5500 4090
rect 5690 4080 5810 4090
rect 5960 4080 6360 4090
rect 6430 4080 6460 4090
rect 6490 4080 6500 4090
rect 6510 4080 6650 4090
rect 7520 4080 7550 4090
rect 9600 4080 9610 4090
rect 9650 4080 9690 4090
rect 9730 4080 9840 4090
rect 9890 4080 9940 4090
rect 3110 4070 3130 4080
rect 3180 4070 3220 4080
rect 3250 4070 3270 4080
rect 4060 4070 4120 4080
rect 4440 4070 4550 4080
rect 4830 4070 4840 4080
rect 4870 4070 4910 4080
rect 5030 4070 5080 4080
rect 5490 4070 5500 4080
rect 5710 4070 5840 4080
rect 5910 4070 5920 4080
rect 5930 4070 5940 4080
rect 5950 4070 6340 4080
rect 6420 4070 6460 4080
rect 6490 4070 6500 4080
rect 6510 4070 6650 4080
rect 7560 4070 7600 4080
rect 9200 4070 9210 4080
rect 9600 4070 9620 4080
rect 9630 4070 9760 4080
rect 9770 4070 9790 4080
rect 9910 4070 9940 4080
rect 3020 4060 3030 4070
rect 3140 4060 3150 4070
rect 3180 4060 3220 4070
rect 3250 4060 3260 4070
rect 4060 4060 4130 4070
rect 4210 4060 4220 4070
rect 4450 4060 4550 4070
rect 4820 4060 4830 4070
rect 4880 4060 4900 4070
rect 5020 4060 5080 4070
rect 5490 4060 5500 4070
rect 5720 4060 6320 4070
rect 6410 4060 6470 4070
rect 6490 4060 6500 4070
rect 6510 4060 6540 4070
rect 6560 4060 6660 4070
rect 6680 4060 6700 4070
rect 7600 4060 7640 4070
rect 9210 4060 9220 4070
rect 9590 4060 9610 4070
rect 9660 4060 9730 4070
rect 9930 4060 9990 4070
rect 3060 4050 3070 4060
rect 3090 4050 3110 4060
rect 3160 4050 3220 4060
rect 3250 4050 3270 4060
rect 4060 4050 4130 4060
rect 4170 4050 4180 4060
rect 4200 4050 4250 4060
rect 4470 4050 4540 4060
rect 4800 4050 4810 4060
rect 4870 4050 4900 4060
rect 5030 4050 5040 4060
rect 5050 4050 5080 4060
rect 5490 4050 5500 4060
rect 5730 4050 6310 4060
rect 6400 4050 6470 4060
rect 6490 4050 6500 4060
rect 6510 4050 6550 4060
rect 6570 4050 6690 4060
rect 7200 4050 7210 4060
rect 7630 4050 7640 4060
rect 7650 4050 7660 4060
rect 9210 4050 9220 4060
rect 9580 4050 9600 4060
rect 9950 4050 9990 4060
rect 2970 4040 2980 4050
rect 3070 4040 3100 4050
rect 3110 4040 3140 4050
rect 3170 4040 3180 4050
rect 3200 4040 3230 4050
rect 3240 4040 3250 4050
rect 4050 4040 4100 4050
rect 4170 4040 4270 4050
rect 4290 4040 4300 4050
rect 4470 4040 4540 4050
rect 4790 4040 4800 4050
rect 4870 4040 4900 4050
rect 5040 4040 5080 4050
rect 5490 4040 5500 4050
rect 5750 4040 6300 4050
rect 6390 4040 6480 4050
rect 6490 4040 6500 4050
rect 6510 4040 6540 4050
rect 6570 4040 6670 4050
rect 7190 4040 7200 4050
rect 7680 4040 7690 4050
rect 8630 4040 8640 4050
rect 8660 4040 8670 4050
rect 9210 4040 9220 4050
rect 9570 4040 9590 4050
rect 9970 4040 9990 4050
rect 3100 4030 3150 4040
rect 3180 4030 3230 4040
rect 3240 4030 3260 4040
rect 4050 4030 4090 4040
rect 4170 4030 4310 4040
rect 4480 4030 4540 4040
rect 4860 4030 4910 4040
rect 5030 4030 5090 4040
rect 5420 4030 5430 4040
rect 5490 4030 5500 4040
rect 5760 4030 6290 4040
rect 6390 4030 6480 4040
rect 6490 4030 6500 4040
rect 6510 4030 6540 4040
rect 6590 4030 6650 4040
rect 7180 4030 7200 4040
rect 7700 4030 7710 4040
rect 8550 4030 8610 4040
rect 9560 4030 9580 4040
rect 3120 4020 3160 4030
rect 3180 4020 3230 4030
rect 3240 4020 3270 4030
rect 4040 4020 4080 4030
rect 4150 4020 4170 4030
rect 4180 4020 4320 4030
rect 4480 4020 4550 4030
rect 4760 4020 4770 4030
rect 4830 4020 4910 4030
rect 5010 4020 5100 4030
rect 5420 4020 5430 4030
rect 5490 4020 5500 4030
rect 5820 4020 6250 4030
rect 6400 4020 6500 4030
rect 6520 4020 6590 4030
rect 6600 4020 6630 4030
rect 7160 4020 7200 4030
rect 7720 4020 7730 4030
rect 8560 4020 8620 4030
rect 9560 4020 9570 4030
rect 3120 4010 3170 4020
rect 3190 4010 3230 4020
rect 3240 4010 3260 4020
rect 4040 4010 4070 4020
rect 4170 4010 4330 4020
rect 4500 4010 4550 4020
rect 4740 4010 4750 4020
rect 4820 4010 4860 4020
rect 4880 4010 4900 4020
rect 5020 4010 5100 4020
rect 5410 4010 5430 4020
rect 5490 4010 5500 4020
rect 5910 4010 5920 4020
rect 5940 4010 6010 4020
rect 6020 4010 6240 4020
rect 6410 4010 6510 4020
rect 6580 4010 6610 4020
rect 7010 4010 7020 4020
rect 7130 4010 7150 4020
rect 7160 4010 7190 4020
rect 7730 4010 7740 4020
rect 7750 4010 7760 4020
rect 8450 4010 8460 4020
rect 8480 4010 8500 4020
rect 8540 4010 8550 4020
rect 8570 4010 8610 4020
rect 8690 4010 8700 4020
rect 8770 4010 8780 4020
rect 9550 4010 9560 4020
rect 3130 4000 3170 4010
rect 3190 4000 3200 4010
rect 3210 4000 3220 4010
rect 3240 4000 3260 4010
rect 4030 4000 4070 4010
rect 4160 4000 4330 4010
rect 4500 4000 4550 4010
rect 4790 4000 4840 4010
rect 4880 4000 4890 4010
rect 5020 4000 5100 4010
rect 5410 4000 5420 4010
rect 5490 4000 5500 4010
rect 5960 4000 5970 4010
rect 6010 4000 6080 4010
rect 6100 4000 6220 4010
rect 6400 4000 6580 4010
rect 7010 4000 7030 4010
rect 7140 4000 7180 4010
rect 7760 4000 7780 4010
rect 8470 4000 8490 4010
rect 8560 4000 8570 4010
rect 8580 4000 8620 4010
rect 8640 4000 8650 4010
rect 8710 4000 8720 4010
rect 3120 3990 3130 4000
rect 3150 3990 3170 4000
rect 3180 3990 3220 4000
rect 3260 3990 3270 4000
rect 4030 3990 4070 4000
rect 4150 3990 4340 4000
rect 4500 3990 4560 4000
rect 4770 3990 4810 4000
rect 4860 3990 4880 4000
rect 5060 3990 5110 4000
rect 5410 3990 5420 4000
rect 6110 3990 6130 4000
rect 6190 3990 6200 4000
rect 6400 3990 6580 4000
rect 7020 3990 7030 4000
rect 7130 3990 7170 4000
rect 7790 3990 7810 4000
rect 8350 3990 8360 4000
rect 8480 3990 8490 4000
rect 8520 3990 8530 4000
rect 8620 3990 8660 4000
rect 8720 3990 8730 4000
rect 3190 3980 3220 3990
rect 3240 3980 3250 3990
rect 3260 3980 3270 3990
rect 4020 3980 4050 3990
rect 4140 3980 4220 3990
rect 4250 3980 4350 3990
rect 4510 3980 4560 3990
rect 4610 3980 4620 3990
rect 4670 3980 4680 3990
rect 4710 3980 4730 3990
rect 4740 3980 4790 3990
rect 4850 3980 4860 3990
rect 5070 3980 5120 3990
rect 5450 3980 5470 3990
rect 5480 3980 5490 3990
rect 6400 3980 6580 3990
rect 7020 3980 7030 3990
rect 7130 3980 7160 3990
rect 7810 3980 7820 3990
rect 7830 3980 7840 3990
rect 8330 3980 8340 3990
rect 8450 3980 8460 3990
rect 8490 3980 8500 3990
rect 8620 3980 8700 3990
rect 8730 3980 8760 3990
rect 3140 3970 3150 3980
rect 3160 3970 3170 3980
rect 3200 3970 3230 3980
rect 3240 3970 3250 3980
rect 4010 3970 4050 3980
rect 4130 3970 4200 3980
rect 4280 3970 4350 3980
rect 4520 3970 4560 3980
rect 4580 3970 4630 3980
rect 4650 3970 4760 3980
rect 4840 3970 4850 3980
rect 5080 3970 5120 3980
rect 5410 3970 5490 3980
rect 6400 3970 6580 3980
rect 7020 3970 7040 3980
rect 7120 3970 7160 3980
rect 7840 3970 7870 3980
rect 8400 3970 8410 3980
rect 8450 3970 8480 3980
rect 8500 3970 8510 3980
rect 8570 3970 8580 3980
rect 8630 3970 8680 3980
rect 8700 3970 8710 3980
rect 8740 3970 8750 3980
rect 3140 3960 3150 3970
rect 3160 3960 3170 3970
rect 3200 3960 3210 3970
rect 3250 3960 3270 3970
rect 4010 3960 4040 3970
rect 4120 3960 4160 3970
rect 4290 3960 4350 3970
rect 4520 3960 4650 3970
rect 4660 3960 4720 3970
rect 4810 3960 4830 3970
rect 5100 3960 5130 3970
rect 5410 3960 5480 3970
rect 6400 3960 6580 3970
rect 7020 3960 7040 3970
rect 7110 3960 7160 3970
rect 7860 3960 7870 3970
rect 7880 3960 7890 3970
rect 8230 3960 8240 3970
rect 8270 3960 8280 3970
rect 8330 3960 8340 3970
rect 8440 3960 8490 3970
rect 8510 3960 8520 3970
rect 8560 3960 8580 3970
rect 8650 3960 8730 3970
rect 3130 3950 3160 3960
rect 3190 3950 3230 3960
rect 3260 3950 3270 3960
rect 3990 3950 4030 3960
rect 4100 3950 4150 3960
rect 4300 3950 4350 3960
rect 4530 3950 4650 3960
rect 4660 3950 4700 3960
rect 4790 3950 4810 3960
rect 5100 3950 5140 3960
rect 5420 3950 5430 3960
rect 5450 3950 5470 3960
rect 6400 3950 6580 3960
rect 7110 3950 7160 3960
rect 7890 3950 7910 3960
rect 8230 3950 8250 3960
rect 8290 3950 8300 3960
rect 8330 3950 8340 3960
rect 8480 3950 8490 3960
rect 8500 3950 8520 3960
rect 8660 3950 8670 3960
rect 8680 3950 8720 3960
rect 8730 3950 8750 3960
rect 3130 3940 3150 3950
rect 3190 3940 3200 3950
rect 3240 3940 3250 3950
rect 3260 3940 3270 3950
rect 3980 3940 4010 3950
rect 4100 3940 4140 3950
rect 4300 3940 4350 3950
rect 4530 3940 4700 3950
rect 4770 3940 4810 3950
rect 5120 3940 5150 3950
rect 6400 3940 6590 3950
rect 7110 3940 7160 3950
rect 7910 3940 7930 3950
rect 8140 3940 8270 3950
rect 8320 3940 8330 3950
rect 8640 3940 8650 3950
rect 8660 3940 8670 3950
rect 8680 3940 8690 3950
rect 8710 3940 8720 3950
rect 9650 3940 9670 3950
rect 9680 3940 9690 3950
rect 9720 3940 9730 3950
rect 9990 3940 9990 3950
rect 3140 3930 3160 3940
rect 3240 3930 3250 3940
rect 3960 3930 4000 3940
rect 4080 3930 4120 3940
rect 4310 3930 4360 3940
rect 4530 3930 4780 3940
rect 5130 3930 5160 3940
rect 6400 3930 6590 3940
rect 7120 3930 7150 3940
rect 7930 3930 7950 3940
rect 8120 3930 8200 3940
rect 8240 3930 8260 3940
rect 8280 3930 8290 3940
rect 8320 3930 8330 3940
rect 8340 3930 8350 3940
rect 8410 3930 8420 3940
rect 8460 3930 8470 3940
rect 8500 3930 8510 3940
rect 8560 3930 8580 3940
rect 8680 3930 8730 3940
rect 9660 3930 9680 3940
rect 9740 3930 9750 3940
rect 3180 3920 3200 3930
rect 3240 3920 3250 3930
rect 3950 3920 3980 3930
rect 4070 3920 4110 3930
rect 4320 3920 4360 3930
rect 4530 3920 4740 3930
rect 5140 3920 5170 3930
rect 6400 3920 6590 3930
rect 7140 3920 7150 3930
rect 7960 3920 7970 3930
rect 8040 3920 8050 3930
rect 8160 3920 8170 3930
rect 8180 3920 8190 3930
rect 8200 3920 8210 3930
rect 8250 3920 8260 3930
rect 8330 3920 8340 3930
rect 8430 3920 8440 3930
rect 8450 3920 8470 3930
rect 8560 3920 8570 3930
rect 8690 3920 8710 3930
rect 9610 3920 9630 3930
rect 9750 3920 9760 3930
rect 9940 3920 9950 3930
rect 3180 3910 3190 3920
rect 3220 3910 3260 3920
rect 3940 3910 3970 3920
rect 4060 3910 4090 3920
rect 4320 3910 4370 3920
rect 4530 3910 4660 3920
rect 4670 3910 4680 3920
rect 4690 3910 4700 3920
rect 5130 3910 5180 3920
rect 6410 3910 6600 3920
rect 7140 3910 7150 3920
rect 7970 3910 8010 3920
rect 8050 3910 8060 3920
rect 8200 3910 8210 3920
rect 8260 3910 8270 3920
rect 8310 3910 8320 3920
rect 8480 3910 8500 3920
rect 8510 3910 8520 3920
rect 9600 3910 9610 3920
rect 9770 3910 9780 3920
rect 3180 3900 3190 3910
rect 3220 3900 3240 3910
rect 3930 3900 3970 3910
rect 4050 3900 4090 3910
rect 4330 3900 4380 3910
rect 4540 3900 4630 3910
rect 5140 3900 5180 3910
rect 6410 3900 6600 3910
rect 8260 3900 8270 3910
rect 8330 3900 8340 3910
rect 8480 3900 8500 3910
rect 8710 3900 8720 3910
rect 3920 3890 3950 3900
rect 4020 3890 4080 3900
rect 4330 3890 4380 3900
rect 4540 3890 4640 3900
rect 5150 3890 5190 3900
rect 6410 3890 6600 3900
rect 7130 3890 7140 3900
rect 8060 3890 8070 3900
rect 8440 3890 8470 3900
rect 8540 3890 8550 3900
rect 8660 3890 8690 3900
rect 8710 3890 8720 3900
rect 9490 3890 9500 3900
rect 9550 3890 9560 3900
rect 9750 3890 9760 3900
rect 3140 3880 3220 3890
rect 3910 3880 3950 3890
rect 4000 3880 4050 3890
rect 4330 3880 4390 3890
rect 4550 3880 4640 3890
rect 5150 3880 5190 3890
rect 6420 3880 6600 3890
rect 8050 3880 8060 3890
rect 8270 3880 8280 3890
rect 8440 3880 8460 3890
rect 8470 3880 8480 3890
rect 8510 3880 8520 3890
rect 8610 3880 8620 3890
rect 8630 3880 8640 3890
rect 8650 3880 8670 3890
rect 8680 3880 8700 3890
rect 9470 3880 9480 3890
rect 9810 3880 9820 3890
rect 3120 3870 3180 3880
rect 3200 3870 3210 3880
rect 3270 3870 3280 3880
rect 3900 3870 3940 3880
rect 3990 3870 4040 3880
rect 4330 3870 4390 3880
rect 4550 3870 4650 3880
rect 5160 3870 5200 3880
rect 6430 3870 6600 3880
rect 8030 3870 8040 3880
rect 8220 3870 8230 3880
rect 8280 3870 8290 3880
rect 8340 3870 8350 3880
rect 8420 3870 8430 3880
rect 8480 3870 8490 3880
rect 8520 3870 8530 3880
rect 8560 3870 8670 3880
rect 8690 3870 8700 3880
rect 9440 3870 9460 3880
rect 9790 3870 9800 3880
rect 2940 3860 2950 3870
rect 3120 3860 3130 3870
rect 3140 3860 3150 3870
rect 3180 3860 3190 3870
rect 3200 3860 3220 3870
rect 3260 3860 3280 3870
rect 3900 3860 3930 3870
rect 3980 3860 4050 3870
rect 4340 3860 4400 3870
rect 4550 3860 4640 3870
rect 5160 3860 5200 3870
rect 6440 3860 6610 3870
rect 8230 3860 8240 3870
rect 8290 3860 8360 3870
rect 8420 3860 8430 3870
rect 8460 3860 8480 3870
rect 8530 3860 8580 3870
rect 8610 3860 8620 3870
rect 8640 3860 8650 3870
rect 8660 3860 8670 3870
rect 9770 3860 9780 3870
rect 9790 3860 9810 3870
rect 3090 3850 3140 3860
rect 3180 3850 3200 3860
rect 3260 3850 3280 3860
rect 3880 3850 3920 3860
rect 3970 3850 4060 3860
rect 4340 3850 4400 3860
rect 4580 3850 4640 3860
rect 5160 3850 5200 3860
rect 6500 3850 6610 3860
rect 8240 3850 8250 3860
rect 8310 3850 8370 3860
rect 8430 3850 8440 3860
rect 8550 3850 8570 3860
rect 8610 3850 8620 3860
rect 8670 3850 8700 3860
rect 9470 3850 9480 3860
rect 9550 3850 9560 3860
rect 9730 3850 9740 3860
rect 3080 3840 3100 3850
rect 3160 3840 3190 3850
rect 3260 3840 3270 3850
rect 3880 3840 3920 3850
rect 3960 3840 4060 3850
rect 4340 3840 4410 3850
rect 4590 3840 4640 3850
rect 5160 3840 5200 3850
rect 6510 3840 6610 3850
rect 8250 3840 8260 3850
rect 8320 3840 8410 3850
rect 8520 3840 8530 3850
rect 8570 3840 8620 3850
rect 8630 3840 8640 3850
rect 8650 3840 8680 3850
rect 9430 3840 9440 3850
rect 9880 3840 9890 3850
rect 3060 3830 3070 3840
rect 3160 3830 3170 3840
rect 3240 3830 3250 3840
rect 3880 3830 3920 3840
rect 3950 3830 4070 3840
rect 4340 3830 4410 3840
rect 4600 3830 4650 3840
rect 5160 3830 5210 3840
rect 6510 3830 6610 3840
rect 8250 3830 8270 3840
rect 8340 3830 8410 3840
rect 8460 3830 8470 3840
rect 8490 3830 8500 3840
rect 8530 3830 8550 3840
rect 8590 3830 8610 3840
rect 8620 3830 8650 3840
rect 8670 3830 8690 3840
rect 9590 3830 9600 3840
rect 9860 3830 9870 3840
rect 9890 3830 9900 3840
rect 3160 3820 3210 3830
rect 3250 3820 3260 3830
rect 3880 3820 3920 3830
rect 3950 3820 4060 3830
rect 4300 3820 4320 3830
rect 4330 3820 4410 3830
rect 4610 3820 4650 3830
rect 5160 3820 5220 3830
rect 6520 3820 6610 3830
rect 8240 3820 8270 3830
rect 8350 3820 8420 3830
rect 8430 3820 8450 3830
rect 8550 3820 8560 3830
rect 8590 3820 8600 3830
rect 8640 3820 8660 3830
rect 8680 3820 8690 3830
rect 9740 3820 9750 3830
rect 9820 3820 9830 3830
rect 3010 3810 3040 3820
rect 3120 3810 3130 3820
rect 3160 3810 3180 3820
rect 3200 3810 3210 3820
rect 3250 3810 3260 3820
rect 3880 3810 3920 3820
rect 3940 3810 4060 3820
rect 4300 3810 4420 3820
rect 5160 3810 5220 3820
rect 6530 3810 6610 3820
rect 8100 3810 8130 3820
rect 8240 3810 8260 3820
rect 8290 3810 8320 3820
rect 8360 3810 8440 3820
rect 8460 3810 8470 3820
rect 8520 3810 8530 3820
rect 8670 3810 8680 3820
rect 2990 3800 3070 3810
rect 3120 3800 3130 3810
rect 3200 3800 3210 3810
rect 3250 3800 3260 3810
rect 3880 3800 4040 3810
rect 4310 3800 4430 3810
rect 5160 3800 5230 3810
rect 6530 3800 6610 3810
rect 8110 3800 8130 3810
rect 8230 3800 8240 3810
rect 8270 3800 8280 3810
rect 8310 3800 8330 3810
rect 8380 3800 8440 3810
rect 8510 3800 8540 3810
rect 8620 3800 8630 3810
rect 2990 3790 3070 3800
rect 3100 3790 3130 3800
rect 3240 3790 3260 3800
rect 3890 3790 4030 3800
rect 4280 3790 4440 3800
rect 5160 3790 5220 3800
rect 6530 3790 6610 3800
rect 8300 3790 8360 3800
rect 8380 3790 8450 3800
rect 8520 3790 8540 3800
rect 8640 3790 8650 3800
rect 9830 3790 9840 3800
rect 2940 3780 3090 3790
rect 3110 3780 3130 3790
rect 3210 3780 3230 3790
rect 3260 3780 3270 3790
rect 3910 3780 4020 3790
rect 4260 3780 4270 3790
rect 4300 3780 4450 3790
rect 5150 3780 5220 3790
rect 6530 3780 6610 3790
rect 7060 3780 7070 3790
rect 8140 3780 8150 3790
rect 8250 3780 8320 3790
rect 8350 3780 8370 3790
rect 8420 3780 8430 3790
rect 8450 3780 8470 3790
rect 8640 3780 8670 3790
rect 9740 3780 9750 3790
rect 9820 3780 9850 3790
rect 2940 3770 2950 3780
rect 2970 3770 3050 3780
rect 3110 3770 3130 3780
rect 3230 3770 3250 3780
rect 3260 3770 3270 3780
rect 3920 3770 4000 3780
rect 4220 3770 4450 3780
rect 4870 3770 4900 3780
rect 5150 3770 5230 3780
rect 6540 3770 6610 3780
rect 8140 3770 8150 3780
rect 8220 3770 8260 3780
rect 8370 3770 8380 3780
rect 8520 3770 8530 3780
rect 8630 3770 8660 3780
rect 9730 3770 9750 3780
rect 9760 3770 9770 3780
rect 9860 3770 9890 3780
rect 2940 3760 3030 3770
rect 3050 3760 3080 3770
rect 3100 3760 3120 3770
rect 3260 3760 3270 3770
rect 3940 3760 3990 3770
rect 4200 3760 4210 3770
rect 4220 3760 4450 3770
rect 4840 3760 4930 3770
rect 5150 3760 5230 3770
rect 6530 3760 6610 3770
rect 8150 3760 8220 3770
rect 8380 3760 8390 3770
rect 8490 3760 8500 3770
rect 8530 3760 8540 3770
rect 8630 3760 8660 3770
rect 9730 3760 9740 3770
rect 9790 3760 9810 3770
rect 9900 3760 9910 3770
rect 2940 3750 3020 3760
rect 3040 3750 3060 3760
rect 3190 3750 3210 3760
rect 3220 3750 3240 3760
rect 3930 3750 3980 3760
rect 4200 3750 4450 3760
rect 4810 3750 4950 3760
rect 5140 3750 5240 3760
rect 6530 3750 6610 3760
rect 7040 3750 7050 3760
rect 8390 3750 8400 3760
rect 8510 3750 8520 3760
rect 8640 3750 8650 3760
rect 9790 3750 9800 3760
rect 2950 3740 3020 3750
rect 3030 3740 3060 3750
rect 3110 3740 3120 3750
rect 3210 3740 3250 3750
rect 3260 3740 3270 3750
rect 3930 3740 3970 3750
rect 4100 3740 4110 3750
rect 4180 3740 4440 3750
rect 4780 3740 4970 3750
rect 5130 3740 5240 3750
rect 6530 3740 6610 3750
rect 8170 3740 8180 3750
rect 8400 3740 8410 3750
rect 8520 3740 8530 3750
rect 8560 3740 8570 3750
rect 9670 3740 9680 3750
rect 9870 3740 9880 3750
rect 2990 3730 3070 3740
rect 3100 3730 3120 3740
rect 3180 3730 3190 3740
rect 3230 3730 3280 3740
rect 3920 3730 3950 3740
rect 4070 3730 4090 3740
rect 4160 3730 4220 3740
rect 4250 3730 4440 3740
rect 4780 3730 4990 3740
rect 5110 3730 5250 3740
rect 6540 3730 6610 3740
rect 8180 3730 8190 3740
rect 8410 3730 8430 3740
rect 9680 3730 9690 3740
rect 9870 3730 9880 3740
rect 9920 3730 9930 3740
rect 9980 3730 9990 3740
rect 2960 3720 3050 3730
rect 3110 3720 3120 3730
rect 3170 3720 3180 3730
rect 3220 3720 3260 3730
rect 3270 3720 3280 3730
rect 3910 3720 3940 3730
rect 4060 3720 4070 3730
rect 4140 3720 4200 3730
rect 4250 3720 4440 3730
rect 4780 3720 4850 3730
rect 4870 3720 5060 3730
rect 5080 3720 5270 3730
rect 6530 3720 6610 3730
rect 7020 3720 7030 3730
rect 8180 3720 8200 3730
rect 8430 3720 8440 3730
rect 8530 3720 8540 3730
rect 8590 3720 8600 3730
rect 9790 3720 9800 3730
rect 9820 3720 9830 3730
rect 9870 3720 9880 3730
rect 2910 3710 2920 3720
rect 3000 3710 3030 3720
rect 3040 3710 3080 3720
rect 3100 3710 3110 3720
rect 3180 3710 3250 3720
rect 3270 3710 3280 3720
rect 3890 3710 3950 3720
rect 4040 3710 4060 3720
rect 4130 3710 4180 3720
rect 4250 3710 4450 3720
rect 4780 3710 4830 3720
rect 4910 3710 5270 3720
rect 6540 3710 6610 3720
rect 8370 3710 8380 3720
rect 8440 3710 8460 3720
rect 9600 3710 9610 3720
rect 9700 3710 9710 3720
rect 9720 3710 9730 3720
rect 9960 3710 9990 3720
rect 3030 3700 3090 3710
rect 3110 3700 3160 3710
rect 3170 3700 3180 3710
rect 3190 3700 3260 3710
rect 3300 3700 3310 3710
rect 3880 3700 3940 3710
rect 4030 3700 4050 3710
rect 4080 3700 4150 3710
rect 4230 3700 4440 3710
rect 4810 3700 4840 3710
rect 4940 3700 5270 3710
rect 6540 3700 6610 3710
rect 8250 3700 8270 3710
rect 8290 3700 8350 3710
rect 8370 3700 8390 3710
rect 8460 3700 8470 3710
rect 9560 3700 9570 3710
rect 9590 3700 9620 3710
rect 9960 3700 9970 3710
rect 3060 3690 3090 3700
rect 3170 3690 3220 3700
rect 3250 3690 3270 3700
rect 3280 3690 3290 3700
rect 3300 3690 3310 3700
rect 3890 3690 3930 3700
rect 4020 3690 4050 3700
rect 4070 3690 4120 3700
rect 4220 3690 4260 3700
rect 4280 3690 4450 3700
rect 4810 3690 4850 3700
rect 4960 3690 5280 3700
rect 6550 3690 6600 3700
rect 7000 3690 7010 3700
rect 8200 3690 8210 3700
rect 8320 3690 8330 3700
rect 8370 3690 8390 3700
rect 8480 3690 8490 3700
rect 9540 3690 9570 3700
rect 9590 3690 9630 3700
rect 9830 3690 9840 3700
rect 9860 3690 9870 3700
rect 9940 3690 9970 3700
rect 3080 3680 3090 3690
rect 3180 3680 3220 3690
rect 3300 3680 3310 3690
rect 3890 3680 3920 3690
rect 4000 3680 4040 3690
rect 4060 3680 4090 3690
rect 4200 3680 4230 3690
rect 4310 3680 4440 3690
rect 4810 3680 4870 3690
rect 5000 3680 5280 3690
rect 6550 3680 6600 3690
rect 6990 3680 7000 3690
rect 8320 3680 8330 3690
rect 8360 3680 8380 3690
rect 8550 3680 8560 3690
rect 9520 3680 9550 3690
rect 9580 3680 9640 3690
rect 9830 3680 9840 3690
rect 3090 3670 3110 3680
rect 3120 3670 3140 3680
rect 3170 3670 3210 3680
rect 3240 3670 3260 3680
rect 3280 3670 3290 3680
rect 3310 3670 3320 3680
rect 3990 3670 4080 3680
rect 4180 3670 4220 3680
rect 4320 3670 4450 3680
rect 4810 3670 4880 3680
rect 5030 3670 5280 3680
rect 6550 3670 6600 3680
rect 6980 3670 6990 3680
rect 8390 3670 8400 3680
rect 8510 3670 8520 3680
rect 9510 3670 9520 3680
rect 9570 3670 9650 3680
rect 9840 3670 9850 3680
rect 9920 3670 9930 3680
rect 3110 3660 3170 3670
rect 3180 3660 3210 3670
rect 3230 3660 3290 3670
rect 3310 3660 3320 3670
rect 3980 3660 4070 3670
rect 4110 3660 4180 3670
rect 4320 3660 4440 3670
rect 4810 3660 4910 3670
rect 5100 3660 5290 3670
rect 6550 3660 6600 3670
rect 6960 3660 6980 3670
rect 8560 3660 8570 3670
rect 8590 3660 8610 3670
rect 9570 3660 9580 3670
rect 9620 3660 9660 3670
rect 3140 3650 3170 3660
rect 3180 3650 3200 3660
rect 3230 3650 3290 3660
rect 3970 3650 4100 3660
rect 4340 3650 4440 3660
rect 4810 3650 4920 3660
rect 5130 3650 5290 3660
rect 6540 3650 6600 3660
rect 6960 3650 6970 3660
rect 8310 3650 8320 3660
rect 8350 3650 8370 3660
rect 8380 3650 8390 3660
rect 8550 3650 8560 3660
rect 9550 3650 9570 3660
rect 9640 3650 9680 3660
rect 9930 3650 9940 3660
rect 3170 3640 3180 3650
rect 3240 3640 3260 3650
rect 3960 3640 4050 3650
rect 4340 3640 4420 3650
rect 4810 3640 4840 3650
rect 4870 3640 4940 3650
rect 5130 3640 5300 3650
rect 6540 3640 6590 3650
rect 6950 3640 6960 3650
rect 8320 3640 8340 3650
rect 8360 3640 8390 3650
rect 8550 3640 8570 3650
rect 9530 3640 9550 3650
rect 9650 3640 9680 3650
rect 9890 3640 9900 3650
rect 3190 3630 3200 3640
rect 3230 3630 3250 3640
rect 3270 3630 3290 3640
rect 3330 3630 3340 3640
rect 3960 3630 4040 3640
rect 4330 3630 4400 3640
rect 4800 3630 4850 3640
rect 4870 3630 4950 3640
rect 5130 3630 5290 3640
rect 6540 3630 6600 3640
rect 6950 3630 6960 3640
rect 8340 3630 8350 3640
rect 8360 3630 8370 3640
rect 8550 3630 8560 3640
rect 9520 3630 9540 3640
rect 9590 3630 9600 3640
rect 9660 3630 9690 3640
rect 9860 3630 9870 3640
rect 9910 3630 9920 3640
rect 3200 3620 3210 3630
rect 3240 3620 3250 3630
rect 3260 3620 3290 3630
rect 3950 3620 4040 3630
rect 4270 3620 4280 3630
rect 4330 3620 4420 3630
rect 4800 3620 4960 3630
rect 5130 3620 5300 3630
rect 6540 3620 6590 3630
rect 6940 3620 6950 3630
rect 8250 3620 8260 3630
rect 8340 3620 8370 3630
rect 8520 3620 8530 3630
rect 8550 3620 8560 3630
rect 9510 3620 9530 3630
rect 9580 3620 9620 3630
rect 9660 3620 9690 3630
rect 9900 3620 9910 3630
rect 9940 3620 9950 3630
rect 3210 3610 3230 3620
rect 3260 3610 3280 3620
rect 3940 3610 4050 3620
rect 4340 3610 4430 3620
rect 4800 3610 4970 3620
rect 5130 3610 5300 3620
rect 6530 3610 6590 3620
rect 6930 3610 6940 3620
rect 8340 3610 8360 3620
rect 9500 3610 9520 3620
rect 9570 3610 9650 3620
rect 9660 3610 9700 3620
rect 9940 3610 9950 3620
rect 3350 3600 3370 3610
rect 3930 3600 4050 3610
rect 4340 3600 4440 3610
rect 4780 3600 4850 3610
rect 4880 3600 4990 3610
rect 5130 3600 5300 3610
rect 6520 3600 6590 3610
rect 8340 3600 8360 3610
rect 8520 3600 8530 3610
rect 9460 3600 9500 3610
rect 9560 3600 9680 3610
rect 9690 3600 9700 3610
rect 9940 3600 9950 3610
rect 3300 3590 3310 3600
rect 3340 3590 3350 3600
rect 3930 3590 4060 3600
rect 4340 3590 4450 3600
rect 4730 3590 4740 3600
rect 4760 3590 4790 3600
rect 4820 3590 4850 3600
rect 4910 3590 5040 3600
rect 5130 3590 5300 3600
rect 6510 3590 6590 3600
rect 6920 3590 6930 3600
rect 8340 3590 8380 3600
rect 8420 3590 8430 3600
rect 9440 3590 9470 3600
rect 9550 3590 9580 3600
rect 9610 3590 9670 3600
rect 9680 3590 9690 3600
rect 9750 3590 9760 3600
rect 9990 3590 9990 3600
rect 3310 3580 3320 3590
rect 3930 3580 4060 3590
rect 4310 3580 4330 3590
rect 4350 3580 4470 3590
rect 4700 3580 4770 3590
rect 4820 3580 4850 3590
rect 4920 3580 4930 3590
rect 4970 3580 5060 3590
rect 5130 3580 5300 3590
rect 6510 3580 6580 3590
rect 6910 3580 6920 3590
rect 8300 3580 8310 3590
rect 8330 3580 8350 3590
rect 8360 3580 8370 3590
rect 8380 3580 8400 3590
rect 9300 3580 9370 3590
rect 9380 3580 9390 3590
rect 9400 3580 9410 3590
rect 9420 3580 9450 3590
rect 9540 3580 9560 3590
rect 9630 3580 9660 3590
rect 9730 3580 9740 3590
rect 9750 3580 9760 3590
rect 3260 3570 3270 3580
rect 3940 3570 4060 3580
rect 4310 3570 4470 3580
rect 4690 3570 4750 3580
rect 4810 3570 4850 3580
rect 4990 3570 5070 3580
rect 5140 3570 5300 3580
rect 6510 3570 6580 3580
rect 6900 3570 6910 3580
rect 8310 3570 8320 3580
rect 8360 3570 8390 3580
rect 8440 3570 8460 3580
rect 8500 3570 8510 3580
rect 9260 3570 9430 3580
rect 9540 3570 9550 3580
rect 9630 3570 9660 3580
rect 9670 3570 9680 3580
rect 9740 3570 9750 3580
rect 3260 3560 3290 3570
rect 3310 3560 3320 3570
rect 3350 3560 3360 3570
rect 3980 3560 4050 3570
rect 4290 3560 4480 3570
rect 4680 3560 4710 3570
rect 4720 3560 4730 3570
rect 4810 3560 4840 3570
rect 4990 3560 5080 3570
rect 5130 3560 5300 3570
rect 6510 3560 6580 3570
rect 8370 3560 8380 3570
rect 8400 3560 8420 3570
rect 8450 3560 8460 3570
rect 8500 3560 8510 3570
rect 8820 3560 8830 3570
rect 9250 3560 9410 3570
rect 9530 3560 9540 3570
rect 9630 3560 9670 3570
rect 9720 3560 9740 3570
rect 3270 3550 3280 3560
rect 3980 3550 4040 3560
rect 4280 3550 4490 3560
rect 4670 3550 4690 3560
rect 4810 3550 4840 3560
rect 5000 3550 5100 3560
rect 5140 3550 5300 3560
rect 6510 3550 6580 3560
rect 8330 3550 8340 3560
rect 8390 3550 8400 3560
rect 8410 3550 8420 3560
rect 8500 3550 8510 3560
rect 9230 3550 9300 3560
rect 9320 3550 9370 3560
rect 9510 3550 9530 3560
rect 9630 3550 9660 3560
rect 9710 3550 9720 3560
rect 3280 3540 3290 3550
rect 3330 3540 3340 3550
rect 3360 3540 3370 3550
rect 3380 3540 3390 3550
rect 3980 3540 4050 3550
rect 4270 3540 4490 3550
rect 4650 3540 4690 3550
rect 4790 3540 4830 3550
rect 5010 3540 5050 3550
rect 5070 3540 5110 3550
rect 5140 3540 5300 3550
rect 6500 3540 6590 3550
rect 6870 3540 6880 3550
rect 8410 3540 8420 3550
rect 8490 3540 8500 3550
rect 9210 3540 9280 3550
rect 9500 3540 9520 3550
rect 9630 3540 9650 3550
rect 9660 3540 9690 3550
rect 3300 3530 3310 3540
rect 3340 3530 3350 3540
rect 3990 3530 4050 3540
rect 4260 3530 4490 3540
rect 4630 3530 4680 3540
rect 4780 3530 4830 3540
rect 5000 3530 5040 3540
rect 5080 3530 5110 3540
rect 5140 3530 5300 3540
rect 6480 3530 6580 3540
rect 6870 3530 6880 3540
rect 8340 3530 8350 3540
rect 8490 3530 8500 3540
rect 9180 3530 9270 3540
rect 9480 3530 9500 3540
rect 9620 3530 9670 3540
rect 3320 3520 3330 3530
rect 3370 3520 3380 3530
rect 3390 3520 3400 3530
rect 3990 3520 4050 3530
rect 4260 3520 4340 3530
rect 4360 3520 4500 3530
rect 4600 3520 4670 3530
rect 4780 3520 4830 3530
rect 5000 3520 5020 3530
rect 5070 3520 5110 3530
rect 5130 3520 5310 3530
rect 6470 3520 6580 3530
rect 6860 3520 6870 3530
rect 8380 3520 8400 3530
rect 9180 3520 9260 3530
rect 9460 3520 9480 3530
rect 9590 3520 9630 3530
rect 3390 3510 3400 3520
rect 3990 3510 4060 3520
rect 4240 3510 4330 3520
rect 4370 3510 4530 3520
rect 4570 3510 4670 3520
rect 4780 3510 4820 3520
rect 4990 3510 5010 3520
rect 5070 3510 5310 3520
rect 6470 3510 6580 3520
rect 6850 3510 6860 3520
rect 8410 3510 8430 3520
rect 9170 3510 9230 3520
rect 9240 3510 9250 3520
rect 9440 3510 9460 3520
rect 9570 3510 9620 3520
rect 9640 3510 9660 3520
rect 3310 3500 3320 3510
rect 3380 3500 3390 3510
rect 3990 3500 4070 3510
rect 4220 3500 4320 3510
rect 4370 3500 4640 3510
rect 4770 3500 4820 3510
rect 4980 3500 4990 3510
rect 5060 3500 5310 3510
rect 6480 3500 6580 3510
rect 8380 3500 8390 3510
rect 8410 3500 8430 3510
rect 9150 3500 9210 3510
rect 9420 3500 9430 3510
rect 9570 3500 9600 3510
rect 9630 3500 9640 3510
rect 2490 3490 2590 3500
rect 3360 3490 3370 3500
rect 3390 3490 3410 3500
rect 3980 3490 4070 3500
rect 4210 3490 4300 3500
rect 4370 3490 4500 3500
rect 4570 3490 4600 3500
rect 4760 3490 4810 3500
rect 4960 3490 4980 3500
rect 5060 3490 5310 3500
rect 6480 3490 6580 3500
rect 6830 3490 6850 3500
rect 8410 3490 8440 3500
rect 9150 3490 9200 3500
rect 9390 3490 9410 3500
rect 9550 3490 9580 3500
rect 9630 3490 9640 3500
rect 2450 3480 2480 3490
rect 2510 3480 2530 3490
rect 2600 3480 2610 3490
rect 2620 3480 2640 3490
rect 2650 3480 2660 3490
rect 2670 3480 2680 3490
rect 3370 3480 3380 3490
rect 3980 3480 4070 3490
rect 4210 3480 4300 3490
rect 4380 3480 4490 3490
rect 4750 3480 4810 3490
rect 4950 3480 4960 3490
rect 5050 3480 5310 3490
rect 6470 3480 6570 3490
rect 6830 3480 6840 3490
rect 8410 3480 8420 3490
rect 8440 3480 8450 3490
rect 9130 3480 9190 3490
rect 9380 3480 9400 3490
rect 9540 3480 9570 3490
rect 9630 3480 9640 3490
rect 2410 3470 2420 3480
rect 2680 3470 2700 3480
rect 3330 3470 3340 3480
rect 3410 3470 3420 3480
rect 3990 3470 4070 3480
rect 4200 3470 4280 3480
rect 4390 3470 4480 3480
rect 4740 3470 4800 3480
rect 4930 3470 4940 3480
rect 5050 3470 5310 3480
rect 6460 3470 6570 3480
rect 6820 3470 6830 3480
rect 8420 3470 8430 3480
rect 8450 3470 8470 3480
rect 8530 3470 8550 3480
rect 9120 3470 9170 3480
rect 9340 3470 9410 3480
rect 9530 3470 9560 3480
rect 9620 3470 9640 3480
rect 2380 3460 2410 3470
rect 2710 3460 2750 3470
rect 2770 3460 2780 3470
rect 3410 3460 3420 3470
rect 4000 3460 4070 3470
rect 4190 3460 4270 3470
rect 4410 3460 4460 3470
rect 4740 3460 4800 3470
rect 4910 3460 4930 3470
rect 5040 3460 5050 3470
rect 5090 3460 5310 3470
rect 6450 3460 6570 3470
rect 8450 3460 8460 3470
rect 8470 3460 8480 3470
rect 8550 3460 8560 3470
rect 9100 3460 9160 3470
rect 9310 3460 9330 3470
rect 9380 3460 9430 3470
rect 9480 3460 9490 3470
rect 9500 3460 9540 3470
rect 9610 3460 9630 3470
rect 2360 3450 2370 3460
rect 2720 3450 2730 3460
rect 2750 3450 2760 3460
rect 2800 3450 2810 3460
rect 4000 3450 4080 3460
rect 4170 3450 4270 3460
rect 4420 3450 4440 3460
rect 4750 3450 4790 3460
rect 4880 3450 4910 3460
rect 5030 3450 5040 3460
rect 5110 3450 5310 3460
rect 6440 3450 6570 3460
rect 6800 3450 6810 3460
rect 8460 3450 8470 3460
rect 9090 3450 9160 3460
rect 9290 3450 9300 3460
rect 9420 3450 9530 3460
rect 9600 3450 9640 3460
rect 2320 3440 2350 3450
rect 2740 3440 2750 3450
rect 2830 3440 2870 3450
rect 4000 3440 4080 3450
rect 4150 3440 4270 3450
rect 4750 3440 4790 3450
rect 4850 3440 4880 3450
rect 5030 3440 5040 3450
rect 5120 3440 5150 3450
rect 5170 3440 5300 3450
rect 6380 3440 6390 3450
rect 6430 3440 6560 3450
rect 8470 3440 8490 3450
rect 9080 3440 9160 3450
rect 9270 3440 9280 3450
rect 9430 3440 9520 3450
rect 9600 3440 9610 3450
rect 2290 3430 2310 3440
rect 2740 3430 2750 3440
rect 2870 3430 2890 3440
rect 4000 3430 4080 3440
rect 4140 3430 4270 3440
rect 4360 3430 4380 3440
rect 4750 3430 4780 3440
rect 4830 3430 4860 3440
rect 5120 3430 5150 3440
rect 5180 3430 5300 3440
rect 6380 3430 6390 3440
rect 6430 3430 6560 3440
rect 6780 3430 6790 3440
rect 8490 3430 8500 3440
rect 9070 3430 9150 3440
rect 9250 3430 9260 3440
rect 9430 3430 9450 3440
rect 9460 3430 9510 3440
rect 9580 3430 9600 3440
rect 2260 3420 2290 3430
rect 2880 3420 2900 3430
rect 4000 3420 4090 3430
rect 4120 3420 4270 3430
rect 4350 3420 4390 3430
rect 4750 3420 4840 3430
rect 5120 3420 5150 3430
rect 5180 3420 5300 3430
rect 6370 3420 6380 3430
rect 6410 3420 6550 3430
rect 8540 3420 8550 3430
rect 9040 3420 9150 3430
rect 9230 3420 9240 3430
rect 9420 3420 9440 3430
rect 9470 3420 9510 3430
rect 9580 3420 9590 3430
rect 2250 3410 2280 3420
rect 4010 3410 4260 3420
rect 4350 3410 4390 3420
rect 4740 3410 4780 3420
rect 5130 3410 5150 3420
rect 5180 3410 5310 3420
rect 6400 3410 6550 3420
rect 6760 3410 6770 3420
rect 8540 3410 8550 3420
rect 9030 3410 9070 3420
rect 9220 3410 9230 3420
rect 9400 3410 9440 3420
rect 9480 3410 9510 3420
rect 9570 3410 9580 3420
rect 9650 3410 9670 3420
rect 2240 3400 2260 3410
rect 2880 3400 2970 3410
rect 4010 3400 4260 3410
rect 4350 3400 4420 3410
rect 4720 3400 4740 3410
rect 4940 3400 4980 3410
rect 5130 3400 5150 3410
rect 5180 3400 5300 3410
rect 6400 3400 6540 3410
rect 6750 3400 6760 3410
rect 9020 3400 9060 3410
rect 9210 3400 9220 3410
rect 9400 3400 9430 3410
rect 9560 3400 9570 3410
rect 9650 3400 9700 3410
rect 9770 3400 9780 3410
rect 2230 3390 2250 3400
rect 2810 3390 2830 3400
rect 2920 3390 2990 3400
rect 4010 3390 4260 3400
rect 4350 3390 4420 3400
rect 4700 3390 4740 3400
rect 4930 3390 4990 3400
rect 5130 3390 5150 3400
rect 5190 3390 5300 3400
rect 6380 3390 6530 3400
rect 6740 3390 6750 3400
rect 9010 3390 9070 3400
rect 9190 3390 9200 3400
rect 9400 3390 9420 3400
rect 9550 3390 9560 3400
rect 9650 3390 9700 3400
rect 2220 3380 2240 3390
rect 2980 3380 3000 3390
rect 4020 3380 4260 3390
rect 4360 3380 4430 3390
rect 4440 3380 4460 3390
rect 4470 3380 4480 3390
rect 4680 3380 4720 3390
rect 4910 3380 4940 3390
rect 4950 3380 4990 3390
rect 5140 3380 5150 3390
rect 5190 3380 5300 3390
rect 6380 3380 6530 3390
rect 8530 3380 8540 3390
rect 9020 3380 9090 3390
rect 9180 3380 9190 3390
rect 9400 3380 9430 3390
rect 9540 3380 9550 3390
rect 9650 3380 9710 3390
rect 2210 3370 2230 3380
rect 3010 3370 3020 3380
rect 3510 3370 3520 3380
rect 4020 3370 4250 3380
rect 4360 3370 4500 3380
rect 4650 3370 4710 3380
rect 4910 3370 4930 3380
rect 4960 3370 4990 3380
rect 5140 3370 5150 3380
rect 5190 3370 5300 3380
rect 6370 3370 6520 3380
rect 9030 3370 9100 3380
rect 9170 3370 9180 3380
rect 9410 3370 9420 3380
rect 9530 3370 9540 3380
rect 9660 3370 9700 3380
rect 9820 3370 9830 3380
rect 2190 3360 2210 3370
rect 3030 3360 3050 3370
rect 3510 3360 3530 3370
rect 4040 3360 4240 3370
rect 4360 3360 4520 3370
rect 4610 3360 4700 3370
rect 4900 3360 4930 3370
rect 4950 3360 5000 3370
rect 5190 3360 5300 3370
rect 6360 3360 6520 3370
rect 9060 3360 9080 3370
rect 9160 3360 9170 3370
rect 9410 3360 9430 3370
rect 9520 3360 9530 3370
rect 9660 3360 9720 3370
rect 2190 3350 2200 3360
rect 3050 3350 3060 3360
rect 3520 3350 3530 3360
rect 4060 3350 4070 3360
rect 4080 3350 4230 3360
rect 4360 3350 4430 3360
rect 4450 3350 4680 3360
rect 4880 3350 4930 3360
rect 4940 3350 4980 3360
rect 4990 3350 5000 3360
rect 5190 3350 5290 3360
rect 6340 3350 6520 3360
rect 8520 3350 8530 3360
rect 9060 3350 9080 3360
rect 9150 3350 9160 3360
rect 9410 3350 9440 3360
rect 9510 3350 9520 3360
rect 9650 3350 9730 3360
rect 2180 3340 2190 3350
rect 3060 3340 3070 3350
rect 3520 3340 3530 3350
rect 4150 3340 4230 3350
rect 4350 3340 4420 3350
rect 4480 3340 4630 3350
rect 4870 3340 4930 3350
rect 4940 3340 5000 3350
rect 5190 3340 5290 3350
rect 6340 3340 6520 3350
rect 9040 3340 9060 3350
rect 9400 3340 9430 3350
rect 9500 3340 9510 3350
rect 9640 3340 9720 3350
rect 2170 3330 2180 3340
rect 3070 3330 3080 3340
rect 3530 3330 3540 3340
rect 3580 3330 3590 3340
rect 4170 3330 4210 3340
rect 4350 3330 4410 3340
rect 4500 3330 4530 3340
rect 4540 3330 4580 3340
rect 4860 3330 4930 3340
rect 4940 3330 4990 3340
rect 5190 3330 5290 3340
rect 6340 3330 6510 3340
rect 6660 3330 6670 3340
rect 8510 3330 8520 3340
rect 8980 3330 9010 3340
rect 9330 3330 9430 3340
rect 9640 3330 9690 3340
rect 9700 3330 9720 3340
rect 2160 3320 2180 3330
rect 3080 3320 3090 3330
rect 3530 3320 3540 3330
rect 4170 3320 4190 3330
rect 4200 3320 4210 3330
rect 4350 3320 4410 3330
rect 4530 3320 4550 3330
rect 4850 3320 4920 3330
rect 4940 3320 4990 3330
rect 5190 3320 5290 3330
rect 6310 3320 6510 3330
rect 6650 3320 6660 3330
rect 8490 3320 8520 3330
rect 8940 3320 8980 3330
rect 9010 3320 9020 3330
rect 9330 3320 9420 3330
rect 9490 3320 9500 3330
rect 9630 3320 9660 3330
rect 2160 3310 2180 3320
rect 3090 3310 3100 3320
rect 3540 3310 3550 3320
rect 4180 3310 4190 3320
rect 4350 3310 4390 3320
rect 4510 3310 4540 3320
rect 4830 3310 4980 3320
rect 5010 3310 5020 3320
rect 5190 3310 5290 3320
rect 6300 3310 6520 3320
rect 6640 3310 6650 3320
rect 8510 3310 8520 3320
rect 8920 3310 9010 3320
rect 9020 3310 9050 3320
rect 9330 3310 9340 3320
rect 9370 3310 9410 3320
rect 9480 3310 9490 3320
rect 9630 3310 9650 3320
rect 2140 3300 2170 3310
rect 3100 3300 3110 3310
rect 3520 3300 3530 3310
rect 3540 3300 3580 3310
rect 4340 3300 4400 3310
rect 4490 3300 4520 3310
rect 4780 3300 4810 3310
rect 4820 3300 4920 3310
rect 4930 3300 4980 3310
rect 5010 3300 5020 3310
rect 5200 3300 5290 3310
rect 6240 3300 6270 3310
rect 6290 3300 6530 3310
rect 6630 3300 6650 3310
rect 8490 3300 8510 3310
rect 8920 3300 8970 3310
rect 9020 3300 9060 3310
rect 9470 3300 9490 3310
rect 9610 3300 9630 3310
rect 2140 3290 2170 3300
rect 3110 3290 3120 3300
rect 3520 3290 3530 3300
rect 4340 3290 4400 3300
rect 4410 3290 4420 3300
rect 4440 3290 4500 3300
rect 4760 3290 4810 3300
rect 4820 3290 4910 3300
rect 4930 3290 4970 3300
rect 5200 3290 5290 3300
rect 6250 3290 6520 3300
rect 6600 3290 6640 3300
rect 8920 3290 9040 3300
rect 9460 3290 9470 3300
rect 9600 3290 9620 3300
rect 9750 3290 9760 3300
rect 2130 3280 2150 3290
rect 3110 3280 3120 3290
rect 4340 3280 4480 3290
rect 4760 3280 4800 3290
rect 4810 3280 4900 3290
rect 4920 3280 4950 3290
rect 4960 3280 4970 3290
rect 5000 3280 5010 3290
rect 5200 3280 5290 3290
rect 6240 3280 6530 3290
rect 6580 3280 6590 3290
rect 6620 3280 6640 3290
rect 8860 3280 8950 3290
rect 8960 3280 8970 3290
rect 9010 3280 9030 3290
rect 9450 3280 9460 3290
rect 9590 3280 9610 3290
rect 9740 3280 9750 3290
rect 2120 3270 2150 3280
rect 4350 3270 4460 3280
rect 4750 3270 4900 3280
rect 4920 3270 4950 3280
rect 5000 3270 5010 3280
rect 5200 3270 5280 3280
rect 6240 3270 6520 3280
rect 6560 3270 6570 3280
rect 6620 3270 6640 3280
rect 8470 3270 8500 3280
rect 8830 3270 8930 3280
rect 8970 3270 9030 3280
rect 9070 3270 9080 3280
rect 9090 3270 9100 3280
rect 9320 3270 9330 3280
rect 9440 3270 9460 3280
rect 9560 3270 9600 3280
rect 9730 3270 9740 3280
rect 2120 3260 2140 3270
rect 3120 3260 3130 3270
rect 4370 3260 4430 3270
rect 4760 3260 4780 3270
rect 4790 3260 4900 3270
rect 4920 3260 4940 3270
rect 5000 3260 5010 3270
rect 5200 3260 5280 3270
rect 6250 3260 6520 3270
rect 6540 3260 6550 3270
rect 6610 3260 6630 3270
rect 8480 3260 8510 3270
rect 8820 3260 8900 3270
rect 8910 3260 8930 3270
rect 8990 3260 9030 3270
rect 9050 3260 9060 3270
rect 9090 3260 9100 3270
rect 9120 3260 9130 3270
rect 9310 3260 9330 3270
rect 9440 3260 9460 3270
rect 9520 3260 9580 3270
rect 9720 3260 9730 3270
rect 2120 3250 2130 3260
rect 3570 3250 3580 3260
rect 3590 3250 3600 3260
rect 4670 3250 4720 3260
rect 4780 3250 4900 3260
rect 4910 3250 4940 3260
rect 5000 3250 5010 3260
rect 5200 3250 5280 3260
rect 6250 3250 6530 3260
rect 6610 3250 6630 3260
rect 8830 3250 8890 3260
rect 8990 3250 9010 3260
rect 9120 3250 9130 3260
rect 9300 3250 9320 3260
rect 9330 3250 9340 3260
rect 9430 3250 9570 3260
rect 9710 3250 9720 3260
rect 2110 3240 2130 3250
rect 3130 3240 3140 3250
rect 3580 3240 3590 3250
rect 4660 3240 4730 3250
rect 4760 3240 4890 3250
rect 4900 3240 4940 3250
rect 4990 3240 5000 3250
rect 5200 3240 5280 3250
rect 6250 3240 6510 3250
rect 6610 3240 6620 3250
rect 8450 3240 8460 3250
rect 8830 3240 8850 3250
rect 8990 3240 9000 3250
rect 9080 3240 9090 3250
rect 9130 3240 9150 3250
rect 9290 3240 9310 3250
rect 9330 3240 9350 3250
rect 9420 3240 9520 3250
rect 2100 3230 2140 3240
rect 4660 3230 4920 3240
rect 4990 3230 5000 3240
rect 5200 3230 5270 3240
rect 6260 3230 6490 3240
rect 6610 3230 6620 3240
rect 9000 3230 9010 3240
rect 9080 3230 9090 3240
rect 9130 3230 9170 3240
rect 9280 3230 9300 3240
rect 9320 3230 9350 3240
rect 9420 3230 9490 3240
rect 9990 3230 9990 3240
rect 2100 3220 2140 3230
rect 3140 3220 3150 3230
rect 4660 3220 4680 3230
rect 4700 3220 4920 3230
rect 4980 3220 5000 3230
rect 5210 3220 5270 3230
rect 6270 3220 6480 3230
rect 6610 3220 6620 3230
rect 8950 3220 8960 3230
rect 8980 3220 8990 3230
rect 9070 3220 9080 3230
rect 9160 3220 9250 3230
rect 9270 3220 9290 3230
rect 9300 3220 9340 3230
rect 9410 3220 9480 3230
rect 9640 3220 9660 3230
rect 2090 3210 2140 3220
rect 3590 3210 3600 3220
rect 4650 3210 4910 3220
rect 4980 3210 5000 3220
rect 5210 3210 5260 3220
rect 6270 3210 6460 3220
rect 8920 3210 8940 3220
rect 8960 3210 8970 3220
rect 9060 3210 9070 3220
rect 9170 3210 9240 3220
rect 9250 3210 9280 3220
rect 9300 3210 9330 3220
rect 9400 3210 9470 3220
rect 9930 3210 9940 3220
rect 9970 3210 9980 3220
rect 2090 3200 2130 3210
rect 3150 3200 3160 3210
rect 4620 3200 4900 3210
rect 4970 3200 5000 3210
rect 5210 3200 5270 3210
rect 6290 3200 6430 3210
rect 8860 3200 8900 3210
rect 8930 3200 8940 3210
rect 9040 3200 9060 3210
rect 9190 3200 9200 3210
rect 9280 3200 9330 3210
rect 9400 3200 9470 3210
rect 9660 3200 9670 3210
rect 9910 3200 9960 3210
rect 2090 3190 2130 3200
rect 4600 3190 4890 3200
rect 4970 3190 5000 3200
rect 5210 3190 5270 3200
rect 6290 3190 6400 3200
rect 8760 3190 8820 3200
rect 8890 3190 8900 3200
rect 9010 3190 9040 3200
rect 9280 3190 9320 3200
rect 9390 3190 9460 3200
rect 9590 3190 9600 3200
rect 9640 3190 9670 3200
rect 9900 3190 9910 3200
rect 9930 3190 9940 3200
rect 2080 3180 2130 3190
rect 3160 3180 3170 3190
rect 4550 3180 4580 3190
rect 4590 3180 4860 3190
rect 4870 3180 4880 3190
rect 4960 3180 5010 3190
rect 5210 3180 5260 3190
rect 6290 3180 6360 3190
rect 8990 3180 9020 3190
rect 9280 3180 9290 3190
rect 9380 3180 9460 3190
rect 9600 3180 9640 3190
rect 9650 3180 9660 3190
rect 9940 3180 9950 3190
rect 2080 3170 2120 3180
rect 4240 3170 4250 3180
rect 4260 3170 4290 3180
rect 4570 3170 4580 3180
rect 4590 3170 4850 3180
rect 4860 3170 4880 3180
rect 4960 3170 5010 3180
rect 5210 3170 5260 3180
rect 6310 3170 6340 3180
rect 8960 3170 8980 3180
rect 9390 3170 9460 3180
rect 9550 3170 9560 3180
rect 9640 3170 9650 3180
rect 2080 3160 2120 3170
rect 4230 3160 4300 3170
rect 4370 3160 4380 3170
rect 4560 3160 4570 3170
rect 4590 3160 4620 3170
rect 4630 3160 4870 3170
rect 4950 3160 5010 3170
rect 5210 3160 5260 3170
rect 8910 3160 8950 3170
rect 9380 3160 9440 3170
rect 9550 3160 9590 3170
rect 9880 3160 9890 3170
rect 9960 3160 9970 3170
rect 2080 3150 2120 3160
rect 4230 3150 4310 3160
rect 4350 3150 4400 3160
rect 4560 3150 4580 3160
rect 4600 3150 4620 3160
rect 4630 3150 4860 3160
rect 4950 3150 5000 3160
rect 5210 3150 5260 3160
rect 8870 3150 8910 3160
rect 8950 3150 8980 3160
rect 9400 3150 9420 3160
rect 9550 3150 9590 3160
rect 9870 3150 9890 3160
rect 2080 3140 2120 3150
rect 3160 3140 3180 3150
rect 4230 3140 4320 3150
rect 4350 3140 4420 3150
rect 4570 3140 4590 3150
rect 4640 3140 4850 3150
rect 4940 3140 5000 3150
rect 5200 3140 5250 3150
rect 8800 3140 8810 3150
rect 8820 3140 8870 3150
rect 8930 3140 8970 3150
rect 9030 3140 9080 3150
rect 9560 3140 9600 3150
rect 9860 3140 9890 3150
rect 2080 3130 2110 3140
rect 3160 3130 3170 3140
rect 4230 3130 4330 3140
rect 4340 3130 4420 3140
rect 4430 3130 4440 3140
rect 4580 3130 4590 3140
rect 4650 3130 4830 3140
rect 4940 3130 5000 3140
rect 5200 3130 5250 3140
rect 8790 3130 8840 3140
rect 8890 3130 8950 3140
rect 9010 3130 9070 3140
rect 9560 3130 9570 3140
rect 9590 3130 9610 3140
rect 9880 3130 9920 3140
rect 2070 3120 2110 3130
rect 3160 3120 3170 3130
rect 4230 3120 4420 3130
rect 4450 3120 4460 3130
rect 4580 3120 4620 3130
rect 4650 3120 4820 3130
rect 4930 3120 4990 3130
rect 5190 3120 5250 3130
rect 8770 3120 8820 3130
rect 8840 3120 8880 3130
rect 8910 3120 8930 3130
rect 8990 3120 9060 3130
rect 9560 3120 9570 3130
rect 9840 3120 9850 3130
rect 9880 3120 9930 3130
rect 2070 3110 2110 3120
rect 3150 3110 3170 3120
rect 4240 3110 4420 3120
rect 4460 3110 4470 3120
rect 4590 3110 4770 3120
rect 4780 3110 4810 3120
rect 4930 3110 4980 3120
rect 5190 3110 5240 3120
rect 8720 3110 8780 3120
rect 8800 3110 8810 3120
rect 8900 3110 8920 3120
rect 8970 3110 9000 3120
rect 9020 3110 9050 3120
rect 9230 3110 9280 3120
rect 9550 3110 9570 3120
rect 9890 3110 9930 3120
rect 2070 3100 2110 3110
rect 3160 3100 3170 3110
rect 3860 3100 3870 3110
rect 3880 3100 3890 3110
rect 4240 3100 4430 3110
rect 4470 3100 4480 3110
rect 4600 3100 4630 3110
rect 4640 3100 4780 3110
rect 4930 3100 4990 3110
rect 5180 3100 5240 3110
rect 8380 3100 8390 3110
rect 8430 3100 8450 3110
rect 8870 3100 8900 3110
rect 8950 3100 8980 3110
rect 9010 3100 9040 3110
rect 9230 3100 9270 3110
rect 9280 3100 9290 3110
rect 9820 3100 9830 3110
rect 9930 3100 9940 3110
rect 2070 3090 2110 3100
rect 3160 3090 3170 3100
rect 3880 3090 3890 3100
rect 3900 3090 3910 3100
rect 4250 3090 4430 3100
rect 4480 3090 4490 3100
rect 4620 3090 4760 3100
rect 4920 3090 4990 3100
rect 5180 3090 5240 3100
rect 8380 3090 8390 3100
rect 8410 3090 8420 3100
rect 8860 3090 8880 3100
rect 8930 3090 8960 3100
rect 9010 3090 9030 3100
rect 9810 3090 9820 3100
rect 9890 3090 9900 3100
rect 9930 3090 9940 3100
rect 2070 3080 2110 3090
rect 3150 3080 3160 3090
rect 3900 3080 3910 3090
rect 4270 3080 4400 3090
rect 4410 3080 4460 3090
rect 4470 3080 4500 3090
rect 4920 3080 4980 3090
rect 5170 3080 5230 3090
rect 8440 3080 8450 3090
rect 8840 3080 8870 3090
rect 8910 3080 8950 3090
rect 9000 3080 9020 3090
rect 9520 3080 9530 3090
rect 9800 3080 9810 3090
rect 9890 3080 9900 3090
rect 9930 3080 9940 3090
rect 2060 3070 2110 3080
rect 3150 3070 3170 3080
rect 3900 3070 3910 3080
rect 4270 3070 4510 3080
rect 4910 3070 4980 3080
rect 5160 3070 5210 3080
rect 8390 3070 8400 3080
rect 8440 3070 8450 3080
rect 8830 3070 8880 3080
rect 8890 3070 8920 3080
rect 8970 3070 9000 3080
rect 9510 3070 9520 3080
rect 9790 3070 9800 3080
rect 9890 3070 9900 3080
rect 9960 3070 9970 3080
rect 2060 3060 2110 3070
rect 3140 3060 3160 3070
rect 4290 3060 4520 3070
rect 4900 3060 4990 3070
rect 5160 3060 5210 3070
rect 8420 3060 8430 3070
rect 8440 3060 8450 3070
rect 8790 3060 8910 3070
rect 8950 3060 8970 3070
rect 9510 3060 9520 3070
rect 2060 3050 2110 3060
rect 3140 3050 3150 3060
rect 3770 3050 3780 3060
rect 4300 3050 4530 3060
rect 4900 3050 5000 3060
rect 5150 3050 5210 3060
rect 8440 3050 8450 3060
rect 8760 3050 8870 3060
rect 8920 3050 8950 3060
rect 9510 3050 9530 3060
rect 9900 3050 9910 3060
rect 9990 3050 9990 3060
rect 2050 3040 2100 3050
rect 3130 3040 3150 3050
rect 3750 3040 3790 3050
rect 3890 3040 3910 3050
rect 4310 3040 4360 3050
rect 4400 3040 4530 3050
rect 4890 3040 5000 3050
rect 5130 3040 5210 3050
rect 8430 3040 8440 3050
rect 8720 3040 8730 3050
rect 8750 3040 8840 3050
rect 8900 3040 8930 3050
rect 9500 3040 9510 3050
rect 9900 3040 9910 3050
rect 2050 3030 2100 3040
rect 3130 3030 3150 3040
rect 3770 3030 3780 3040
rect 3880 3030 3920 3040
rect 4320 3030 4360 3040
rect 4400 3030 4530 3040
rect 4890 3030 5010 3040
rect 5120 3030 5210 3040
rect 8430 3030 8450 3040
rect 8640 3030 8650 3040
rect 8660 3030 8910 3040
rect 9500 3030 9510 3040
rect 2040 3020 2100 3030
rect 3130 3020 3150 3030
rect 3890 3020 3910 3030
rect 3920 3020 3930 3030
rect 4340 3020 4370 3030
rect 4410 3020 4470 3030
rect 4890 3020 5030 3030
rect 5080 3020 5090 3030
rect 5110 3020 5200 3030
rect 8440 3020 8450 3030
rect 8630 3020 8900 3030
rect 9490 3020 9500 3030
rect 9910 3020 9920 3030
rect 2040 3010 2090 3020
rect 3130 3010 3150 3020
rect 4350 3010 4380 3020
rect 4420 3010 4460 3020
rect 4890 3010 5100 3020
rect 5120 3010 5200 3020
rect 8340 3010 8350 3020
rect 8400 3010 8410 3020
rect 8440 3010 8450 3020
rect 8590 3010 8600 3020
rect 8620 3010 8880 3020
rect 8920 3010 8930 3020
rect 8940 3010 8950 3020
rect 9930 3010 9940 3020
rect 2040 3000 2090 3010
rect 3130 3000 3150 3010
rect 3870 3000 3880 3010
rect 3900 3000 3910 3010
rect 4360 3000 4390 3010
rect 4430 3000 4460 3010
rect 4890 3000 5190 3010
rect 8600 3000 8740 3010
rect 8770 3000 8900 3010
rect 9750 3000 9770 3010
rect 9940 3000 9960 3010
rect 2040 2990 2090 3000
rect 3130 2990 3150 3000
rect 3870 2990 3880 3000
rect 4370 2990 4410 3000
rect 4430 2990 4460 3000
rect 4880 2990 5190 3000
rect 8330 2990 8340 3000
rect 8450 2990 8460 3000
rect 8570 2990 8710 3000
rect 8850 2990 8910 3000
rect 9460 2990 9470 3000
rect 9770 2990 9780 3000
rect 9880 2990 9960 3000
rect 2040 2980 2080 2990
rect 3130 2980 3150 2990
rect 4090 2980 4100 2990
rect 4370 2980 4470 2990
rect 4900 2980 5190 2990
rect 8400 2980 8410 2990
rect 8560 2980 8710 2990
rect 8860 2980 8920 2990
rect 8940 2980 8950 2990
rect 9460 2980 9470 2990
rect 9790 2980 9800 2990
rect 9870 2980 9950 2990
rect 9960 2980 9970 2990
rect 2040 2970 2080 2980
rect 3120 2970 3140 2980
rect 3890 2970 3900 2980
rect 4000 2970 4010 2980
rect 4060 2970 4070 2980
rect 4390 2970 4480 2980
rect 4900 2970 5180 2980
rect 8550 2970 8710 2980
rect 8850 2970 8920 2980
rect 8930 2970 8950 2980
rect 9800 2970 9810 2980
rect 9830 2970 9870 2980
rect 9890 2970 9910 2980
rect 9940 2970 9960 2980
rect 2040 2960 2080 2970
rect 3120 2960 3140 2970
rect 3890 2960 3900 2970
rect 3990 2960 4000 2970
rect 4390 2960 4490 2970
rect 4910 2960 5180 2970
rect 8550 2960 8730 2970
rect 8750 2960 8760 2970
rect 8830 2960 8930 2970
rect 9810 2960 9820 2970
rect 9890 2960 9910 2970
rect 9940 2960 9950 2970
rect 2040 2950 2080 2960
rect 3120 2950 3130 2960
rect 3890 2950 3900 2960
rect 3980 2950 3990 2960
rect 4000 2950 4010 2960
rect 4050 2950 4060 2960
rect 4160 2950 4170 2960
rect 4420 2950 4500 2960
rect 4900 2950 5170 2960
rect 8550 2950 8900 2960
rect 8910 2950 8930 2960
rect 9690 2950 9720 2960
rect 9910 2950 9930 2960
rect 9940 2950 9950 2960
rect 2040 2940 2090 2950
rect 3120 2940 3130 2950
rect 3840 2940 3850 2950
rect 4150 2940 4160 2950
rect 4170 2940 4180 2950
rect 4430 2940 4510 2950
rect 4950 2940 5160 2950
rect 8300 2940 8310 2950
rect 8550 2940 8820 2950
rect 8890 2940 8910 2950
rect 9680 2940 9700 2950
rect 9730 2940 9740 2950
rect 9920 2940 9930 2950
rect 9950 2940 9960 2950
rect 2040 2930 2080 2940
rect 3110 2930 3140 2940
rect 3830 2930 3850 2940
rect 4000 2930 4010 2940
rect 4080 2930 4090 2940
rect 4440 2930 4520 2940
rect 4930 2930 5160 2940
rect 8550 2930 8750 2940
rect 9430 2930 9440 2940
rect 9680 2930 9700 2940
rect 9950 2930 9960 2940
rect 2040 2920 2080 2930
rect 3110 2920 3130 2930
rect 3910 2920 3930 2930
rect 3950 2920 3960 2930
rect 4100 2920 4110 2930
rect 4440 2920 4530 2930
rect 4930 2920 4940 2930
rect 4960 2920 5150 2930
rect 8540 2920 8690 2930
rect 9420 2920 9430 2930
rect 9670 2920 9700 2930
rect 2030 2910 2080 2920
rect 3110 2910 3130 2920
rect 4470 2910 4540 2920
rect 4930 2910 5150 2920
rect 8280 2910 8290 2920
rect 8500 2910 8670 2920
rect 9150 2910 9170 2920
rect 9660 2910 9720 2920
rect 2020 2900 2080 2910
rect 3100 2900 3130 2910
rect 4480 2900 4540 2910
rect 4940 2900 5120 2910
rect 5130 2900 5140 2910
rect 8500 2900 8640 2910
rect 9150 2900 9190 2910
rect 9410 2900 9420 2910
rect 9650 2900 9730 2910
rect 9900 2900 9970 2910
rect 2020 2890 2070 2900
rect 3100 2890 3130 2900
rect 4230 2890 4240 2900
rect 4490 2890 4540 2900
rect 4950 2890 4960 2900
rect 8270 2890 8280 2900
rect 8500 2890 8630 2900
rect 8790 2890 8800 2900
rect 8810 2890 8830 2900
rect 8860 2890 8880 2900
rect 9140 2890 9200 2900
rect 9640 2890 9730 2900
rect 9900 2890 9920 2900
rect 9960 2890 9980 2900
rect 2020 2880 2070 2890
rect 3100 2880 3120 2890
rect 4000 2880 4010 2890
rect 8260 2880 8270 2890
rect 8500 2880 8620 2890
rect 8710 2880 8880 2890
rect 9110 2880 9200 2890
rect 9390 2880 9400 2890
rect 9650 2880 9750 2890
rect 9920 2880 9930 2890
rect 9950 2880 9990 2890
rect 2020 2870 2070 2880
rect 3100 2870 3130 2880
rect 8500 2870 8620 2880
rect 8650 2870 8680 2880
rect 8690 2870 8840 2880
rect 9100 2870 9180 2880
rect 9660 2870 9740 2880
rect 9920 2870 9930 2880
rect 9940 2870 9960 2880
rect 2020 2860 2060 2870
rect 3110 2860 3150 2870
rect 7420 2860 7430 2870
rect 7480 2860 7490 2870
rect 8500 2860 8640 2870
rect 8650 2860 8800 2870
rect 9100 2860 9180 2870
rect 9360 2860 9370 2870
rect 9680 2860 9740 2870
rect 9950 2860 9970 2870
rect 2020 2850 2060 2860
rect 3110 2850 3150 2860
rect 7270 2850 7280 2860
rect 8240 2850 8250 2860
rect 8500 2850 8630 2860
rect 8710 2850 8740 2860
rect 8910 2850 8930 2860
rect 9090 2850 9180 2860
rect 9360 2850 9370 2860
rect 9690 2850 9740 2860
rect 9930 2850 9940 2860
rect 9950 2850 9970 2860
rect 2020 2840 2050 2850
rect 3110 2840 3150 2850
rect 8230 2840 8240 2850
rect 8510 2840 8620 2850
rect 8850 2840 8920 2850
rect 9080 2840 9180 2850
rect 9710 2840 9740 2850
rect 9940 2840 9990 2850
rect 2010 2830 2050 2840
rect 3090 2830 3100 2840
rect 3110 2830 3150 2840
rect 4080 2830 4100 2840
rect 4150 2830 4160 2840
rect 8520 2830 8610 2840
rect 8820 2830 8910 2840
rect 9070 2830 9180 2840
rect 9390 2830 9400 2840
rect 9720 2830 9750 2840
rect 9940 2830 9950 2840
rect 2010 2820 2040 2830
rect 3050 2820 3150 2830
rect 4070 2820 4080 2830
rect 4250 2820 4260 2830
rect 7210 2820 7220 2830
rect 8530 2820 8610 2830
rect 8790 2820 8910 2830
rect 9060 2820 9180 2830
rect 9230 2820 9260 2830
rect 9410 2820 9420 2830
rect 9600 2820 9610 2830
rect 9630 2820 9640 2830
rect 9660 2820 9670 2830
rect 9730 2820 9770 2830
rect 9970 2820 9980 2830
rect 2020 2810 2050 2820
rect 2900 2810 2920 2820
rect 3030 2810 3110 2820
rect 3990 2810 4000 2820
rect 4070 2810 4090 2820
rect 8210 2810 8220 2820
rect 8510 2810 8520 2820
rect 8530 2810 8610 2820
rect 8740 2810 8890 2820
rect 9060 2810 9160 2820
rect 9220 2810 9290 2820
rect 9360 2810 9370 2820
rect 9570 2810 9590 2820
rect 9600 2810 9610 2820
rect 9650 2810 9660 2820
rect 9680 2810 9690 2820
rect 9730 2810 9780 2820
rect 9920 2810 9930 2820
rect 9980 2810 9990 2820
rect 2010 2800 2060 2810
rect 2250 2800 2270 2810
rect 2290 2800 2390 2810
rect 2840 2800 2850 2810
rect 2860 2800 2970 2810
rect 2990 2800 3000 2810
rect 3010 2800 3100 2810
rect 3980 2800 3990 2810
rect 7550 2800 7560 2810
rect 8200 2800 8210 2810
rect 8500 2800 8620 2810
rect 8720 2800 8850 2810
rect 9060 2800 9150 2810
rect 9220 2800 9290 2810
rect 9350 2800 9360 2810
rect 9380 2800 9390 2810
rect 9590 2800 9600 2810
rect 9660 2800 9670 2810
rect 9760 2800 9780 2810
rect 9990 2800 9990 2810
rect 2010 2790 2080 2800
rect 2220 2790 2410 2800
rect 2810 2790 3100 2800
rect 4170 2790 4180 2800
rect 8500 2790 8620 2800
rect 8700 2790 8710 2800
rect 8720 2790 8800 2800
rect 9040 2790 9130 2800
rect 9220 2790 9290 2800
rect 9340 2790 9350 2800
rect 9400 2790 9410 2800
rect 9600 2790 9620 2800
rect 9950 2790 9990 2800
rect 2010 2780 2080 2790
rect 2220 2780 2430 2790
rect 2800 2780 3100 2790
rect 8500 2780 8630 2790
rect 8660 2780 8670 2790
rect 8680 2780 8760 2790
rect 9030 2780 9090 2790
rect 9200 2780 9210 2790
rect 9220 2780 9280 2790
rect 9380 2780 9430 2790
rect 9610 2780 9620 2790
rect 9670 2780 9680 2790
rect 9970 2780 9990 2790
rect 2000 2770 2080 2780
rect 2210 2770 2430 2780
rect 2790 2770 3100 2780
rect 4260 2770 4270 2780
rect 8510 2770 8630 2780
rect 8650 2770 8660 2780
rect 8670 2770 8730 2780
rect 9020 2770 9030 2780
rect 9050 2770 9070 2780
rect 9180 2770 9290 2780
rect 9330 2770 9340 2780
rect 9390 2770 9400 2780
rect 9410 2770 9440 2780
rect 9500 2770 9510 2780
rect 9680 2770 9690 2780
rect 2030 2760 2090 2770
rect 2200 2760 2440 2770
rect 2780 2760 3110 2770
rect 3940 2760 3950 2770
rect 4260 2760 4270 2770
rect 7610 2760 7620 2770
rect 8170 2760 8180 2770
rect 8530 2760 8640 2770
rect 9020 2760 9060 2770
rect 9170 2760 9180 2770
rect 9200 2760 9290 2770
rect 9420 2760 9470 2770
rect 9520 2760 9530 2770
rect 9710 2760 9730 2770
rect 9910 2760 9920 2770
rect 2040 2750 2080 2760
rect 2180 2750 2450 2760
rect 2780 2750 2990 2760
rect 3030 2750 3040 2760
rect 3100 2750 3110 2760
rect 3940 2750 3950 2760
rect 7620 2750 7630 2760
rect 8570 2750 8640 2760
rect 9010 2750 9020 2760
rect 9210 2750 9270 2760
rect 9420 2750 9460 2760
rect 9540 2750 9550 2760
rect 9700 2750 9730 2760
rect 9740 2750 9750 2760
rect 9900 2750 9910 2760
rect 2040 2740 2070 2750
rect 2220 2740 2460 2750
rect 2770 2740 2980 2750
rect 3100 2740 3140 2750
rect 3940 2740 3950 2750
rect 4170 2740 4190 2750
rect 4200 2740 4220 2750
rect 8150 2740 8160 2750
rect 8580 2740 8640 2750
rect 8980 2740 9030 2750
rect 9210 2740 9260 2750
rect 9310 2740 9320 2750
rect 9420 2740 9440 2750
rect 9500 2740 9510 2750
rect 9620 2740 9630 2750
rect 9720 2740 9750 2750
rect 9890 2740 9910 2750
rect 2030 2730 2080 2740
rect 2260 2730 2460 2740
rect 2770 2730 2950 2740
rect 3100 2730 3150 2740
rect 3930 2730 3940 2740
rect 4220 2730 4250 2740
rect 8570 2730 8660 2740
rect 8980 2730 9020 2740
rect 9210 2730 9230 2740
rect 9380 2730 9400 2740
rect 9420 2730 9430 2740
rect 9530 2730 9540 2740
rect 9590 2730 9600 2740
rect 9730 2730 9740 2740
rect 9890 2730 9900 2740
rect 2030 2720 2080 2730
rect 2270 2720 2470 2730
rect 2760 2720 2940 2730
rect 3110 2720 3150 2730
rect 3920 2720 3930 2730
rect 4210 2720 4250 2730
rect 8580 2720 8650 2730
rect 8980 2720 9000 2730
rect 9300 2720 9310 2730
rect 9380 2720 9390 2730
rect 9410 2720 9420 2730
rect 9550 2720 9560 2730
rect 9610 2720 9620 2730
rect 9690 2720 9700 2730
rect 9730 2720 9740 2730
rect 9890 2720 9900 2730
rect 2020 2710 2080 2720
rect 2280 2710 2470 2720
rect 2760 2710 2950 2720
rect 3110 2710 3150 2720
rect 4220 2710 4250 2720
rect 8550 2710 8650 2720
rect 8980 2710 8990 2720
rect 9290 2710 9300 2720
rect 9350 2710 9360 2720
rect 9570 2710 9580 2720
rect 9630 2710 9640 2720
rect 9660 2710 9670 2720
rect 9710 2710 9740 2720
rect 9810 2710 9820 2720
rect 9890 2710 9900 2720
rect 2020 2700 2050 2710
rect 2270 2700 2470 2710
rect 2750 2700 2950 2710
rect 3110 2700 3150 2710
rect 3920 2700 3930 2710
rect 4230 2700 4240 2710
rect 8560 2700 8650 2710
rect 9370 2700 9390 2710
rect 9590 2700 9600 2710
rect 9650 2700 9660 2710
rect 9710 2700 9730 2710
rect 9900 2700 9910 2710
rect 2020 2690 2050 2700
rect 2220 2690 2470 2700
rect 2750 2690 2800 2700
rect 2820 2690 2950 2700
rect 3110 2690 3130 2700
rect 3920 2690 3930 2700
rect 6980 2690 6990 2700
rect 7160 2690 7170 2700
rect 8110 2690 8120 2700
rect 8540 2690 8550 2700
rect 8560 2690 8640 2700
rect 9280 2690 9300 2700
rect 9610 2690 9620 2700
rect 9670 2690 9680 2700
rect 9910 2690 9930 2700
rect 2000 2680 2040 2690
rect 2200 2680 2480 2690
rect 2740 2680 2790 2690
rect 2830 2680 3060 2690
rect 3090 2680 3130 2690
rect 7160 2680 7170 2690
rect 8100 2680 8110 2690
rect 8510 2680 8530 2690
rect 8550 2680 8570 2690
rect 8580 2680 8640 2690
rect 9270 2680 9280 2690
rect 9630 2680 9640 2690
rect 9690 2680 9700 2690
rect 2000 2670 2030 2680
rect 2160 2670 2260 2680
rect 2410 2670 2480 2680
rect 2740 2670 2790 2680
rect 2860 2670 2920 2680
rect 2990 2670 3130 2680
rect 3910 2670 3920 2680
rect 6950 2670 6960 2680
rect 7160 2670 7170 2680
rect 8540 2670 8550 2680
rect 8560 2670 8570 2680
rect 8580 2670 8650 2680
rect 9710 2670 9720 2680
rect 9950 2670 9960 2680
rect 1990 2660 2030 2670
rect 2140 2660 2210 2670
rect 2420 2660 2480 2670
rect 2740 2660 2770 2670
rect 4240 2660 4250 2670
rect 7160 2660 7180 2670
rect 8520 2660 8560 2670
rect 8590 2660 8640 2670
rect 8780 2660 8830 2670
rect 9670 2660 9680 2670
rect 9730 2660 9740 2670
rect 9960 2660 9970 2670
rect 1990 2650 2020 2660
rect 2090 2650 2170 2660
rect 2440 2650 2480 2660
rect 2740 2650 2770 2660
rect 3910 2650 3920 2660
rect 4190 2650 4200 2660
rect 4260 2650 4270 2660
rect 7140 2650 7150 2660
rect 7170 2650 7190 2660
rect 8500 2650 8550 2660
rect 8590 2650 8660 2660
rect 8760 2650 8770 2660
rect 8790 2650 8850 2660
rect 9690 2650 9700 2660
rect 9750 2650 9760 2660
rect 9970 2650 9980 2660
rect 1990 2640 2030 2650
rect 2070 2640 2130 2650
rect 2440 2640 2480 2650
rect 2730 2640 2760 2650
rect 2970 2640 2980 2650
rect 3020 2640 3040 2650
rect 3910 2640 3930 2650
rect 4180 2640 4200 2650
rect 4260 2640 4270 2650
rect 7130 2640 7170 2650
rect 7180 2640 7190 2650
rect 8500 2640 8520 2650
rect 8530 2640 8550 2650
rect 8600 2640 8660 2650
rect 8750 2640 8770 2650
rect 8780 2640 8870 2650
rect 9210 2640 9220 2650
rect 9710 2640 9720 2650
rect 9770 2640 9780 2650
rect 9880 2640 9890 2650
rect 9930 2640 9940 2650
rect 9950 2640 9960 2650
rect 1980 2630 2110 2640
rect 2220 2630 2250 2640
rect 2440 2630 2480 2640
rect 2730 2630 2760 2640
rect 2940 2630 2970 2640
rect 3050 2630 3060 2640
rect 4190 2630 4200 2640
rect 4230 2630 4240 2640
rect 4260 2630 4270 2640
rect 7130 2630 7220 2640
rect 7240 2630 7250 2640
rect 7700 2630 7710 2640
rect 8430 2630 8470 2640
rect 8510 2630 8520 2640
rect 8540 2630 8550 2640
rect 8600 2630 8730 2640
rect 8740 2630 8890 2640
rect 9730 2630 9740 2640
rect 9790 2630 9800 2640
rect 9840 2630 9850 2640
rect 1980 2620 2090 2630
rect 2190 2620 2200 2630
rect 2250 2620 2270 2630
rect 2430 2620 2490 2630
rect 2730 2620 2760 2630
rect 2920 2620 2940 2630
rect 2980 2620 2990 2630
rect 3000 2620 3020 2630
rect 3030 2620 3080 2630
rect 3930 2620 3940 2630
rect 4190 2620 4200 2630
rect 7140 2620 7220 2630
rect 7240 2620 7260 2630
rect 8410 2620 8480 2630
rect 8520 2620 8560 2630
rect 8590 2620 8610 2630
rect 8620 2620 8900 2630
rect 9810 2620 9820 2630
rect 1970 2610 2070 2620
rect 2180 2610 2190 2620
rect 2200 2610 2220 2620
rect 2430 2610 2480 2620
rect 2730 2610 2760 2620
rect 3050 2610 3080 2620
rect 3940 2610 3950 2620
rect 4200 2610 4210 2620
rect 7130 2610 7230 2620
rect 7240 2610 7260 2620
rect 7270 2610 7280 2620
rect 8400 2610 8490 2620
rect 8530 2610 8570 2620
rect 8580 2610 8910 2620
rect 1970 2600 2060 2610
rect 2430 2600 2480 2610
rect 2730 2600 2760 2610
rect 3940 2600 3950 2610
rect 4200 2600 4210 2610
rect 7130 2600 7140 2610
rect 7150 2600 7200 2610
rect 7230 2600 7280 2610
rect 7720 2600 7730 2610
rect 8400 2600 8490 2610
rect 8550 2600 8870 2610
rect 8900 2600 8940 2610
rect 9190 2600 9200 2610
rect 9850 2600 9880 2610
rect 1970 2590 2040 2600
rect 2430 2590 2470 2600
rect 2730 2590 2770 2600
rect 2810 2590 2820 2600
rect 3940 2590 3950 2600
rect 4090 2590 4100 2600
rect 4200 2590 4210 2600
rect 4250 2590 4260 2600
rect 7130 2590 7200 2600
rect 7230 2590 7290 2600
rect 7730 2590 7740 2600
rect 8400 2590 8500 2600
rect 8560 2590 8860 2600
rect 8940 2590 8960 2600
rect 9190 2590 9200 2600
rect 9800 2590 9810 2600
rect 1970 2580 2040 2590
rect 2420 2580 2460 2590
rect 2730 2580 2810 2590
rect 3950 2580 3960 2590
rect 4190 2580 4200 2590
rect 4230 2580 4240 2590
rect 7100 2580 7150 2590
rect 7160 2580 7210 2590
rect 7240 2580 7270 2590
rect 7280 2580 7290 2590
rect 8400 2580 8490 2590
rect 8500 2580 8510 2590
rect 8520 2580 8540 2590
rect 8580 2580 8860 2590
rect 8940 2580 8970 2590
rect 9180 2580 9190 2590
rect 1940 2570 2020 2580
rect 2420 2570 2450 2580
rect 2730 2570 2830 2580
rect 3910 2570 3920 2580
rect 4040 2570 4050 2580
rect 4090 2570 4110 2580
rect 4180 2570 4220 2580
rect 4230 2570 4240 2580
rect 7100 2570 7160 2580
rect 7170 2570 7210 2580
rect 7250 2570 7270 2580
rect 7290 2570 7300 2580
rect 8400 2570 8870 2580
rect 8940 2570 9000 2580
rect 9320 2570 9330 2580
rect 1940 2560 2010 2570
rect 2420 2560 2430 2570
rect 2730 2560 2830 2570
rect 3930 2560 3950 2570
rect 4070 2560 4080 2570
rect 4100 2560 4110 2570
rect 4170 2560 4180 2570
rect 6840 2560 6850 2570
rect 7110 2560 7140 2570
rect 7160 2560 7170 2570
rect 7180 2560 7220 2570
rect 7290 2560 7310 2570
rect 7980 2560 7990 2570
rect 8400 2560 8490 2570
rect 8500 2560 8580 2570
rect 8630 2560 8880 2570
rect 8940 2560 8980 2570
rect 9000 2560 9020 2570
rect 9180 2560 9190 2570
rect 9310 2560 9320 2570
rect 9390 2560 9400 2570
rect 9940 2560 9960 2570
rect 1940 2550 2000 2560
rect 2420 2550 2430 2560
rect 2740 2550 2800 2560
rect 2890 2550 2900 2560
rect 4010 2550 4020 2560
rect 4030 2550 4040 2560
rect 4060 2550 4070 2560
rect 4150 2550 4160 2560
rect 6830 2550 6840 2560
rect 7120 2550 7140 2560
rect 7170 2550 7180 2560
rect 7190 2550 7220 2560
rect 7300 2550 7320 2560
rect 7970 2550 7980 2560
rect 8400 2550 8490 2560
rect 8500 2550 8580 2560
rect 8640 2550 8890 2560
rect 8930 2550 8980 2560
rect 9010 2550 9030 2560
rect 9180 2550 9190 2560
rect 9340 2550 9360 2560
rect 9420 2550 9430 2560
rect 9490 2550 9500 2560
rect 9960 2550 9970 2560
rect 9980 2550 9990 2560
rect 1940 2540 1990 2550
rect 2420 2540 2430 2550
rect 2740 2540 2790 2550
rect 2890 2540 2900 2550
rect 3990 2540 4010 2550
rect 4030 2540 4060 2550
rect 4070 2540 4080 2550
rect 4100 2540 4110 2550
rect 4120 2540 4160 2550
rect 6820 2540 6830 2550
rect 7130 2540 7160 2550
rect 7180 2540 7190 2550
rect 7210 2540 7230 2550
rect 7300 2540 7330 2550
rect 8390 2540 8580 2550
rect 8590 2540 8660 2550
rect 8670 2540 8890 2550
rect 8910 2540 8990 2550
rect 9340 2540 9350 2550
rect 9380 2540 9410 2550
rect 9470 2540 9480 2550
rect 1940 2530 1980 2540
rect 2750 2530 2760 2540
rect 2820 2530 2830 2540
rect 2950 2530 2970 2540
rect 3010 2530 3030 2540
rect 3040 2530 3110 2540
rect 3960 2530 3970 2540
rect 4050 2530 4060 2540
rect 4110 2530 4130 2540
rect 6810 2530 6820 2540
rect 6830 2530 6840 2540
rect 7160 2530 7180 2540
rect 7190 2530 7210 2540
rect 7230 2530 7240 2540
rect 7310 2530 7340 2540
rect 8390 2530 8670 2540
rect 8680 2530 8900 2540
rect 8910 2530 8990 2540
rect 9170 2530 9180 2540
rect 9480 2530 9520 2540
rect 9990 2530 9990 2540
rect 1940 2520 1970 2530
rect 2400 2520 2410 2530
rect 2840 2520 2860 2530
rect 2900 2520 2920 2530
rect 3100 2520 3140 2530
rect 3970 2520 4050 2530
rect 4060 2520 4070 2530
rect 4080 2520 4090 2530
rect 6800 2520 6810 2530
rect 6830 2520 6850 2530
rect 7210 2520 7250 2530
rect 7310 2520 7340 2530
rect 7780 2520 7790 2530
rect 8390 2520 8880 2530
rect 8890 2520 8990 2530
rect 9490 2520 9510 2530
rect 1950 2510 1970 2520
rect 2110 2510 2160 2520
rect 2240 2510 2250 2520
rect 2270 2510 2300 2520
rect 2380 2510 2390 2520
rect 2870 2510 2900 2520
rect 3120 2510 3190 2520
rect 3980 2510 4000 2520
rect 4010 2510 4020 2520
rect 4070 2510 4090 2520
rect 6830 2510 6850 2520
rect 7190 2510 7200 2520
rect 7220 2510 7260 2520
rect 7320 2510 7340 2520
rect 8390 2510 8690 2520
rect 8700 2510 8830 2520
rect 8860 2510 8870 2520
rect 8900 2510 8980 2520
rect 9160 2510 9170 2520
rect 9410 2510 9420 2520
rect 2010 2500 2020 2510
rect 2040 2500 2070 2510
rect 2090 2500 2120 2510
rect 2200 2500 2320 2510
rect 2350 2500 2370 2510
rect 3120 2500 3200 2510
rect 6820 2500 6830 2510
rect 6840 2500 6860 2510
rect 7210 2500 7220 2510
rect 7230 2500 7270 2510
rect 7330 2500 7350 2510
rect 7900 2500 7910 2510
rect 8390 2500 8830 2510
rect 8890 2500 8970 2510
rect 9160 2500 9170 2510
rect 9270 2500 9280 2510
rect 9430 2500 9440 2510
rect 9600 2500 9610 2510
rect 1980 2490 2000 2500
rect 2060 2490 2120 2500
rect 2230 2490 2360 2500
rect 3100 2490 3190 2500
rect 6780 2490 6790 2500
rect 6810 2490 6860 2500
rect 7220 2490 7230 2500
rect 7260 2490 7270 2500
rect 7330 2490 7360 2500
rect 8390 2490 8750 2500
rect 8760 2490 8840 2500
rect 8890 2490 8940 2500
rect 9150 2490 9160 2500
rect 9580 2490 9590 2500
rect 1950 2480 1980 2490
rect 2180 2480 2190 2490
rect 2200 2480 2310 2490
rect 3070 2480 3150 2490
rect 3200 2480 3210 2490
rect 6790 2480 6870 2490
rect 7230 2480 7240 2490
rect 7350 2480 7370 2490
rect 8390 2480 8780 2490
rect 8790 2480 8940 2490
rect 9140 2480 9160 2490
rect 1940 2470 1970 2480
rect 2190 2470 2250 2480
rect 2300 2470 2310 2480
rect 2920 2470 3130 2480
rect 3200 2470 3220 2480
rect 6770 2470 6870 2480
rect 7240 2470 7250 2480
rect 7350 2470 7380 2480
rect 7810 2470 7820 2480
rect 8390 2470 8770 2480
rect 8800 2470 8950 2480
rect 9130 2470 9160 2480
rect 9240 2470 9250 2480
rect 9720 2470 9730 2480
rect 1930 2460 1960 2470
rect 2280 2460 2330 2470
rect 2930 2460 3110 2470
rect 3190 2460 3230 2470
rect 6770 2460 6870 2470
rect 7250 2460 7260 2470
rect 7360 2460 7430 2470
rect 7820 2460 7830 2470
rect 8390 2460 8970 2470
rect 9100 2460 9160 2470
rect 1930 2450 1950 2460
rect 2060 2450 2140 2460
rect 2230 2450 2320 2460
rect 2960 2450 3070 2460
rect 3200 2450 3230 2460
rect 6760 2450 6880 2460
rect 7260 2450 7280 2460
rect 7360 2450 7440 2460
rect 8390 2450 9150 2460
rect 9480 2450 9490 2460
rect 1920 2440 1940 2450
rect 2060 2440 2140 2450
rect 2180 2440 2310 2450
rect 3200 2440 3240 2450
rect 6760 2440 6770 2450
rect 6800 2440 6890 2450
rect 7380 2440 7440 2450
rect 8390 2440 9150 2450
rect 9680 2440 9690 2450
rect 9740 2440 9750 2450
rect 9760 2440 9770 2450
rect 9780 2440 9790 2450
rect 1920 2430 1960 2440
rect 2100 2430 2140 2440
rect 2230 2430 2290 2440
rect 3210 2430 3240 2440
rect 6760 2430 6780 2440
rect 6810 2430 6910 2440
rect 7290 2430 7300 2440
rect 7390 2430 7420 2440
rect 7430 2430 7450 2440
rect 8390 2430 9160 2440
rect 9220 2430 9230 2440
rect 9500 2430 9520 2440
rect 1920 2420 1960 2430
rect 2130 2420 2270 2430
rect 3210 2420 3250 2430
rect 6850 2420 6920 2430
rect 7310 2420 7320 2430
rect 7430 2420 7450 2430
rect 8400 2420 9160 2430
rect 9210 2420 9220 2430
rect 9270 2420 9280 2430
rect 1910 2410 1960 2420
rect 2150 2410 2220 2420
rect 3210 2410 3240 2420
rect 6850 2410 6930 2420
rect 7330 2410 7340 2420
rect 7430 2410 7460 2420
rect 8390 2410 9160 2420
rect 9200 2410 9210 2420
rect 9220 2410 9230 2420
rect 9260 2410 9270 2420
rect 9340 2410 9360 2420
rect 9370 2410 9380 2420
rect 9390 2410 9400 2420
rect 9670 2410 9680 2420
rect 9690 2410 9700 2420
rect 9800 2410 9810 2420
rect 1910 2400 1970 2410
rect 3220 2400 3240 2410
rect 6870 2400 6970 2410
rect 7350 2400 7360 2410
rect 7440 2400 7470 2410
rect 8390 2400 8950 2410
rect 8960 2400 9160 2410
rect 9170 2400 9180 2410
rect 9240 2400 9250 2410
rect 9330 2400 9340 2410
rect 9390 2400 9400 2410
rect 9570 2400 9580 2410
rect 9810 2400 9820 2410
rect 1910 2390 1970 2400
rect 3220 2390 3250 2400
rect 6890 2390 6990 2400
rect 7440 2390 7480 2400
rect 8390 2390 9160 2400
rect 9520 2390 9550 2400
rect 9580 2390 9590 2400
rect 9670 2390 9680 2400
rect 1910 2380 1970 2390
rect 3220 2380 3250 2390
rect 6900 2380 7010 2390
rect 7020 2380 7040 2390
rect 7380 2380 7390 2390
rect 7450 2380 7490 2390
rect 8400 2380 9160 2390
rect 9260 2380 9270 2390
rect 9390 2380 9400 2390
rect 9460 2380 9470 2390
rect 9520 2380 9530 2390
rect 9570 2380 9580 2390
rect 9820 2380 9850 2390
rect 1910 2370 1970 2380
rect 3220 2370 3250 2380
rect 6900 2370 7090 2380
rect 7390 2370 7400 2380
rect 7460 2370 7500 2380
rect 8410 2370 8700 2380
rect 8710 2370 8740 2380
rect 8760 2370 8860 2380
rect 8900 2370 9150 2380
rect 9460 2370 9470 2380
rect 9580 2370 9590 2380
rect 9690 2370 9700 2380
rect 9820 2370 9830 2380
rect 1910 2360 1950 2370
rect 3230 2360 3260 2370
rect 6900 2360 7090 2370
rect 7410 2360 7420 2370
rect 7480 2360 7510 2370
rect 8420 2360 8670 2370
rect 8760 2360 8850 2370
rect 8860 2360 8870 2370
rect 8890 2360 9150 2370
rect 9330 2360 9340 2370
rect 9370 2360 9380 2370
rect 9470 2360 9480 2370
rect 1910 2350 1960 2360
rect 3230 2350 3260 2360
rect 6920 2350 7150 2360
rect 7420 2350 7430 2360
rect 7480 2350 7510 2360
rect 8430 2350 8510 2360
rect 8530 2350 8650 2360
rect 8760 2350 8870 2360
rect 8890 2350 9150 2360
rect 9210 2350 9220 2360
rect 9240 2350 9250 2360
rect 9310 2350 9320 2360
rect 9480 2350 9490 2360
rect 9570 2350 9590 2360
rect 9600 2350 9610 2360
rect 1900 2340 1950 2350
rect 3230 2340 3260 2350
rect 6940 2340 7170 2350
rect 7440 2340 7450 2350
rect 7490 2340 7520 2350
rect 8540 2340 8660 2350
rect 8750 2340 9140 2350
rect 9230 2340 9240 2350
rect 9640 2340 9650 2350
rect 9770 2340 9780 2350
rect 9790 2340 9800 2350
rect 9850 2340 9860 2350
rect 9920 2340 9930 2350
rect 1900 2330 1950 2340
rect 3230 2330 3260 2340
rect 6950 2330 6960 2340
rect 7010 2330 7180 2340
rect 7500 2330 7530 2340
rect 8560 2330 8660 2340
rect 8750 2330 8850 2340
rect 8860 2330 8930 2340
rect 8980 2330 9140 2340
rect 9280 2330 9290 2340
rect 9410 2330 9420 2340
rect 9430 2330 9440 2340
rect 9540 2330 9550 2340
rect 9770 2330 9800 2340
rect 9910 2330 9930 2340
rect 1900 2320 1940 2330
rect 3230 2320 3260 2330
rect 7030 2320 7210 2330
rect 7510 2320 7550 2330
rect 8370 2320 8380 2330
rect 8570 2320 8660 2330
rect 8750 2320 8840 2330
rect 8880 2320 8920 2330
rect 8980 2320 9140 2330
rect 9430 2320 9440 2330
rect 9500 2320 9510 2330
rect 9530 2320 9540 2330
rect 1900 2310 1930 2320
rect 3230 2310 3260 2320
rect 6750 2310 6760 2320
rect 7060 2310 7230 2320
rect 7540 2310 7590 2320
rect 8570 2310 8660 2320
rect 8740 2310 8830 2320
rect 8960 2310 9130 2320
rect 9220 2310 9230 2320
rect 9430 2310 9440 2320
rect 9830 2310 9840 2320
rect 1900 2300 1930 2310
rect 3240 2300 3260 2310
rect 7080 2300 7180 2310
rect 7200 2300 7240 2310
rect 7260 2300 7270 2310
rect 7560 2300 7590 2310
rect 8580 2300 8660 2310
rect 8720 2300 8830 2310
rect 8930 2300 9140 2310
rect 9360 2300 9370 2310
rect 9480 2300 9500 2310
rect 9830 2300 9840 2310
rect 1890 2290 1930 2300
rect 3240 2290 3270 2300
rect 6410 2290 6420 2300
rect 6750 2290 6760 2300
rect 7220 2290 7270 2300
rect 7330 2290 7340 2300
rect 7580 2290 7620 2300
rect 8590 2290 8660 2300
rect 8720 2290 8860 2300
rect 8900 2290 9140 2300
rect 9200 2290 9210 2300
rect 9480 2290 9490 2300
rect 9520 2290 9590 2300
rect 1880 2280 1930 2290
rect 3250 2280 3270 2290
rect 6410 2280 6420 2290
rect 7230 2280 7290 2290
rect 7320 2280 7340 2290
rect 7360 2280 7400 2290
rect 7490 2280 7500 2290
rect 7590 2280 7620 2290
rect 8590 2280 8670 2290
rect 8720 2280 8860 2290
rect 8870 2280 9140 2290
rect 9490 2280 9500 2290
rect 9570 2280 9580 2290
rect 1880 2270 1930 2280
rect 3250 2270 3270 2280
rect 6410 2270 6430 2280
rect 7260 2270 7290 2280
rect 7300 2270 7320 2280
rect 7330 2270 7420 2280
rect 7480 2270 7500 2280
rect 7610 2270 7630 2280
rect 8600 2270 8680 2280
rect 8690 2270 9150 2280
rect 9530 2270 9540 2280
rect 1880 2260 1930 2270
rect 3250 2260 3270 2270
rect 6400 2260 6430 2270
rect 6760 2260 6770 2270
rect 7280 2260 7320 2270
rect 7330 2260 7360 2270
rect 7400 2260 7430 2270
rect 7500 2260 7510 2270
rect 7620 2260 7630 2270
rect 8610 2260 9130 2270
rect 9540 2260 9550 2270
rect 9870 2260 9880 2270
rect 1870 2250 1930 2260
rect 3250 2250 3280 2260
rect 6400 2250 6440 2260
rect 6750 2250 6770 2260
rect 7290 2250 7320 2260
rect 7330 2250 7360 2260
rect 7410 2250 7440 2260
rect 7500 2250 7510 2260
rect 7630 2250 7640 2260
rect 8640 2250 8890 2260
rect 8910 2250 9010 2260
rect 9020 2250 9110 2260
rect 1870 2240 1910 2250
rect 2690 2240 2720 2250
rect 3250 2240 3280 2250
rect 6400 2240 6440 2250
rect 6760 2240 6780 2250
rect 7300 2240 7310 2250
rect 7390 2240 7430 2250
rect 7500 2240 7510 2250
rect 7630 2240 7650 2250
rect 8650 2240 8870 2250
rect 9030 2240 9080 2250
rect 9250 2240 9260 2250
rect 1870 2230 1910 2240
rect 2650 2230 2730 2240
rect 3250 2230 3280 2240
rect 6400 2230 6440 2240
rect 6760 2230 6780 2240
rect 7380 2230 7400 2240
rect 7420 2230 7430 2240
rect 7500 2230 7510 2240
rect 7640 2230 7660 2240
rect 8680 2230 8720 2240
rect 8800 2230 8860 2240
rect 9020 2230 9060 2240
rect 9270 2230 9280 2240
rect 1870 2220 1910 2230
rect 2490 2220 2510 2230
rect 2610 2220 2740 2230
rect 3250 2220 3280 2230
rect 6400 2220 6460 2230
rect 6760 2220 6790 2230
rect 7380 2220 7400 2230
rect 7500 2220 7510 2230
rect 7650 2220 7680 2230
rect 8830 2220 8850 2230
rect 8990 2220 9030 2230
rect 9300 2220 9310 2230
rect 9570 2220 9580 2230
rect 1870 2210 1910 2220
rect 2470 2210 2640 2220
rect 2690 2210 2750 2220
rect 3250 2210 3280 2220
rect 6400 2210 6440 2220
rect 6450 2210 6460 2220
rect 6760 2210 6790 2220
rect 7380 2210 7400 2220
rect 7490 2210 7510 2220
rect 7660 2210 7690 2220
rect 8840 2210 8870 2220
rect 8970 2210 8990 2220
rect 9320 2210 9330 2220
rect 9590 2210 9600 2220
rect 9810 2210 9820 2220
rect 9980 2210 9990 2220
rect 1870 2200 1910 2210
rect 2470 2200 2620 2210
rect 2700 2200 2770 2210
rect 2820 2200 2850 2210
rect 3250 2200 3280 2210
rect 6400 2200 6440 2210
rect 6780 2200 6800 2210
rect 7420 2200 7430 2210
rect 7480 2200 7510 2210
rect 7680 2200 7710 2210
rect 9350 2200 9360 2210
rect 9960 2200 9970 2210
rect 1870 2190 1910 2200
rect 2450 2190 2600 2200
rect 2750 2190 2860 2200
rect 3240 2190 3280 2200
rect 6390 2190 6440 2200
rect 6460 2190 6470 2200
rect 6770 2190 6820 2200
rect 7390 2190 7400 2200
rect 7410 2190 7430 2200
rect 7470 2190 7500 2200
rect 7690 2190 7730 2200
rect 9680 2190 9700 2200
rect 9950 2190 9960 2200
rect 1860 2180 1910 2190
rect 2280 2180 2310 2190
rect 2420 2180 2450 2190
rect 2490 2180 2580 2190
rect 2770 2180 2810 2190
rect 2820 2180 2860 2190
rect 3240 2180 3280 2190
rect 6390 2180 6440 2190
rect 6460 2180 6470 2190
rect 6770 2180 6800 2190
rect 7390 2180 7440 2190
rect 7450 2180 7490 2190
rect 7710 2180 7740 2190
rect 1860 2170 1910 2180
rect 2260 2170 2310 2180
rect 2350 2170 2430 2180
rect 2510 2170 2560 2180
rect 2840 2170 2860 2180
rect 3240 2170 3270 2180
rect 6390 2170 6460 2180
rect 6470 2170 6480 2180
rect 6770 2170 6810 2180
rect 6820 2170 6830 2180
rect 7390 2170 7420 2180
rect 7440 2170 7470 2180
rect 7730 2170 7750 2180
rect 9960 2170 9970 2180
rect 1860 2160 1910 2170
rect 2250 2160 2300 2170
rect 2350 2160 2420 2170
rect 2530 2160 2550 2170
rect 2840 2160 2860 2170
rect 3230 2160 3270 2170
rect 6390 2160 6450 2170
rect 6460 2160 6480 2170
rect 6770 2160 6820 2170
rect 7400 2160 7410 2170
rect 7450 2160 7460 2170
rect 7750 2160 7780 2170
rect 9980 2160 9990 2170
rect 1860 2150 1920 2160
rect 2240 2150 2300 2160
rect 2350 2150 2400 2160
rect 2830 2150 2840 2160
rect 3230 2150 3280 2160
rect 6390 2150 6450 2160
rect 6460 2150 6490 2160
rect 6770 2150 6820 2160
rect 7310 2150 7320 2160
rect 7750 2150 7840 2160
rect 9440 2150 9450 2160
rect 9570 2150 9580 2160
rect 9980 2150 9990 2160
rect 1860 2140 1920 2150
rect 2230 2140 2290 2150
rect 2360 2140 2380 2150
rect 2820 2140 2830 2150
rect 3230 2140 3280 2150
rect 6380 2140 6440 2150
rect 6460 2140 6480 2150
rect 6790 2140 6830 2150
rect 7840 2140 7850 2150
rect 9290 2140 9300 2150
rect 9460 2140 9470 2150
rect 9560 2140 9570 2150
rect 9940 2140 9950 2150
rect 9980 2140 9990 2150
rect 1860 2130 1930 2140
rect 2220 2130 2290 2140
rect 2360 2130 2390 2140
rect 2730 2130 2760 2140
rect 2800 2130 2820 2140
rect 3220 2130 3270 2140
rect 6380 2130 6440 2140
rect 6450 2130 6480 2140
rect 6790 2130 6850 2140
rect 6860 2130 6870 2140
rect 7310 2130 7320 2140
rect 9240 2130 9250 2140
rect 9310 2130 9320 2140
rect 9680 2130 9690 2140
rect 9910 2130 9920 2140
rect 1860 2120 1930 2130
rect 2220 2120 2280 2130
rect 2370 2120 2410 2130
rect 2660 2120 2800 2130
rect 3220 2120 3270 2130
rect 6380 2120 6440 2130
rect 6450 2120 6470 2130
rect 6790 2120 6870 2130
rect 7310 2120 7320 2130
rect 7860 2120 7870 2130
rect 8380 2120 8390 2130
rect 9500 2120 9510 2130
rect 9580 2120 9590 2130
rect 9690 2120 9710 2130
rect 1870 2110 1940 2120
rect 2210 2110 2270 2120
rect 2380 2110 2490 2120
rect 2520 2110 2560 2120
rect 2640 2110 2670 2120
rect 2740 2110 2770 2120
rect 3220 2110 3260 2120
rect 6380 2110 6430 2120
rect 6450 2110 6480 2120
rect 6790 2110 6870 2120
rect 7300 2110 7320 2120
rect 7860 2110 7880 2120
rect 9650 2110 9670 2120
rect 1870 2100 1930 2110
rect 2210 2100 2260 2110
rect 2400 2100 2430 2110
rect 2540 2100 2570 2110
rect 2630 2100 2640 2110
rect 3220 2100 3260 2110
rect 6380 2100 6430 2110
rect 6450 2100 6490 2110
rect 6780 2100 6890 2110
rect 7300 2100 7320 2110
rect 7870 2100 7880 2110
rect 9360 2100 9370 2110
rect 9610 2100 9620 2110
rect 1870 2090 1940 2100
rect 2200 2090 2260 2100
rect 2550 2090 2580 2100
rect 2600 2090 2620 2100
rect 3200 2090 3260 2100
rect 6390 2090 6430 2100
rect 6450 2090 6490 2100
rect 6790 2090 6860 2100
rect 6870 2090 6900 2100
rect 7310 2090 7320 2100
rect 7870 2090 7880 2100
rect 9370 2090 9380 2100
rect 1870 2080 1940 2090
rect 2180 2080 2250 2090
rect 3200 2080 3260 2090
rect 6380 2080 6490 2090
rect 6790 2080 6910 2090
rect 7300 2080 7320 2090
rect 7880 2080 7900 2090
rect 9350 2080 9360 2090
rect 9450 2080 9460 2090
rect 9700 2080 9710 2090
rect 1870 2070 1940 2080
rect 2180 2070 2240 2080
rect 3190 2070 3260 2080
rect 6380 2070 6430 2080
rect 6440 2070 6490 2080
rect 6800 2070 6920 2080
rect 7300 2070 7320 2080
rect 7890 2070 7900 2080
rect 8380 2070 8390 2080
rect 9690 2070 9700 2080
rect 1860 2060 1960 2070
rect 2170 2060 2230 2070
rect 3180 2060 3250 2070
rect 6390 2060 6500 2070
rect 6800 2060 6930 2070
rect 7300 2060 7320 2070
rect 7900 2060 8000 2070
rect 8380 2060 8390 2070
rect 9210 2060 9220 2070
rect 9270 2060 9300 2070
rect 9680 2060 9690 2070
rect 1860 2050 1960 2060
rect 2160 2050 2220 2060
rect 3170 2050 3250 2060
rect 6390 2050 6490 2060
rect 6800 2050 6950 2060
rect 7300 2050 7320 2060
rect 7900 2050 7960 2060
rect 8000 2050 8010 2060
rect 8380 2050 8390 2060
rect 9150 2050 9160 2060
rect 9210 2050 9230 2060
rect 9510 2050 9540 2060
rect 9550 2050 9600 2060
rect 9670 2050 9680 2060
rect 1860 2040 1980 2050
rect 2150 2040 2220 2050
rect 3160 2040 3240 2050
rect 6380 2040 6480 2050
rect 6800 2040 6970 2050
rect 7300 2040 7320 2050
rect 8380 2040 8390 2050
rect 9150 2040 9160 2050
rect 9480 2040 9490 2050
rect 9620 2040 9650 2050
rect 1860 2030 1990 2040
rect 2100 2030 2210 2040
rect 3150 2030 3240 2040
rect 6380 2030 6470 2040
rect 6810 2030 6980 2040
rect 7290 2030 7320 2040
rect 8380 2030 8390 2040
rect 8470 2030 8480 2040
rect 9140 2030 9150 2040
rect 9470 2030 9480 2040
rect 1860 2020 2000 2030
rect 2080 2020 2200 2030
rect 3130 2020 3230 2030
rect 6370 2020 6470 2030
rect 6820 2020 6980 2030
rect 7280 2020 7330 2030
rect 8000 2020 8010 2030
rect 8380 2020 8390 2030
rect 8440 2020 8510 2030
rect 9110 2020 9150 2030
rect 9340 2020 9350 2030
rect 9360 2020 9370 2030
rect 1860 2010 2010 2020
rect 2040 2010 2200 2020
rect 3120 2010 3230 2020
rect 6360 2010 6470 2020
rect 6820 2010 7010 2020
rect 7280 2010 7330 2020
rect 7990 2010 8000 2020
rect 8380 2010 8390 2020
rect 8440 2010 8520 2020
rect 9080 2010 9150 2020
rect 9210 2010 9280 2020
rect 9390 2010 9400 2020
rect 1870 2000 2010 2010
rect 2020 2000 2200 2010
rect 3120 2000 3230 2010
rect 6360 2000 6480 2010
rect 6830 2000 7020 2010
rect 7280 2000 7330 2010
rect 8380 2000 8390 2010
rect 8440 2000 8540 2010
rect 9070 2000 9090 2010
rect 9110 2000 9190 2010
rect 1860 1990 2190 2000
rect 3110 1990 3220 2000
rect 6360 1990 6480 2000
rect 6830 1990 7040 2000
rect 7280 1990 7320 2000
rect 8450 1990 8550 2000
rect 9110 1990 9140 2000
rect 1860 1980 2180 1990
rect 3110 1980 3220 1990
rect 6360 1980 6480 1990
rect 6830 1980 7050 1990
rect 7280 1980 7320 1990
rect 7980 1980 7990 1990
rect 8450 1980 8550 1990
rect 9080 1980 9100 1990
rect 9110 1980 9140 1990
rect 9650 1980 9660 1990
rect 9670 1980 9680 1990
rect 1860 1970 2180 1980
rect 3100 1970 3220 1980
rect 6360 1970 6410 1980
rect 6420 1970 6460 1980
rect 6830 1970 7070 1980
rect 7280 1970 7320 1980
rect 7810 1970 7840 1980
rect 8450 1970 8570 1980
rect 9060 1970 9130 1980
rect 1860 1960 2180 1970
rect 3110 1960 3220 1970
rect 6360 1960 6410 1970
rect 6430 1960 6470 1970
rect 6830 1960 7090 1970
rect 7270 1960 7330 1970
rect 7820 1960 7860 1970
rect 8450 1960 8590 1970
rect 9030 1960 9130 1970
rect 9670 1960 9680 1970
rect 9920 1960 9930 1970
rect 1850 1950 1860 1960
rect 1870 1950 2170 1960
rect 3100 1950 3220 1960
rect 6370 1950 6410 1960
rect 6430 1950 6470 1960
rect 6840 1950 7140 1960
rect 7160 1950 7180 1960
rect 7220 1950 7330 1960
rect 7830 1950 7870 1960
rect 8450 1950 8640 1960
rect 8660 1950 8670 1960
rect 8690 1950 8710 1960
rect 8870 1950 8890 1960
rect 8990 1950 9130 1960
rect 9670 1950 9680 1960
rect 1860 1940 2170 1950
rect 3110 1940 3220 1950
rect 6370 1940 6480 1950
rect 6830 1940 7140 1950
rect 7150 1940 7330 1950
rect 7840 1940 7890 1950
rect 7950 1940 7960 1950
rect 8450 1940 8770 1950
rect 8810 1940 9130 1950
rect 9660 1940 9670 1950
rect 9680 1940 9690 1950
rect 9850 1940 9860 1950
rect 9940 1940 9990 1950
rect 1860 1930 2170 1940
rect 3030 1930 3040 1940
rect 3110 1930 3220 1940
rect 4550 1930 4600 1940
rect 4790 1930 4800 1940
rect 4830 1930 4840 1940
rect 6380 1930 6480 1940
rect 6830 1930 7330 1940
rect 7840 1930 7890 1940
rect 8450 1930 8830 1940
rect 8900 1930 9130 1940
rect 9640 1930 9650 1940
rect 9850 1930 9860 1940
rect 9870 1930 9880 1940
rect 9990 1930 9990 1940
rect 1860 1920 2160 1930
rect 2650 1920 2720 1930
rect 3010 1920 3030 1930
rect 3110 1920 3230 1930
rect 4500 1920 4510 1930
rect 4590 1920 4600 1930
rect 4780 1920 4790 1930
rect 4850 1920 4860 1930
rect 6380 1920 6490 1930
rect 6830 1920 7330 1930
rect 7830 1920 7900 1930
rect 8450 1920 8800 1930
rect 8930 1920 9130 1930
rect 9680 1920 9690 1930
rect 9860 1920 9870 1930
rect 9910 1920 9920 1930
rect 9980 1920 9990 1930
rect 1860 1910 2160 1920
rect 2600 1910 2660 1920
rect 2690 1910 2760 1920
rect 2850 1910 2880 1920
rect 2890 1910 2900 1920
rect 2990 1910 3040 1920
rect 3110 1910 3250 1920
rect 4530 1910 4550 1920
rect 4800 1910 4810 1920
rect 5020 1910 5060 1920
rect 6390 1910 6470 1920
rect 6840 1910 7330 1920
rect 7840 1910 7910 1920
rect 8370 1910 8380 1920
rect 8450 1910 8690 1920
rect 8960 1910 9120 1920
rect 9600 1910 9610 1920
rect 9630 1910 9670 1920
rect 9880 1910 9890 1920
rect 1860 1900 2160 1910
rect 2450 1900 2600 1910
rect 2730 1900 2930 1910
rect 2980 1900 3030 1910
rect 3110 1900 3270 1910
rect 4400 1900 4410 1910
rect 4860 1900 4870 1910
rect 4970 1900 4980 1910
rect 5040 1900 5050 1910
rect 5100 1900 5110 1910
rect 6830 1900 7340 1910
rect 7850 1900 7910 1910
rect 8370 1900 8380 1910
rect 8450 1900 8680 1910
rect 8960 1900 9120 1910
rect 9590 1900 9600 1910
rect 9610 1900 9640 1910
rect 9670 1900 9680 1910
rect 9730 1900 9740 1910
rect 1860 1890 2160 1900
rect 2430 1890 2460 1900
rect 2740 1890 2950 1900
rect 2970 1890 3020 1900
rect 3110 1890 3270 1900
rect 4360 1890 4370 1900
rect 4400 1890 4410 1900
rect 4630 1890 4650 1900
rect 4770 1890 4780 1900
rect 4790 1890 4800 1900
rect 4970 1890 4980 1900
rect 5060 1890 5070 1900
rect 5130 1890 5140 1900
rect 6830 1890 7340 1900
rect 7850 1890 7910 1900
rect 8450 1890 8660 1900
rect 8980 1890 9120 1900
rect 9580 1890 9620 1900
rect 9670 1890 9680 1900
rect 9750 1890 9760 1900
rect 9960 1890 9970 1900
rect 1870 1880 2160 1890
rect 2410 1880 2450 1890
rect 2780 1880 2800 1890
rect 2820 1880 2950 1890
rect 2970 1880 3020 1890
rect 3110 1880 3270 1890
rect 4550 1880 4560 1890
rect 4570 1880 4580 1890
rect 4630 1880 4640 1890
rect 4980 1880 4990 1890
rect 6830 1880 7340 1890
rect 7850 1880 7920 1890
rect 8450 1880 8640 1890
rect 8990 1880 9120 1890
rect 9240 1880 9250 1890
rect 9580 1880 9610 1890
rect 1860 1870 2160 1880
rect 2390 1870 2430 1880
rect 2830 1870 2950 1880
rect 2970 1870 3010 1880
rect 3110 1870 3270 1880
rect 4330 1870 4340 1880
rect 4540 1870 4550 1880
rect 4630 1870 4640 1880
rect 4990 1870 5000 1880
rect 6830 1870 7340 1880
rect 7850 1870 7920 1880
rect 8450 1870 8630 1880
rect 8990 1870 9120 1880
rect 9140 1870 9150 1880
rect 9200 1870 9210 1880
rect 9250 1870 9260 1880
rect 9570 1870 9600 1880
rect 1870 1860 2170 1870
rect 2370 1860 2400 1870
rect 2840 1860 2950 1870
rect 3120 1860 3260 1870
rect 3270 1860 3280 1870
rect 4300 1860 4330 1870
rect 4380 1860 4390 1870
rect 4400 1860 4410 1870
rect 4490 1860 4500 1870
rect 4630 1860 4640 1870
rect 4760 1860 4770 1870
rect 4850 1860 4860 1870
rect 5010 1860 5020 1870
rect 5030 1860 5040 1870
rect 5090 1860 5120 1870
rect 5200 1860 5210 1870
rect 5230 1860 5240 1870
rect 5260 1860 5270 1870
rect 6840 1860 7340 1870
rect 7850 1860 7930 1870
rect 8450 1860 8630 1870
rect 8990 1860 9120 1870
rect 9300 1860 9310 1870
rect 9340 1860 9360 1870
rect 9420 1860 9430 1870
rect 9520 1860 9530 1870
rect 9980 1860 9990 1870
rect 1870 1850 2170 1860
rect 2230 1850 2280 1860
rect 2290 1850 2330 1860
rect 2340 1850 2390 1860
rect 2860 1850 2870 1860
rect 2890 1850 2950 1860
rect 3120 1850 3280 1860
rect 4290 1850 4300 1860
rect 4360 1850 4370 1860
rect 4380 1850 4390 1860
rect 4490 1850 4500 1860
rect 4630 1850 4640 1860
rect 4850 1850 4860 1860
rect 5180 1850 5190 1860
rect 5230 1850 5240 1860
rect 5290 1850 5300 1860
rect 6840 1850 7340 1860
rect 7850 1850 7920 1860
rect 8450 1850 8630 1860
rect 8980 1850 9120 1860
rect 9210 1850 9230 1860
rect 9250 1850 9290 1860
rect 9360 1850 9370 1860
rect 9970 1850 9980 1860
rect 1880 1840 2170 1850
rect 2210 1840 2370 1850
rect 2890 1840 2960 1850
rect 3120 1840 3280 1850
rect 4350 1840 4360 1850
rect 4630 1840 4640 1850
rect 4770 1840 4780 1850
rect 4850 1840 4860 1850
rect 5010 1840 5020 1850
rect 5030 1840 5040 1850
rect 5170 1840 5180 1850
rect 5260 1840 5270 1850
rect 5300 1840 5310 1850
rect 6830 1840 7340 1850
rect 7860 1840 7920 1850
rect 8360 1840 8370 1850
rect 8450 1840 8630 1850
rect 8980 1840 9110 1850
rect 9230 1840 9240 1850
rect 9770 1840 9780 1850
rect 1870 1830 2180 1840
rect 2200 1830 2350 1840
rect 2900 1830 2950 1840
rect 3130 1830 3270 1840
rect 4580 1830 4590 1840
rect 4630 1830 4640 1840
rect 5190 1830 5200 1840
rect 5310 1830 5320 1840
rect 6840 1830 7340 1840
rect 7860 1830 7930 1840
rect 8450 1830 8630 1840
rect 8960 1830 9110 1840
rect 9300 1830 9310 1840
rect 9370 1830 9380 1840
rect 9410 1830 9420 1840
rect 9690 1830 9700 1840
rect 9770 1830 9780 1840
rect 9960 1830 9970 1840
rect 1870 1820 2160 1830
rect 2190 1820 2320 1830
rect 2910 1820 2960 1830
rect 3130 1820 3270 1830
rect 4280 1820 4290 1830
rect 4490 1820 4500 1830
rect 4630 1820 4640 1830
rect 4810 1820 4820 1830
rect 4870 1820 4880 1830
rect 5160 1820 5170 1830
rect 5320 1820 5330 1830
rect 6400 1820 6410 1830
rect 6840 1820 7340 1830
rect 7850 1820 7940 1830
rect 8450 1820 8630 1830
rect 8950 1820 9110 1830
rect 9200 1820 9210 1830
rect 9280 1820 9290 1830
rect 9420 1820 9430 1830
rect 9690 1820 9700 1830
rect 9990 1820 9990 1830
rect 1880 1810 2150 1820
rect 2190 1810 2290 1820
rect 2900 1810 2950 1820
rect 3130 1810 3270 1820
rect 4280 1810 4290 1820
rect 4560 1810 4570 1820
rect 4590 1810 4600 1820
rect 4640 1810 4650 1820
rect 4760 1810 4770 1820
rect 4820 1810 4830 1820
rect 4870 1810 4880 1820
rect 5000 1810 5010 1820
rect 5310 1810 5320 1820
rect 6380 1810 6410 1820
rect 6840 1810 7340 1820
rect 7860 1810 7950 1820
rect 8460 1810 8630 1820
rect 8930 1810 9110 1820
rect 9300 1810 9330 1820
rect 9950 1810 9960 1820
rect 1890 1800 2140 1810
rect 2190 1800 2250 1810
rect 2810 1800 2930 1810
rect 3150 1800 3270 1810
rect 4490 1800 4500 1810
rect 4550 1800 4560 1810
rect 4580 1800 4590 1810
rect 4620 1800 4630 1810
rect 4740 1800 4750 1810
rect 5020 1800 5030 1810
rect 5050 1800 5060 1810
rect 5070 1800 5080 1810
rect 5150 1800 5160 1810
rect 5170 1800 5180 1810
rect 5330 1800 5340 1810
rect 6370 1800 6420 1810
rect 6840 1800 7340 1810
rect 7860 1800 7940 1810
rect 8460 1800 8620 1810
rect 8930 1800 9110 1810
rect 9280 1800 9290 1810
rect 9300 1800 9310 1810
rect 9320 1800 9370 1810
rect 9770 1800 9780 1810
rect 1880 1790 2080 1800
rect 2100 1790 2110 1800
rect 2200 1790 2240 1800
rect 2780 1790 2820 1800
rect 3150 1790 3260 1800
rect 4280 1790 4290 1800
rect 4370 1790 4390 1800
rect 4490 1790 4500 1800
rect 4630 1790 4640 1800
rect 4800 1790 4820 1800
rect 6370 1790 6420 1800
rect 6840 1790 7340 1800
rect 7850 1790 7940 1800
rect 8460 1790 8620 1800
rect 8930 1790 9110 1800
rect 9220 1790 9230 1800
rect 9260 1790 9270 1800
rect 9280 1790 9290 1800
rect 9320 1790 9340 1800
rect 9460 1790 9470 1800
rect 9600 1790 9620 1800
rect 9930 1790 9940 1800
rect 9970 1790 9980 1800
rect 1880 1780 2080 1790
rect 2190 1780 2260 1790
rect 2760 1780 2820 1790
rect 3160 1780 3260 1790
rect 4190 1780 4200 1790
rect 4280 1780 4290 1790
rect 4350 1780 4360 1790
rect 4370 1780 4400 1790
rect 4490 1780 4500 1790
rect 4620 1780 4630 1790
rect 4730 1780 4740 1790
rect 4750 1780 4760 1790
rect 4830 1780 4840 1790
rect 4990 1780 5000 1790
rect 5140 1780 5150 1790
rect 6370 1780 6420 1790
rect 6840 1780 7340 1790
rect 7860 1780 7940 1790
rect 8350 1780 8360 1790
rect 8470 1780 8620 1790
rect 8910 1780 9100 1790
rect 9240 1780 9250 1790
rect 9270 1780 9280 1790
rect 9310 1780 9340 1790
rect 9690 1780 9700 1790
rect 1880 1770 2050 1780
rect 2190 1770 2320 1780
rect 2330 1770 2360 1780
rect 2370 1770 2380 1780
rect 2630 1770 2650 1780
rect 2660 1770 2800 1780
rect 3160 1770 3260 1780
rect 4200 1770 4210 1780
rect 4280 1770 4290 1780
rect 4340 1770 4360 1780
rect 4490 1770 4500 1780
rect 4610 1770 4620 1780
rect 4830 1770 4840 1780
rect 5010 1770 5020 1780
rect 5060 1770 5070 1780
rect 5310 1770 5320 1780
rect 5410 1770 5420 1780
rect 5430 1770 5460 1780
rect 6370 1770 6420 1780
rect 6850 1770 7070 1780
rect 7080 1770 7090 1780
rect 7100 1770 7350 1780
rect 7860 1770 7930 1780
rect 8350 1770 8360 1780
rect 8480 1770 8620 1780
rect 8900 1770 9100 1780
rect 9230 1770 9240 1780
rect 9320 1770 9340 1780
rect 9690 1770 9700 1780
rect 9960 1770 9970 1780
rect 1890 1760 2040 1770
rect 2200 1760 2300 1770
rect 2360 1760 2400 1770
rect 2530 1760 2780 1770
rect 3170 1760 3250 1770
rect 4280 1760 4290 1770
rect 4490 1760 4500 1770
rect 4780 1760 4790 1770
rect 5040 1760 5050 1770
rect 5130 1760 5140 1770
rect 5250 1760 5260 1770
rect 5350 1760 5360 1770
rect 5400 1760 5410 1770
rect 5430 1760 5450 1770
rect 6360 1760 6410 1770
rect 6840 1760 7040 1770
rect 7110 1760 7350 1770
rect 7860 1760 7940 1770
rect 8490 1760 8500 1770
rect 8520 1760 8610 1770
rect 8920 1760 9100 1770
rect 9220 1760 9240 1770
rect 9360 1760 9370 1770
rect 9380 1760 9390 1770
rect 9420 1760 9430 1770
rect 9830 1760 9850 1770
rect 9920 1760 9930 1770
rect 9960 1760 9970 1770
rect 1890 1750 2030 1760
rect 2210 1750 2240 1760
rect 2370 1750 2430 1760
rect 2530 1750 2760 1760
rect 3170 1750 3260 1760
rect 4290 1750 4300 1760
rect 4490 1750 4500 1760
rect 4540 1750 4550 1760
rect 4560 1750 4570 1760
rect 4720 1750 4730 1760
rect 4740 1750 4750 1760
rect 4860 1750 4870 1760
rect 5130 1750 5140 1760
rect 5150 1750 5160 1760
rect 5300 1750 5310 1760
rect 5350 1750 5360 1760
rect 5450 1750 5460 1760
rect 5480 1750 5490 1760
rect 6370 1750 6410 1760
rect 6840 1750 7050 1760
rect 7110 1750 7350 1760
rect 7860 1750 7940 1760
rect 8490 1750 8610 1760
rect 8920 1750 9090 1760
rect 9210 1750 9230 1760
rect 9370 1750 9390 1760
rect 9410 1750 9420 1760
rect 9700 1750 9710 1760
rect 1900 1740 2030 1750
rect 2390 1740 2440 1750
rect 2500 1740 2730 1750
rect 3150 1740 3250 1750
rect 4370 1740 4380 1750
rect 4570 1740 4580 1750
rect 4620 1740 4630 1750
rect 4860 1740 4870 1750
rect 4880 1740 4890 1750
rect 4980 1740 4990 1750
rect 5380 1740 5390 1750
rect 5500 1740 5510 1750
rect 6370 1740 6410 1750
rect 6840 1740 7040 1750
rect 7120 1740 7350 1750
rect 7860 1740 7940 1750
rect 8500 1740 8610 1750
rect 8910 1740 9090 1750
rect 9390 1740 9420 1750
rect 9550 1740 9560 1750
rect 9830 1740 9840 1750
rect 9950 1740 9960 1750
rect 1900 1730 2040 1740
rect 2410 1730 2710 1740
rect 3150 1730 3240 1740
rect 4220 1730 4230 1740
rect 4360 1730 4370 1740
rect 4550 1730 4560 1740
rect 4710 1730 4720 1740
rect 4880 1730 4890 1740
rect 5000 1730 5010 1740
rect 5030 1730 5040 1740
rect 5120 1730 5130 1740
rect 5140 1730 5150 1740
rect 5290 1730 5300 1740
rect 5340 1730 5350 1740
rect 5380 1730 5390 1740
rect 5480 1730 5490 1740
rect 5510 1730 5520 1740
rect 6380 1730 6390 1740
rect 6840 1730 7020 1740
rect 7030 1730 7040 1740
rect 7130 1730 7350 1740
rect 7860 1730 7950 1740
rect 8340 1730 8350 1740
rect 8510 1730 8600 1740
rect 8910 1730 9090 1740
rect 9390 1730 9410 1740
rect 9570 1730 9580 1740
rect 9780 1730 9790 1740
rect 9910 1730 9920 1740
rect 1900 1720 2020 1730
rect 2030 1720 2040 1730
rect 2440 1720 2690 1730
rect 3140 1720 3240 1730
rect 4180 1720 4230 1730
rect 4880 1720 4890 1730
rect 5260 1720 5270 1730
rect 5370 1720 5380 1730
rect 5490 1720 5500 1730
rect 5520 1720 5530 1730
rect 6840 1720 7010 1730
rect 7150 1720 7350 1730
rect 7860 1720 7950 1730
rect 8340 1720 8350 1730
rect 8500 1720 8600 1730
rect 8900 1720 9090 1730
rect 9540 1720 9580 1730
rect 9790 1720 9800 1730
rect 9860 1720 9870 1730
rect 9930 1720 9940 1730
rect 1910 1710 2020 1720
rect 2030 1710 2040 1720
rect 2460 1710 2670 1720
rect 3140 1710 3240 1720
rect 4070 1710 4090 1720
rect 4150 1710 4230 1720
rect 4290 1710 4300 1720
rect 4760 1710 4770 1720
rect 4990 1710 5000 1720
rect 5110 1710 5120 1720
rect 5250 1710 5260 1720
rect 5280 1710 5290 1720
rect 5390 1710 5400 1720
rect 6850 1710 7010 1720
rect 7150 1710 7350 1720
rect 7860 1710 7950 1720
rect 8500 1710 8610 1720
rect 8870 1710 9090 1720
rect 9200 1710 9220 1720
rect 9320 1710 9330 1720
rect 9650 1710 9660 1720
rect 9700 1710 9710 1720
rect 1920 1700 2020 1710
rect 2030 1700 2050 1710
rect 2480 1700 2580 1710
rect 2600 1700 2660 1710
rect 3130 1700 3230 1710
rect 4070 1700 4100 1710
rect 4120 1700 4240 1710
rect 4290 1700 4300 1710
rect 4490 1700 4500 1710
rect 4570 1700 4580 1710
rect 4700 1700 4710 1710
rect 4720 1700 4730 1710
rect 4810 1700 4820 1710
rect 5130 1700 5140 1710
rect 5220 1700 5230 1710
rect 5320 1700 5330 1710
rect 5360 1700 5370 1710
rect 5430 1700 5440 1710
rect 6840 1700 7010 1710
rect 7120 1700 7350 1710
rect 7860 1700 7950 1710
rect 8510 1700 8610 1710
rect 8850 1700 9080 1710
rect 9320 1700 9330 1710
rect 1920 1690 2030 1700
rect 2480 1690 2570 1700
rect 2600 1690 2660 1700
rect 3120 1690 3220 1700
rect 4070 1690 4240 1700
rect 4480 1690 4490 1700
rect 4640 1690 4650 1700
rect 4750 1690 4760 1700
rect 4810 1690 4820 1700
rect 4830 1690 4840 1700
rect 4960 1690 4970 1700
rect 5240 1690 5250 1700
rect 5270 1690 5280 1700
rect 5350 1690 5360 1700
rect 5380 1690 5390 1700
rect 5420 1690 5430 1700
rect 5520 1690 5530 1700
rect 6850 1690 7020 1700
rect 7130 1690 7340 1700
rect 7870 1690 7950 1700
rect 8510 1690 8610 1700
rect 8850 1690 9080 1700
rect 9350 1690 9360 1700
rect 9790 1690 9800 1700
rect 1920 1680 2030 1690
rect 2480 1680 2540 1690
rect 2550 1680 2560 1690
rect 2590 1680 2660 1690
rect 3110 1680 3220 1690
rect 4080 1680 4250 1690
rect 4290 1680 4310 1690
rect 4480 1680 4490 1690
rect 4600 1680 4610 1690
rect 4660 1680 4670 1690
rect 4710 1680 4720 1690
rect 4820 1680 4830 1690
rect 4980 1680 4990 1690
rect 5100 1680 5110 1690
rect 5210 1680 5220 1690
rect 5340 1680 5350 1690
rect 5370 1680 5380 1690
rect 5410 1680 5420 1690
rect 5460 1680 5470 1690
rect 5480 1680 5490 1690
rect 6850 1680 7020 1690
rect 7130 1680 7340 1690
rect 7870 1680 7960 1690
rect 8510 1680 8620 1690
rect 8860 1680 9080 1690
rect 9110 1680 9120 1690
rect 9350 1680 9370 1690
rect 9700 1680 9710 1690
rect 9880 1680 9890 1690
rect 1930 1670 2040 1680
rect 2470 1670 2570 1680
rect 2580 1670 2590 1680
rect 2600 1670 2660 1680
rect 2710 1670 2720 1680
rect 3110 1670 3210 1680
rect 4080 1670 4170 1680
rect 4180 1670 4240 1680
rect 4300 1670 4310 1680
rect 4400 1670 4410 1680
rect 4440 1670 4450 1680
rect 4480 1670 4500 1680
rect 4690 1670 4700 1680
rect 4710 1670 4720 1680
rect 4760 1670 4770 1680
rect 5010 1670 5020 1680
rect 5230 1670 5240 1680
rect 5260 1670 5270 1680
rect 5430 1670 5440 1680
rect 5460 1670 5470 1680
rect 5550 1670 5560 1680
rect 6840 1670 7020 1680
rect 7140 1670 7350 1680
rect 7870 1670 7970 1680
rect 8330 1670 8340 1680
rect 8510 1670 8620 1680
rect 8840 1670 9080 1680
rect 9200 1670 9210 1680
rect 9530 1670 9550 1680
rect 1930 1660 2050 1670
rect 2450 1660 2720 1670
rect 3100 1660 3210 1670
rect 4080 1660 4160 1670
rect 4170 1660 4260 1670
rect 4300 1660 4310 1670
rect 4370 1660 4390 1670
rect 4490 1660 4500 1670
rect 4690 1660 4700 1670
rect 4730 1660 4740 1670
rect 4830 1660 4860 1670
rect 5200 1660 5210 1670
rect 5460 1660 5470 1670
rect 5550 1660 5560 1670
rect 6840 1660 7010 1670
rect 7140 1660 7350 1670
rect 7870 1660 7970 1670
rect 8520 1660 8630 1670
rect 8830 1660 9080 1670
rect 9530 1660 9540 1670
rect 9610 1660 9630 1670
rect 9670 1660 9690 1670
rect 9790 1660 9800 1670
rect 9960 1660 9970 1670
rect 1940 1650 2050 1660
rect 2420 1650 2740 1660
rect 3100 1650 3200 1660
rect 4100 1650 4130 1660
rect 4190 1650 4250 1660
rect 4350 1650 4370 1660
rect 4500 1650 4510 1660
rect 4520 1650 4530 1660
rect 4830 1650 4840 1660
rect 5020 1650 5030 1660
rect 5100 1650 5110 1660
rect 5190 1650 5200 1660
rect 5250 1650 5260 1660
rect 5300 1650 5320 1660
rect 6840 1650 7000 1660
rect 7140 1650 7350 1660
rect 7870 1650 7970 1660
rect 8510 1650 8630 1660
rect 8830 1650 9080 1660
rect 9620 1650 9630 1660
rect 9660 1650 9680 1660
rect 9950 1650 9960 1660
rect 1940 1640 2060 1650
rect 2420 1640 2730 1650
rect 3090 1640 3200 1650
rect 4090 1640 4100 1650
rect 4200 1640 4270 1650
rect 4480 1640 4490 1650
rect 4530 1640 4540 1650
rect 4860 1640 4870 1650
rect 5000 1640 5010 1650
rect 5100 1640 5110 1650
rect 5210 1640 5220 1650
rect 5300 1640 5310 1650
rect 5400 1640 5410 1650
rect 5430 1640 5440 1650
rect 5480 1640 5490 1650
rect 5520 1640 5530 1650
rect 5560 1640 5570 1650
rect 6830 1640 7000 1650
rect 7150 1640 7350 1650
rect 7870 1640 7980 1650
rect 8430 1640 8450 1650
rect 8480 1640 8490 1650
rect 8500 1640 8620 1650
rect 8630 1640 8650 1650
rect 8820 1640 9080 1650
rect 9220 1640 9230 1650
rect 9860 1640 9870 1650
rect 9890 1640 9900 1650
rect 9950 1640 9970 1650
rect 1940 1630 2070 1640
rect 2390 1630 2750 1640
rect 2760 1630 2770 1640
rect 3090 1630 3190 1640
rect 4210 1630 4270 1640
rect 4300 1630 4310 1640
rect 4420 1630 4430 1640
rect 4500 1630 4510 1640
rect 4520 1630 4530 1640
rect 4980 1630 4990 1640
rect 5170 1630 5180 1640
rect 5200 1630 5210 1640
rect 5470 1630 5480 1640
rect 5540 1630 5550 1640
rect 5560 1630 5570 1640
rect 6840 1630 7000 1640
rect 7150 1630 7350 1640
rect 7870 1630 7970 1640
rect 8320 1630 8330 1640
rect 8430 1630 8450 1640
rect 8470 1630 8620 1640
rect 8630 1630 8650 1640
rect 8820 1630 9080 1640
rect 9810 1630 9820 1640
rect 9840 1630 9860 1640
rect 1950 1620 2070 1630
rect 2370 1620 2750 1630
rect 2760 1620 2770 1630
rect 3070 1620 3190 1630
rect 4210 1620 4280 1630
rect 4300 1620 4310 1630
rect 4410 1620 4440 1630
rect 5100 1620 5110 1630
rect 5320 1620 5330 1630
rect 5420 1620 5430 1630
rect 5450 1620 5470 1630
rect 5560 1620 5570 1630
rect 5620 1620 5640 1630
rect 6840 1620 7000 1630
rect 7140 1620 7360 1630
rect 7880 1620 7970 1630
rect 8320 1620 8330 1630
rect 8430 1620 8640 1630
rect 8790 1620 8800 1630
rect 8810 1620 9070 1630
rect 9260 1620 9270 1630
rect 9710 1620 9720 1630
rect 9730 1620 9740 1630
rect 9800 1620 9820 1630
rect 9940 1620 9950 1630
rect 1950 1610 2080 1620
rect 2380 1610 2750 1620
rect 3060 1610 3170 1620
rect 4220 1610 4280 1620
rect 4300 1610 4310 1620
rect 4350 1610 4360 1620
rect 4380 1610 4390 1620
rect 5130 1610 5140 1620
rect 5250 1610 5260 1620
rect 5280 1610 5290 1620
rect 5310 1610 5320 1620
rect 5530 1610 5540 1620
rect 5600 1610 5620 1620
rect 5650 1610 5660 1620
rect 6830 1610 7000 1620
rect 7140 1610 7350 1620
rect 7880 1610 7960 1620
rect 8430 1610 8640 1620
rect 8660 1610 8700 1620
rect 8790 1610 9070 1620
rect 9220 1610 9230 1620
rect 9240 1610 9250 1620
rect 9370 1610 9380 1620
rect 9420 1610 9430 1620
rect 9700 1610 9710 1620
rect 9840 1610 9850 1620
rect 9940 1610 9950 1620
rect 1960 1600 2090 1610
rect 2370 1600 2730 1610
rect 3060 1600 3170 1610
rect 4220 1600 4280 1610
rect 4300 1600 4310 1610
rect 5210 1600 5220 1610
rect 5240 1600 5250 1610
rect 5400 1600 5410 1610
rect 5480 1600 5490 1610
rect 5540 1600 5550 1610
rect 5580 1600 5590 1610
rect 5670 1600 5680 1610
rect 6840 1600 7000 1610
rect 7140 1600 7360 1610
rect 7880 1600 7950 1610
rect 7960 1600 7970 1610
rect 8440 1600 8610 1610
rect 8630 1600 8640 1610
rect 8660 1600 8710 1610
rect 8780 1600 9070 1610
rect 9120 1600 9130 1610
rect 9420 1600 9430 1610
rect 9930 1600 9940 1610
rect 1970 1590 2100 1600
rect 2370 1590 2720 1600
rect 3050 1590 3160 1600
rect 4220 1590 4280 1600
rect 4310 1590 4320 1600
rect 5130 1590 5140 1600
rect 5230 1590 5240 1600
rect 5460 1590 5470 1600
rect 5640 1590 5660 1600
rect 6830 1590 7000 1600
rect 7010 1590 7030 1600
rect 7130 1590 7360 1600
rect 7880 1590 7950 1600
rect 7960 1590 7970 1600
rect 8450 1590 8600 1600
rect 8610 1590 8620 1600
rect 8660 1590 8740 1600
rect 8750 1590 8760 1600
rect 8770 1590 9070 1600
rect 9920 1590 9940 1600
rect 1970 1580 2110 1590
rect 2370 1580 2710 1590
rect 3030 1580 3150 1590
rect 4220 1580 4280 1590
rect 5210 1580 5220 1590
rect 5290 1580 5300 1590
rect 5400 1580 5410 1590
rect 5450 1580 5460 1590
rect 5520 1580 5540 1590
rect 5570 1580 5580 1590
rect 5590 1580 5600 1590
rect 5660 1580 5670 1590
rect 6840 1580 7030 1590
rect 7130 1580 7360 1590
rect 7880 1580 7970 1590
rect 8310 1580 8320 1590
rect 8450 1580 8620 1590
rect 8670 1580 9070 1590
rect 9310 1580 9330 1590
rect 9960 1580 9970 1590
rect 9980 1580 9990 1590
rect 1970 1570 2110 1580
rect 2370 1570 2700 1580
rect 3000 1570 3140 1580
rect 4230 1570 4280 1580
rect 5250 1570 5260 1580
rect 5330 1570 5340 1580
rect 5460 1570 5470 1580
rect 5510 1570 5520 1580
rect 5700 1570 5710 1580
rect 6840 1570 7000 1580
rect 7150 1570 7360 1580
rect 7880 1570 7970 1580
rect 8450 1570 8610 1580
rect 8660 1570 9070 1580
rect 9330 1570 9340 1580
rect 9910 1570 9920 1580
rect 9940 1570 9950 1580
rect 1980 1560 2140 1570
rect 2380 1560 2680 1570
rect 2990 1560 3140 1570
rect 4220 1560 4280 1570
rect 4960 1560 4970 1570
rect 5270 1560 5280 1570
rect 5380 1560 5390 1570
rect 5410 1560 5420 1570
rect 5490 1560 5520 1570
rect 5560 1560 5570 1570
rect 5580 1560 5590 1570
rect 5630 1560 5640 1570
rect 6830 1560 7000 1570
rect 7160 1560 7370 1570
rect 7890 1560 7990 1570
rect 8450 1560 8580 1570
rect 8600 1560 8620 1570
rect 8660 1560 9070 1570
rect 9720 1560 9730 1570
rect 9800 1560 9810 1570
rect 9850 1560 9860 1570
rect 1990 1550 2140 1560
rect 2440 1550 2520 1560
rect 2960 1550 3120 1560
rect 4120 1550 4130 1560
rect 4240 1550 4280 1560
rect 5260 1550 5280 1560
rect 5310 1550 5320 1560
rect 5370 1550 5380 1560
rect 5430 1550 5440 1560
rect 5450 1550 5460 1560
rect 5480 1550 5500 1560
rect 5560 1550 5570 1560
rect 5610 1550 5620 1560
rect 6840 1550 7000 1560
rect 7180 1550 7370 1560
rect 7890 1550 8000 1560
rect 8300 1550 8310 1560
rect 8460 1550 8590 1560
rect 8670 1550 9070 1560
rect 9800 1550 9810 1560
rect 9900 1550 9910 1560
rect 2000 1540 2160 1550
rect 2950 1540 3110 1550
rect 4240 1540 4270 1550
rect 4320 1540 4330 1550
rect 5270 1540 5280 1550
rect 5300 1540 5310 1550
rect 5320 1540 5330 1550
rect 5560 1540 5570 1550
rect 5700 1540 5710 1550
rect 6830 1540 6980 1550
rect 6990 1540 7000 1550
rect 7180 1540 7370 1550
rect 7880 1540 8000 1550
rect 8300 1540 8310 1550
rect 8440 1540 8580 1550
rect 8660 1540 9060 1550
rect 9580 1540 9600 1550
rect 9840 1540 9850 1550
rect 9900 1540 9920 1550
rect 2010 1530 2170 1540
rect 2940 1530 3100 1540
rect 4250 1530 4270 1540
rect 5720 1530 5730 1540
rect 6830 1530 6980 1540
rect 7170 1530 7370 1540
rect 7880 1530 8000 1540
rect 8450 1530 8620 1540
rect 8670 1530 9060 1540
rect 9470 1530 9490 1540
rect 9530 1530 9540 1540
rect 9890 1530 9910 1540
rect 2010 1520 2180 1530
rect 2930 1520 3090 1530
rect 4250 1520 4260 1530
rect 5310 1520 5320 1530
rect 5600 1520 5610 1530
rect 5720 1520 5730 1530
rect 6830 1520 6990 1530
rect 7170 1520 7190 1530
rect 7220 1520 7370 1530
rect 7880 1520 8010 1530
rect 8450 1520 8650 1530
rect 8670 1520 9000 1530
rect 9010 1520 9070 1530
rect 9890 1520 9910 1530
rect 9950 1520 9960 1530
rect 2020 1510 2190 1520
rect 2920 1510 3080 1520
rect 4140 1510 4150 1520
rect 4240 1510 4250 1520
rect 5600 1510 5610 1520
rect 5620 1510 5630 1520
rect 5700 1510 5710 1520
rect 6820 1510 6990 1520
rect 7210 1510 7370 1520
rect 7890 1510 8020 1520
rect 8290 1510 8300 1520
rect 8450 1510 8650 1520
rect 8670 1510 9000 1520
rect 9010 1510 9060 1520
rect 9180 1510 9210 1520
rect 9500 1510 9510 1520
rect 9700 1510 9710 1520
rect 9780 1510 9790 1520
rect 9880 1510 9890 1520
rect 9930 1510 9940 1520
rect 9960 1510 9970 1520
rect 2020 1500 2210 1510
rect 2920 1500 3070 1510
rect 4140 1500 4250 1510
rect 4340 1500 4350 1510
rect 5450 1500 5460 1510
rect 5600 1500 5610 1510
rect 5620 1500 5630 1510
rect 6820 1500 6980 1510
rect 7200 1500 7370 1510
rect 7880 1500 8020 1510
rect 8290 1500 8300 1510
rect 8450 1500 8640 1510
rect 8680 1500 9060 1510
rect 9230 1500 9240 1510
rect 9360 1500 9370 1510
rect 9410 1500 9430 1510
rect 9590 1500 9600 1510
rect 9820 1500 9830 1510
rect 9960 1500 9970 1510
rect 2040 1490 2210 1500
rect 2910 1490 3060 1500
rect 4140 1490 4250 1500
rect 5450 1490 5460 1500
rect 5500 1490 5510 1500
rect 5600 1490 5610 1500
rect 5620 1490 5630 1500
rect 6820 1490 6960 1500
rect 6970 1490 6980 1500
rect 7190 1490 7200 1500
rect 7220 1490 7370 1500
rect 7890 1490 8000 1500
rect 8450 1490 8640 1500
rect 8670 1490 8680 1500
rect 8690 1490 9070 1500
rect 9190 1490 9200 1500
rect 9230 1490 9240 1500
rect 9810 1490 9820 1500
rect 9890 1490 9900 1500
rect 9930 1490 9940 1500
rect 2040 1480 2220 1490
rect 2900 1480 2950 1490
rect 2960 1480 2980 1490
rect 3010 1480 3050 1490
rect 4150 1480 4260 1490
rect 5450 1480 5480 1490
rect 5490 1480 5510 1490
rect 5600 1480 5610 1490
rect 5620 1480 5630 1490
rect 5670 1480 5680 1490
rect 5690 1480 5700 1490
rect 6820 1480 6960 1490
rect 7230 1480 7240 1490
rect 7250 1480 7370 1490
rect 7890 1480 7990 1490
rect 8270 1480 8290 1490
rect 8450 1480 8610 1490
rect 8670 1480 8680 1490
rect 8720 1480 9070 1490
rect 9210 1480 9220 1490
rect 9230 1480 9240 1490
rect 9340 1480 9350 1490
rect 9570 1480 9580 1490
rect 9860 1480 9870 1490
rect 9890 1480 9900 1490
rect 2060 1470 2220 1480
rect 2890 1470 2940 1480
rect 3000 1470 3020 1480
rect 4140 1470 4260 1480
rect 4350 1470 4360 1480
rect 5450 1470 5460 1480
rect 5500 1470 5510 1480
rect 5600 1470 5610 1480
rect 5620 1470 5630 1480
rect 5680 1470 5690 1480
rect 5730 1470 5740 1480
rect 6810 1470 6960 1480
rect 7260 1470 7370 1480
rect 7900 1470 8000 1480
rect 8270 1470 8280 1480
rect 8450 1470 8590 1480
rect 8690 1470 8700 1480
rect 8720 1470 9070 1480
rect 9210 1470 9230 1480
rect 9590 1470 9600 1480
rect 9800 1470 9810 1480
rect 9860 1470 9880 1480
rect 2070 1460 2230 1470
rect 2880 1460 2920 1470
rect 4160 1460 4270 1470
rect 5570 1460 5580 1470
rect 5600 1460 5610 1470
rect 5620 1460 5630 1470
rect 6810 1460 6930 1470
rect 7250 1460 7370 1470
rect 7900 1460 8010 1470
rect 8270 1460 8280 1470
rect 8450 1460 8590 1470
rect 8750 1460 9070 1470
rect 9090 1460 9100 1470
rect 9520 1460 9530 1470
rect 9640 1460 9650 1470
rect 900 1450 940 1460
rect 2080 1450 2240 1460
rect 2870 1450 2910 1460
rect 4150 1450 4270 1460
rect 5460 1450 5470 1460
rect 5490 1450 5500 1460
rect 5550 1450 5560 1460
rect 5600 1450 5610 1460
rect 5620 1450 5630 1460
rect 5700 1450 5710 1460
rect 6810 1450 6930 1460
rect 7230 1450 7360 1460
rect 7370 1450 7380 1460
rect 7900 1450 8010 1460
rect 8260 1450 8280 1460
rect 8450 1450 8590 1460
rect 8700 1450 8710 1460
rect 8720 1450 9070 1460
rect 9080 1450 9110 1460
rect 9640 1450 9650 1460
rect 9950 1450 9960 1460
rect 880 1440 890 1450
rect 920 1440 930 1450
rect 940 1440 970 1450
rect 2080 1440 2240 1450
rect 2850 1440 2910 1450
rect 4150 1440 4280 1450
rect 5490 1440 5500 1450
rect 5600 1440 5610 1450
rect 5620 1440 5630 1450
rect 6810 1440 6920 1450
rect 7230 1440 7250 1450
rect 7260 1440 7380 1450
rect 7900 1440 8010 1450
rect 8260 1440 8280 1450
rect 8440 1440 8590 1450
rect 8620 1440 8630 1450
rect 8690 1440 9110 1450
rect 9340 1440 9350 1450
rect 9360 1440 9370 1450
rect 9390 1440 9410 1450
rect 9600 1440 9610 1450
rect 9780 1440 9790 1450
rect 9950 1440 9970 1450
rect 2100 1430 2250 1440
rect 2850 1430 2890 1440
rect 4160 1430 4290 1440
rect 5490 1430 5500 1440
rect 5600 1430 5610 1440
rect 6810 1430 6880 1440
rect 6900 1430 6910 1440
rect 7260 1430 7380 1440
rect 7890 1430 8010 1440
rect 8240 1430 8270 1440
rect 8440 1430 8580 1440
rect 8610 1430 8640 1440
rect 8700 1430 9070 1440
rect 9080 1430 9110 1440
rect 9350 1430 9360 1440
rect 9510 1430 9560 1440
rect 9580 1430 9590 1440
rect 9840 1430 9850 1440
rect 860 1420 870 1430
rect 2120 1420 2260 1430
rect 2840 1420 2890 1430
rect 4170 1420 4290 1430
rect 5470 1420 5480 1430
rect 5490 1420 5500 1430
rect 5520 1420 5540 1430
rect 5560 1420 5570 1430
rect 6810 1420 6860 1430
rect 7270 1420 7370 1430
rect 7910 1420 8010 1430
rect 8230 1420 8270 1430
rect 8440 1420 8590 1430
rect 8610 1420 8680 1430
rect 8690 1420 9070 1430
rect 9080 1420 9110 1430
rect 9350 1420 9370 1430
rect 9490 1420 9500 1430
rect 9550 1420 9560 1430
rect 9580 1420 9590 1430
rect 9610 1420 9620 1430
rect 9730 1420 9740 1430
rect 9830 1420 9840 1430
rect 2120 1410 2270 1420
rect 2830 1410 2870 1420
rect 4170 1410 4290 1420
rect 5450 1410 5460 1420
rect 5500 1410 5510 1420
rect 5550 1410 5560 1420
rect 5590 1410 5600 1420
rect 5610 1410 5620 1420
rect 6810 1410 6860 1420
rect 7270 1410 7370 1420
rect 7910 1410 7990 1420
rect 8060 1410 8070 1420
rect 8220 1410 8270 1420
rect 8460 1410 8600 1420
rect 8620 1410 9110 1420
rect 9240 1410 9250 1420
rect 9410 1410 9420 1420
rect 9500 1410 9510 1420
rect 9530 1410 9540 1420
rect 9640 1410 9650 1420
rect 9690 1410 9700 1420
rect 9930 1410 9950 1420
rect 9970 1410 9990 1420
rect 2130 1400 2290 1410
rect 2820 1400 2870 1410
rect 4170 1400 4310 1410
rect 5520 1400 5540 1410
rect 6810 1400 6860 1410
rect 7270 1400 7380 1410
rect 7910 1400 7990 1410
rect 8040 1400 8050 1410
rect 8210 1400 8260 1410
rect 8440 1400 8460 1410
rect 8470 1400 9110 1410
rect 9290 1400 9310 1410
rect 9590 1400 9600 1410
rect 9620 1400 9640 1410
rect 9870 1400 9880 1410
rect 9940 1400 9950 1410
rect 9960 1400 9990 1410
rect 2150 1390 2300 1400
rect 2810 1390 2860 1400
rect 4170 1390 4320 1400
rect 5460 1390 5470 1400
rect 5580 1390 5590 1400
rect 6820 1390 6850 1400
rect 7260 1390 7380 1400
rect 7910 1390 8010 1400
rect 8170 1390 8180 1400
rect 8200 1390 8260 1400
rect 8440 1390 9110 1400
rect 9260 1390 9270 1400
rect 9280 1390 9290 1400
rect 9300 1390 9310 1400
rect 9590 1390 9600 1400
rect 9620 1390 9640 1400
rect 9810 1390 9830 1400
rect 9860 1390 9870 1400
rect 9940 1390 9950 1400
rect 9990 1390 9990 1400
rect 2160 1380 2310 1390
rect 2800 1380 2850 1390
rect 4170 1380 4330 1390
rect 5570 1380 5580 1390
rect 6820 1380 6850 1390
rect 7270 1380 7390 1390
rect 7910 1380 8010 1390
rect 8190 1380 8250 1390
rect 8460 1380 9110 1390
rect 9210 1380 9220 1390
rect 9540 1380 9550 1390
rect 9620 1380 9650 1390
rect 9810 1380 9830 1390
rect 9920 1380 9930 1390
rect 2170 1370 2320 1380
rect 2780 1370 2840 1380
rect 4180 1370 4210 1380
rect 4240 1370 4330 1380
rect 5500 1370 5510 1380
rect 5560 1370 5570 1380
rect 5590 1370 5600 1380
rect 6820 1370 6860 1380
rect 7270 1370 7380 1380
rect 7920 1370 8010 1380
rect 8170 1370 8240 1380
rect 8460 1370 9110 1380
rect 9200 1370 9210 1380
rect 9280 1370 9290 1380
rect 9520 1370 9550 1380
rect 9570 1370 9610 1380
rect 9800 1370 9810 1380
rect 9820 1370 9830 1380
rect 9870 1370 9920 1380
rect 9930 1370 9950 1380
rect 2180 1360 2340 1370
rect 2770 1360 2820 1370
rect 4180 1360 4200 1370
rect 4260 1360 4340 1370
rect 5580 1360 5590 1370
rect 6820 1360 6850 1370
rect 7260 1360 7390 1370
rect 7920 1360 8010 1370
rect 8160 1360 8230 1370
rect 8440 1360 9110 1370
rect 9260 1360 9270 1370
rect 9310 1360 9330 1370
rect 9460 1360 9470 1370
rect 9590 1360 9620 1370
rect 9820 1360 9830 1370
rect 9900 1360 9920 1370
rect 9960 1360 9970 1370
rect 2190 1350 2370 1360
rect 2760 1350 2820 1360
rect 3600 1350 3610 1360
rect 4190 1350 4200 1360
rect 4260 1350 4340 1360
rect 5490 1350 5500 1360
rect 6820 1350 6850 1360
rect 7260 1350 7380 1360
rect 7920 1350 8020 1360
rect 8150 1350 8210 1360
rect 8440 1350 9120 1360
rect 9260 1350 9270 1360
rect 9590 1350 9610 1360
rect 9690 1350 9700 1360
rect 9790 1350 9800 1360
rect 2220 1340 2240 1350
rect 2250 1340 2390 1350
rect 2730 1340 2800 1350
rect 4190 1340 4200 1350
rect 4270 1340 4340 1350
rect 6820 1340 6850 1350
rect 7270 1340 7280 1350
rect 7290 1340 7380 1350
rect 7920 1340 8040 1350
rect 8130 1340 8200 1350
rect 8430 1340 9120 1350
rect 9600 1340 9620 1350
rect 9640 1340 9650 1350
rect 9670 1340 9680 1350
rect 9950 1340 9960 1350
rect 2220 1330 2410 1340
rect 2720 1330 2790 1340
rect 4190 1330 4220 1340
rect 4270 1330 4330 1340
rect 4400 1330 4410 1340
rect 6820 1330 6850 1340
rect 7290 1330 7380 1340
rect 7910 1330 8050 1340
rect 8110 1330 8190 1340
rect 8440 1330 9120 1340
rect 9480 1330 9490 1340
rect 9620 1330 9630 1340
rect 9720 1330 9730 1340
rect 9770 1330 9780 1340
rect 9960 1330 9990 1340
rect 2230 1320 2290 1330
rect 2300 1320 2440 1330
rect 2700 1320 2770 1330
rect 3520 1320 3530 1330
rect 3650 1320 3660 1330
rect 4190 1320 4290 1330
rect 6820 1320 6850 1330
rect 7300 1320 7380 1330
rect 7920 1320 8010 1330
rect 8030 1320 8060 1330
rect 8080 1320 8190 1330
rect 8440 1320 9090 1330
rect 9100 1320 9120 1330
rect 9390 1320 9400 1330
rect 9450 1320 9470 1330
rect 2260 1310 2280 1320
rect 2340 1310 2530 1320
rect 2660 1310 2750 1320
rect 4200 1310 4290 1320
rect 6820 1310 6850 1320
rect 7280 1310 7290 1320
rect 7310 1310 7380 1320
rect 7920 1310 8020 1320
rect 8030 1310 8180 1320
rect 8420 1310 8440 1320
rect 8460 1310 9080 1320
rect 9100 1310 9120 1320
rect 9660 1310 9680 1320
rect 9920 1310 9940 1320
rect 2270 1300 2280 1310
rect 2360 1300 2720 1310
rect 4200 1300 4290 1310
rect 6830 1300 6850 1310
rect 7310 1300 7380 1310
rect 7920 1300 8180 1310
rect 8420 1300 8430 1310
rect 8440 1300 9080 1310
rect 9840 1300 9850 1310
rect 9980 1300 9990 1310
rect 2400 1290 2710 1300
rect 4200 1290 4250 1300
rect 4260 1290 4290 1300
rect 6820 1290 6850 1300
rect 7290 1290 7300 1300
rect 7310 1290 7380 1300
rect 7920 1290 8170 1300
rect 8430 1290 9080 1300
rect 9130 1290 9140 1300
rect 9590 1290 9600 1300
rect 9610 1290 9620 1300
rect 9830 1290 9860 1300
rect 2430 1280 2680 1290
rect 3700 1280 3710 1290
rect 4200 1280 4240 1290
rect 4270 1280 4290 1290
rect 5690 1280 5700 1290
rect 6820 1280 6850 1290
rect 7290 1280 7380 1290
rect 7920 1280 8180 1290
rect 8440 1280 9080 1290
rect 9120 1280 9130 1290
rect 9480 1280 9500 1290
rect 9830 1280 9840 1290
rect 9950 1280 9960 1290
rect 2440 1270 2490 1280
rect 2500 1270 2660 1280
rect 4200 1270 4210 1280
rect 4420 1270 4430 1280
rect 5690 1270 5700 1280
rect 6820 1270 6850 1280
rect 7300 1270 7380 1280
rect 7920 1270 8170 1280
rect 8450 1270 8990 1280
rect 9000 1270 9070 1280
rect 9460 1270 9470 1280
rect 9490 1270 9500 1280
rect 9690 1270 9700 1280
rect 9890 1270 9910 1280
rect 4200 1260 4210 1270
rect 5340 1260 5350 1270
rect 5440 1260 5450 1270
rect 6820 1260 6850 1270
rect 7290 1260 7380 1270
rect 7920 1260 8180 1270
rect 8450 1260 9070 1270
rect 9310 1260 9330 1270
rect 9400 1260 9450 1270
rect 9880 1260 9900 1270
rect 9940 1260 9950 1270
rect 3510 1250 3610 1260
rect 3620 1250 3650 1260
rect 5240 1250 5250 1260
rect 5270 1250 5280 1260
rect 5290 1250 5330 1260
rect 5390 1250 5410 1260
rect 5420 1250 5450 1260
rect 5670 1250 5680 1260
rect 6820 1250 6850 1260
rect 7300 1250 7380 1260
rect 7940 1250 8180 1260
rect 8460 1250 8980 1260
rect 8990 1250 9010 1260
rect 9020 1250 9070 1260
rect 9130 1250 9140 1260
rect 9590 1250 9610 1260
rect 9630 1250 9640 1260
rect 9730 1250 9740 1260
rect 3510 1240 3670 1250
rect 5150 1240 5160 1250
rect 5190 1240 5200 1250
rect 5290 1240 5300 1250
rect 5310 1240 5320 1250
rect 5380 1240 5400 1250
rect 5420 1240 5440 1250
rect 6830 1240 6850 1250
rect 7300 1240 7380 1250
rect 7400 1240 7410 1250
rect 7940 1240 8180 1250
rect 8460 1240 8900 1250
rect 8910 1240 8940 1250
rect 9000 1240 9010 1250
rect 9020 1240 9070 1250
rect 9290 1240 9320 1250
rect 9610 1240 9630 1250
rect 9720 1240 9730 1250
rect 9910 1240 9940 1250
rect 3520 1230 3540 1240
rect 3590 1230 3680 1240
rect 3760 1230 3770 1240
rect 4430 1230 4440 1240
rect 5060 1230 5070 1240
rect 5140 1230 5160 1240
rect 5180 1230 5190 1240
rect 5250 1230 5260 1240
rect 5280 1230 5290 1240
rect 5300 1230 5320 1240
rect 5330 1230 5340 1240
rect 5380 1230 5390 1240
rect 5400 1230 5410 1240
rect 5430 1230 5450 1240
rect 6830 1230 6860 1240
rect 7300 1230 7390 1240
rect 7950 1230 8180 1240
rect 8400 1230 8410 1240
rect 8450 1230 8940 1240
rect 9020 1230 9030 1240
rect 9040 1230 9070 1240
rect 9130 1230 9140 1240
rect 9490 1230 9500 1240
rect 9510 1230 9520 1240
rect 9620 1230 9630 1240
rect 9900 1230 9960 1240
rect 3520 1220 3530 1230
rect 3660 1220 3690 1230
rect 3780 1220 3790 1230
rect 5030 1220 5050 1230
rect 5070 1220 5080 1230
rect 5110 1220 5130 1230
rect 5140 1220 5150 1230
rect 5180 1220 5190 1230
rect 5200 1220 5210 1230
rect 5220 1220 5230 1230
rect 5320 1220 5330 1230
rect 5350 1220 5360 1230
rect 5370 1220 5380 1230
rect 5400 1220 5410 1230
rect 5440 1220 5460 1230
rect 6760 1220 6770 1230
rect 6830 1220 6850 1230
rect 7300 1220 7390 1230
rect 7950 1220 8180 1230
rect 8400 1220 8410 1230
rect 8450 1220 8880 1230
rect 8900 1220 8920 1230
rect 8970 1220 8980 1230
rect 9010 1220 9060 1230
rect 9110 1220 9120 1230
rect 9130 1220 9140 1230
rect 9490 1220 9500 1230
rect 9610 1220 9620 1230
rect 9950 1220 9960 1230
rect 3530 1210 3540 1220
rect 3660 1210 3700 1220
rect 4990 1210 5000 1220
rect 5020 1210 5040 1220
rect 5060 1210 5070 1220
rect 5100 1210 5130 1220
rect 5140 1210 5150 1220
rect 5210 1210 5230 1220
rect 5240 1210 5250 1220
rect 5270 1210 5280 1220
rect 5310 1210 5330 1220
rect 5350 1210 5400 1220
rect 5410 1210 5420 1220
rect 5450 1210 5460 1220
rect 6740 1210 6790 1220
rect 6830 1210 6860 1220
rect 7300 1210 7380 1220
rect 7950 1210 8180 1220
rect 8410 1210 8430 1220
rect 8440 1210 8900 1220
rect 8950 1210 8980 1220
rect 9000 1210 9070 1220
rect 9110 1210 9120 1220
rect 9310 1210 9320 1220
rect 9880 1210 9910 1220
rect 3670 1200 3720 1210
rect 3810 1200 3820 1210
rect 4210 1200 4220 1210
rect 4870 1200 4890 1210
rect 4990 1200 5000 1210
rect 5020 1200 5030 1210
rect 5070 1200 5080 1210
rect 5110 1200 5130 1210
rect 5140 1200 5160 1210
rect 5180 1200 5200 1210
rect 5210 1200 5250 1210
rect 5260 1200 5290 1210
rect 5300 1200 5310 1210
rect 5320 1200 5370 1210
rect 5400 1200 5420 1210
rect 5440 1200 5450 1210
rect 6730 1200 6790 1210
rect 6830 1200 6860 1210
rect 7300 1200 7380 1210
rect 7950 1200 8180 1210
rect 8380 1200 8860 1210
rect 8950 1200 8970 1210
rect 8990 1200 9000 1210
rect 9020 1200 9040 1210
rect 9060 1200 9070 1210
rect 9110 1200 9120 1210
rect 9310 1200 9320 1210
rect 9530 1200 9540 1210
rect 9570 1200 9590 1210
rect 9600 1200 9620 1210
rect 9650 1200 9660 1210
rect 9850 1200 9860 1210
rect 9890 1200 9910 1210
rect 9920 1200 9930 1210
rect 9940 1200 9950 1210
rect 3540 1190 3550 1200
rect 3680 1190 3730 1200
rect 4210 1190 4220 1200
rect 4770 1190 4780 1200
rect 4800 1190 4810 1200
rect 4830 1190 4840 1200
rect 4850 1190 4870 1200
rect 4880 1190 4900 1200
rect 5010 1190 5050 1200
rect 5060 1190 5070 1200
rect 5120 1190 5130 1200
rect 5140 1190 5150 1200
rect 5180 1190 5210 1200
rect 5220 1190 5230 1200
rect 6720 1190 6790 1200
rect 6830 1190 6850 1200
rect 7300 1190 7380 1200
rect 7950 1190 8180 1200
rect 8400 1190 8420 1200
rect 8430 1190 8500 1200
rect 8520 1190 8810 1200
rect 8850 1190 8860 1200
rect 8960 1190 8980 1200
rect 8990 1190 9040 1200
rect 9110 1190 9120 1200
rect 9280 1190 9300 1200
rect 9320 1190 9330 1200
rect 9500 1190 9510 1200
rect 9820 1190 9830 1200
rect 9840 1190 9850 1200
rect 3550 1180 3560 1190
rect 3700 1180 3750 1190
rect 4730 1180 4770 1190
rect 4810 1180 4840 1190
rect 4850 1180 4860 1190
rect 4870 1180 4890 1190
rect 5030 1180 5050 1190
rect 5070 1180 5080 1190
rect 5120 1180 5130 1190
rect 6710 1180 6790 1190
rect 6830 1180 6860 1190
rect 7300 1180 7380 1190
rect 7950 1180 8180 1190
rect 8380 1180 8410 1190
rect 8430 1180 8470 1190
rect 8480 1180 8550 1190
rect 8570 1180 8750 1190
rect 8770 1180 8810 1190
rect 9000 1180 9020 1190
rect 9110 1180 9120 1190
rect 9140 1180 9150 1190
rect 9360 1180 9380 1190
rect 9600 1180 9610 1190
rect 790 1170 810 1180
rect 3560 1170 3570 1180
rect 3720 1170 3750 1180
rect 4600 1170 4620 1180
rect 4640 1170 4650 1180
rect 4680 1170 4690 1180
rect 4700 1170 4710 1180
rect 4730 1170 4740 1180
rect 4770 1170 4780 1180
rect 4800 1170 4810 1180
rect 4850 1170 4860 1180
rect 4880 1170 4900 1180
rect 5000 1170 5010 1180
rect 5040 1170 5050 1180
rect 5070 1170 5080 1180
rect 6690 1170 6750 1180
rect 6760 1170 6790 1180
rect 6830 1170 6860 1180
rect 7300 1170 7380 1180
rect 7960 1170 8180 1180
rect 8370 1170 8410 1180
rect 8450 1170 8750 1180
rect 8790 1170 8800 1180
rect 9110 1170 9120 1180
rect 9540 1170 9550 1180
rect 790 1160 820 1170
rect 3570 1160 3580 1170
rect 3730 1160 3750 1170
rect 4450 1160 4460 1170
rect 4570 1160 4580 1170
rect 4600 1160 4610 1170
rect 4670 1160 4680 1170
rect 4700 1160 4720 1170
rect 4730 1160 4740 1170
rect 4780 1160 4790 1170
rect 4800 1160 4810 1170
rect 4820 1160 4840 1170
rect 4850 1160 4860 1170
rect 4890 1160 4900 1170
rect 4990 1160 5000 1170
rect 6670 1160 6710 1170
rect 6750 1160 6800 1170
rect 6830 1160 6860 1170
rect 7300 1160 7380 1170
rect 7960 1160 8170 1170
rect 8380 1160 8410 1170
rect 8430 1160 8520 1170
rect 8530 1160 8540 1170
rect 8550 1160 8730 1170
rect 8770 1160 8790 1170
rect 9110 1160 9120 1170
rect 9140 1160 9150 1170
rect 9590 1160 9600 1170
rect 9630 1160 9640 1170
rect 9680 1160 9700 1170
rect 9840 1160 9870 1170
rect 780 1150 830 1160
rect 3740 1150 3760 1160
rect 3880 1150 3890 1160
rect 4220 1150 4230 1160
rect 4450 1150 4460 1160
rect 4600 1150 4610 1160
rect 4670 1150 4680 1160
rect 4700 1150 4720 1160
rect 4730 1150 4740 1160
rect 4770 1150 4780 1160
rect 4800 1150 4810 1160
rect 4820 1150 4830 1160
rect 4840 1150 4860 1160
rect 4870 1150 4880 1160
rect 4890 1150 4900 1160
rect 6660 1150 6690 1160
rect 6770 1150 6790 1160
rect 6830 1150 6860 1160
rect 7300 1150 7380 1160
rect 7950 1150 8090 1160
rect 8100 1150 8170 1160
rect 8380 1150 8400 1160
rect 8430 1150 8720 1160
rect 8750 1150 8780 1160
rect 9110 1150 9120 1160
rect 9550 1150 9560 1160
rect 9850 1150 9860 1160
rect 780 1140 830 1150
rect 3740 1140 3750 1150
rect 4220 1140 4230 1150
rect 4600 1140 4620 1150
rect 4640 1140 4650 1150
rect 4670 1140 4680 1150
rect 4710 1140 4720 1150
rect 4730 1140 4740 1150
rect 4750 1140 4760 1150
rect 4780 1140 4790 1150
rect 4810 1140 4830 1150
rect 4840 1140 4860 1150
rect 4880 1140 4890 1150
rect 6640 1140 6670 1150
rect 6780 1140 6800 1150
rect 6830 1140 6850 1150
rect 7310 1140 7380 1150
rect 7950 1140 8090 1150
rect 8100 1140 8170 1150
rect 8380 1140 8510 1150
rect 8520 1140 8710 1150
rect 8760 1140 8770 1150
rect 9110 1140 9120 1150
rect 9520 1140 9530 1150
rect 9550 1140 9560 1150
rect 9710 1140 9720 1150
rect 9830 1140 9840 1150
rect 9850 1140 9860 1150
rect 9890 1140 9920 1150
rect 9930 1140 9940 1150
rect 9980 1140 9990 1150
rect 770 1130 830 1140
rect 3740 1130 3750 1140
rect 4220 1130 4240 1140
rect 4600 1130 4610 1140
rect 4620 1130 4630 1140
rect 4640 1130 4650 1140
rect 4670 1130 4680 1140
rect 4700 1130 4710 1140
rect 4720 1130 4730 1140
rect 4740 1130 4760 1140
rect 4770 1130 4790 1140
rect 6630 1130 6650 1140
rect 6770 1130 6800 1140
rect 6830 1130 6860 1140
rect 7310 1130 7380 1140
rect 7960 1130 8070 1140
rect 8100 1130 8170 1140
rect 8380 1130 8680 1140
rect 9110 1130 9120 1140
rect 9710 1130 9720 1140
rect 9820 1130 9830 1140
rect 9880 1130 9890 1140
rect 770 1120 830 1130
rect 3730 1120 3760 1130
rect 3920 1120 3930 1130
rect 4230 1120 4240 1130
rect 4570 1120 4590 1130
rect 4600 1120 4610 1130
rect 4620 1120 4630 1130
rect 6610 1120 6630 1130
rect 6780 1120 6800 1130
rect 6840 1120 6860 1130
rect 7310 1120 7380 1130
rect 7960 1120 8070 1130
rect 8100 1120 8170 1130
rect 8360 1120 8410 1130
rect 8420 1120 8460 1130
rect 8480 1120 8550 1130
rect 8560 1120 8570 1130
rect 8580 1120 8600 1130
rect 8630 1120 8680 1130
rect 9110 1120 9120 1130
rect 9550 1120 9560 1130
rect 9870 1120 9880 1130
rect 770 1110 830 1120
rect 3720 1110 3770 1120
rect 4460 1110 4470 1120
rect 4570 1110 4580 1120
rect 6590 1110 6620 1120
rect 6780 1110 6800 1120
rect 6840 1110 6860 1120
rect 7300 1110 7380 1120
rect 7960 1110 8060 1120
rect 8090 1110 8160 1120
rect 8350 1110 8460 1120
rect 8470 1110 8480 1120
rect 8490 1110 8540 1120
rect 8550 1110 8680 1120
rect 9110 1110 9120 1120
rect 9350 1110 9360 1120
rect 9550 1110 9570 1120
rect 9820 1110 9840 1120
rect 9870 1110 9880 1120
rect 9900 1110 9910 1120
rect 9990 1110 9990 1120
rect 760 1100 830 1110
rect 3630 1100 3640 1110
rect 3710 1100 3780 1110
rect 3950 1100 3960 1110
rect 6570 1100 6610 1110
rect 6780 1100 6800 1110
rect 6840 1100 6860 1110
rect 7300 1100 7390 1110
rect 7950 1100 8060 1110
rect 8090 1100 8160 1110
rect 8350 1100 8360 1110
rect 8370 1100 8420 1110
rect 8440 1100 8480 1110
rect 8490 1100 8620 1110
rect 8630 1100 8670 1110
rect 9110 1100 9120 1110
rect 9400 1100 9410 1110
rect 9550 1100 9560 1110
rect 9600 1100 9610 1110
rect 9650 1100 9670 1110
rect 9860 1100 9870 1110
rect 9990 1100 9990 1110
rect 760 1090 830 1100
rect 1550 1090 1620 1100
rect 3710 1090 3840 1100
rect 6560 1090 6580 1100
rect 6780 1090 6800 1100
rect 6830 1090 6850 1100
rect 7310 1090 7380 1100
rect 7960 1090 8070 1100
rect 8090 1090 8160 1100
rect 8350 1090 8410 1100
rect 8440 1090 8450 1100
rect 8460 1090 8550 1100
rect 8560 1090 8660 1100
rect 9110 1090 9120 1100
rect 9240 1090 9250 1100
rect 9270 1090 9280 1100
rect 9410 1090 9420 1100
rect 9540 1090 9550 1100
rect 9640 1090 9650 1100
rect 9850 1090 9870 1100
rect 9920 1090 9930 1100
rect 9940 1090 9950 1100
rect 760 1080 820 1090
rect 1530 1080 1630 1090
rect 3650 1080 3660 1090
rect 3700 1080 3850 1090
rect 3980 1080 3990 1090
rect 4470 1080 4480 1090
rect 6540 1080 6580 1090
rect 6780 1080 6800 1090
rect 6840 1080 6860 1090
rect 7310 1080 7380 1090
rect 7960 1080 8060 1090
rect 8090 1080 8160 1090
rect 8350 1080 8370 1090
rect 8390 1080 8400 1090
rect 8420 1080 8440 1090
rect 8460 1080 8550 1090
rect 8580 1080 8660 1090
rect 9110 1080 9120 1090
rect 9150 1080 9160 1090
rect 9180 1080 9190 1090
rect 9360 1080 9370 1090
rect 9580 1080 9590 1090
rect 9630 1080 9650 1090
rect 760 1070 820 1080
rect 1520 1070 1630 1080
rect 2160 1070 2180 1080
rect 3670 1070 3860 1080
rect 6520 1070 6580 1080
rect 6780 1070 6800 1080
rect 6840 1070 6860 1080
rect 7300 1070 7390 1080
rect 7960 1070 8070 1080
rect 8080 1070 8160 1080
rect 8360 1070 8370 1080
rect 8380 1070 8390 1080
rect 8400 1070 8410 1080
rect 8430 1070 8440 1080
rect 8460 1070 8500 1080
rect 8520 1070 8550 1080
rect 8570 1070 8590 1080
rect 8610 1070 8660 1080
rect 9110 1070 9140 1080
rect 9160 1070 9170 1080
rect 9360 1070 9370 1080
rect 9830 1070 9840 1080
rect 750 1060 810 1070
rect 1510 1060 1630 1070
rect 2090 1060 2100 1070
rect 2110 1060 2160 1070
rect 3680 1060 3770 1070
rect 3810 1060 3870 1070
rect 6500 1060 6560 1070
rect 6780 1060 6800 1070
rect 6840 1060 6860 1070
rect 7300 1060 7390 1070
rect 7960 1060 8060 1070
rect 8080 1060 8150 1070
rect 8390 1060 8400 1070
rect 8410 1060 8450 1070
rect 8470 1060 8560 1070
rect 8570 1060 8650 1070
rect 9100 1060 9140 1070
rect 9530 1060 9540 1070
rect 9880 1060 9890 1070
rect 9910 1060 9920 1070
rect 750 1050 810 1060
rect 1500 1050 1520 1060
rect 1530 1050 1600 1060
rect 2080 1050 2210 1060
rect 3690 1050 3760 1060
rect 3820 1050 3870 1060
rect 6480 1050 6560 1060
rect 6780 1050 6800 1060
rect 6840 1050 6850 1060
rect 7300 1050 7390 1060
rect 7960 1050 8050 1060
rect 8070 1050 8150 1060
rect 8320 1050 8330 1060
rect 8360 1050 8390 1060
rect 8400 1050 8440 1060
rect 8450 1050 8480 1060
rect 8490 1050 8560 1060
rect 8620 1050 8640 1060
rect 9110 1050 9120 1060
rect 9350 1050 9360 1060
rect 9620 1050 9630 1060
rect 9840 1050 9850 1060
rect 9890 1050 9900 1060
rect 9920 1050 9930 1060
rect 9940 1050 9950 1060
rect 9990 1050 9990 1060
rect 750 1040 810 1050
rect 1490 1040 1520 1050
rect 2070 1040 2220 1050
rect 3690 1040 3750 1050
rect 3840 1040 3870 1050
rect 4040 1040 4050 1050
rect 4550 1040 4560 1050
rect 6470 1040 6560 1050
rect 6780 1040 6800 1050
rect 6840 1040 6860 1050
rect 7320 1040 7390 1050
rect 7970 1040 8050 1050
rect 8070 1040 8150 1050
rect 8380 1040 8480 1050
rect 8490 1040 8500 1050
rect 8510 1040 8550 1050
rect 8640 1040 8650 1050
rect 9100 1040 9110 1050
rect 9240 1040 9250 1050
rect 9360 1040 9370 1050
rect 9560 1040 9570 1050
rect 9710 1040 9720 1050
rect 9850 1040 9870 1050
rect 9940 1040 9950 1050
rect 740 1030 810 1040
rect 1480 1030 1520 1040
rect 2060 1030 2210 1040
rect 3700 1030 3730 1040
rect 3850 1030 3870 1040
rect 4060 1030 4070 1040
rect 4220 1030 4230 1040
rect 4580 1030 4590 1040
rect 6450 1030 6550 1040
rect 6790 1030 6810 1040
rect 6840 1030 6870 1040
rect 7320 1030 7390 1040
rect 7970 1030 8050 1040
rect 8070 1030 8140 1040
rect 8370 1030 8480 1040
rect 8490 1030 8550 1040
rect 8630 1030 8650 1040
rect 9110 1030 9120 1040
rect 9330 1030 9340 1040
rect 9710 1030 9720 1040
rect 9910 1030 9920 1040
rect 9930 1030 9950 1040
rect 9980 1030 9990 1040
rect 740 1020 800 1030
rect 1470 1020 1510 1030
rect 2050 1020 2220 1030
rect 2250 1020 2260 1030
rect 3710 1020 3730 1030
rect 3850 1020 3870 1030
rect 4070 1020 4080 1030
rect 6450 1020 6540 1030
rect 6790 1020 6810 1030
rect 6840 1020 6860 1030
rect 7320 1020 7390 1030
rect 7970 1020 8050 1030
rect 8070 1020 8140 1030
rect 8350 1020 8480 1030
rect 8490 1020 8550 1030
rect 8630 1020 8650 1030
rect 9100 1020 9120 1030
rect 9240 1020 9260 1030
rect 9510 1020 9520 1030
rect 9550 1020 9560 1030
rect 9720 1020 9730 1030
rect 9850 1020 9870 1030
rect 9930 1020 9940 1030
rect 9960 1020 9970 1030
rect 740 1010 800 1020
rect 1450 1010 1490 1020
rect 2040 1010 2230 1020
rect 2240 1010 2280 1020
rect 3720 1010 3730 1020
rect 3840 1010 3870 1020
rect 4090 1010 4100 1020
rect 4650 1010 4660 1020
rect 6450 1010 6540 1020
rect 6790 1010 6810 1020
rect 6840 1010 6860 1020
rect 7310 1010 7390 1020
rect 7970 1010 8140 1020
rect 8350 1010 8520 1020
rect 8550 1010 8560 1020
rect 8590 1010 8650 1020
rect 9100 1010 9120 1020
rect 9220 1010 9250 1020
rect 730 1000 800 1010
rect 1450 1000 1490 1010
rect 2030 1000 2040 1010
rect 2050 1000 2290 1010
rect 3730 1000 3740 1010
rect 3830 1000 3870 1010
rect 4670 1000 4680 1010
rect 6460 1000 6540 1010
rect 6790 1000 6810 1010
rect 6840 1000 6860 1010
rect 7310 1000 7400 1010
rect 7970 1000 8140 1010
rect 8340 1000 8500 1010
rect 8530 1000 8540 1010
rect 8550 1000 8560 1010
rect 8600 1000 8660 1010
rect 9100 1000 9120 1010
rect 9220 1000 9240 1010
rect 9650 1000 9660 1010
rect 9920 1000 9930 1010
rect 730 990 790 1000
rect 1430 990 1480 1000
rect 2040 990 2300 1000
rect 2460 990 2480 1000
rect 2590 990 2620 1000
rect 2670 990 2730 1000
rect 3740 990 3750 1000
rect 3830 990 3890 1000
rect 4120 990 4130 1000
rect 6460 990 6540 1000
rect 6790 990 6810 1000
rect 6840 990 6870 1000
rect 7310 990 7400 1000
rect 7970 990 8140 1000
rect 8340 990 8360 1000
rect 8370 990 8570 1000
rect 9110 990 9120 1000
rect 9220 990 9260 1000
rect 9420 990 9430 1000
rect 9490 990 9500 1000
rect 9530 990 9540 1000
rect 9730 990 9740 1000
rect 9950 990 9970 1000
rect 720 980 790 990
rect 1420 980 1470 990
rect 2030 980 2300 990
rect 2340 980 2390 990
rect 2420 980 2530 990
rect 2560 980 2660 990
rect 2670 980 2740 990
rect 3740 980 3760 990
rect 3820 980 3890 990
rect 4140 980 4150 990
rect 4720 980 4730 990
rect 6460 980 6540 990
rect 6790 980 6810 990
rect 6840 980 6860 990
rect 7310 980 7400 990
rect 7970 980 8140 990
rect 8370 980 8560 990
rect 9110 980 9120 990
rect 9150 980 9160 990
rect 9220 980 9250 990
rect 9410 980 9420 990
rect 9530 980 9540 990
rect 9690 980 9700 990
rect 9730 980 9750 990
rect 9870 980 9900 990
rect 720 970 780 980
rect 1410 970 1460 980
rect 2040 970 2740 980
rect 3760 970 3780 980
rect 3830 970 3880 980
rect 4170 970 4190 980
rect 4740 970 4750 980
rect 6460 970 6540 980
rect 6790 970 6810 980
rect 6840 970 6860 980
rect 7310 970 7400 980
rect 7970 970 8130 980
rect 8370 970 8570 980
rect 9100 970 9120 980
rect 9480 970 9490 980
rect 9720 970 9730 980
rect 9780 970 9790 980
rect 9810 970 9820 980
rect 9870 970 9920 980
rect 9950 970 9960 980
rect 720 960 780 970
rect 1400 960 1460 970
rect 2030 960 2720 970
rect 3760 960 3800 970
rect 3830 960 3870 970
rect 5610 960 5620 970
rect 5640 960 5660 970
rect 5700 960 5720 970
rect 5730 960 5760 970
rect 5800 960 5810 970
rect 6470 960 6540 970
rect 6800 960 6820 970
rect 6840 960 6860 970
rect 7310 960 7390 970
rect 7970 960 8130 970
rect 8360 960 8560 970
rect 9110 960 9120 970
rect 9200 960 9220 970
rect 9770 960 9780 970
rect 9810 960 9820 970
rect 9830 960 9850 970
rect 710 950 780 960
rect 1390 950 1440 960
rect 2030 950 2730 960
rect 3780 950 3790 960
rect 3830 950 3870 960
rect 5380 950 5400 960
rect 5410 950 5420 960
rect 5430 950 5440 960
rect 5510 950 5530 960
rect 5550 950 5560 960
rect 5600 950 5630 960
rect 5640 950 5650 960
rect 5700 950 5710 960
rect 5730 950 5740 960
rect 5750 950 5760 960
rect 5770 950 5800 960
rect 6470 950 6540 960
rect 6800 950 6820 960
rect 6840 950 6860 960
rect 7310 950 7390 960
rect 7970 950 8130 960
rect 8370 950 8540 960
rect 8550 950 8570 960
rect 9110 950 9120 960
rect 9470 950 9480 960
rect 9850 950 9860 960
rect 710 940 780 950
rect 1370 940 1420 950
rect 2030 940 2730 950
rect 3790 940 3870 950
rect 5330 940 5350 950
rect 5380 940 5400 950
rect 5420 940 5450 950
rect 5470 940 5490 950
rect 5550 940 5570 950
rect 5600 940 5610 950
rect 5620 940 5630 950
rect 5650 940 5660 950
rect 5710 940 5720 950
rect 5730 940 5740 950
rect 5750 940 5760 950
rect 5770 940 5780 950
rect 5800 940 5810 950
rect 6470 940 6560 950
rect 6800 940 6820 950
rect 6840 940 6880 950
rect 7320 940 7390 950
rect 7980 940 8120 950
rect 8370 940 8570 950
rect 9110 940 9120 950
rect 9190 940 9200 950
rect 9210 940 9220 950
rect 9510 940 9520 950
rect 700 930 770 940
rect 1360 930 1410 940
rect 2030 930 2730 940
rect 3800 930 3870 940
rect 4810 930 4820 940
rect 5330 930 5350 940
rect 5410 930 5420 940
rect 5430 930 5450 940
rect 5460 930 5470 940
rect 5500 930 5510 940
rect 5530 930 5540 940
rect 5550 930 5560 940
rect 5640 930 5670 940
rect 5680 930 5690 940
rect 5710 930 5720 940
rect 5730 930 5740 940
rect 5750 930 5760 940
rect 5780 930 5790 940
rect 5800 930 5810 940
rect 6470 930 6550 940
rect 6810 930 6820 940
rect 6850 930 6880 940
rect 7320 930 7390 940
rect 7980 930 8130 940
rect 8370 930 8420 940
rect 8430 930 8580 940
rect 9110 930 9120 940
rect 9190 930 9210 940
rect 9500 930 9510 940
rect 9800 930 9810 940
rect 700 920 710 930
rect 720 920 780 930
rect 1350 920 1400 930
rect 2030 920 2730 930
rect 3810 920 3880 930
rect 4820 920 4830 930
rect 5330 920 5350 930
rect 5380 920 5390 930
rect 5410 920 5430 930
rect 5440 920 5450 930
rect 5460 920 5470 930
rect 5500 920 5510 930
rect 5540 920 5550 930
rect 5610 920 5630 930
rect 5660 920 5670 930
rect 5730 920 5740 930
rect 5750 920 5760 930
rect 5780 920 5790 930
rect 5800 920 5810 930
rect 6470 920 6560 930
rect 6810 920 6820 930
rect 6850 920 6880 930
rect 7310 920 7390 930
rect 7980 920 8130 930
rect 8380 920 8400 930
rect 8410 920 8420 930
rect 8430 920 8580 930
rect 8720 920 8740 930
rect 9110 920 9120 930
rect 9210 920 9240 930
rect 710 910 770 920
rect 1330 910 1390 920
rect 2030 910 2720 920
rect 3810 910 3890 920
rect 4630 910 4640 920
rect 5340 910 5350 920
rect 5390 910 5400 920
rect 5410 910 5430 920
rect 5440 910 5450 920
rect 5460 910 5490 920
rect 5500 910 5510 920
rect 5540 910 5560 920
rect 5610 910 5620 920
rect 5660 910 5670 920
rect 5710 910 5720 920
rect 5730 910 5760 920
rect 5780 910 5790 920
rect 6470 910 6560 920
rect 6810 910 6820 920
rect 6850 910 6890 920
rect 7320 910 7390 920
rect 7980 910 8130 920
rect 8400 910 8520 920
rect 8540 910 8590 920
rect 8710 910 8750 920
rect 9100 910 9110 920
rect 9490 910 9500 920
rect 9660 910 9670 920
rect 690 900 700 910
rect 710 900 770 910
rect 1320 900 1390 910
rect 2030 900 2710 910
rect 3830 900 3900 910
rect 3980 900 4040 910
rect 4620 900 4640 910
rect 5340 900 5350 910
rect 5370 900 5390 910
rect 5410 900 5430 910
rect 5440 900 5450 910
rect 5460 900 5470 910
rect 5500 900 5510 910
rect 5550 900 5560 910
rect 5570 900 5580 910
rect 5610 900 5620 910
rect 5640 900 5670 910
rect 5700 900 5720 910
rect 6470 900 6560 910
rect 6810 900 6830 910
rect 6850 900 6870 910
rect 7310 900 7380 910
rect 7980 900 8130 910
rect 8410 900 8430 910
rect 8440 900 8590 910
rect 8710 900 8720 910
rect 9100 900 9110 910
rect 9540 900 9550 910
rect 690 890 700 900
rect 710 890 770 900
rect 1310 890 1380 900
rect 2030 890 2710 900
rect 3840 890 3920 900
rect 3930 890 4050 900
rect 4620 890 4630 900
rect 5370 890 5380 900
rect 5410 890 5440 900
rect 5460 890 5470 900
rect 5480 890 5490 900
rect 5500 890 5520 900
rect 5550 890 5560 900
rect 5600 890 5610 900
rect 5620 890 5630 900
rect 5650 890 5660 900
rect 6470 890 6570 900
rect 6810 890 6830 900
rect 6850 890 6880 900
rect 7300 890 7380 900
rect 7990 890 8130 900
rect 8430 890 8610 900
rect 8700 890 8720 900
rect 9100 890 9110 900
rect 680 880 690 890
rect 700 880 770 890
rect 1300 880 1380 890
rect 2040 880 2700 890
rect 3850 880 4050 890
rect 4610 880 4620 890
rect 5350 880 5360 890
rect 5390 880 5400 890
rect 5410 880 5430 890
rect 5460 880 5470 890
rect 5480 880 5490 890
rect 5530 880 5540 890
rect 5610 880 5620 890
rect 6470 880 6570 890
rect 6810 880 6830 890
rect 6850 880 6880 890
rect 7290 880 7380 890
rect 7990 880 8130 890
rect 8430 880 8650 890
rect 8680 880 8720 890
rect 680 870 760 880
rect 1290 870 1370 880
rect 2040 870 2690 880
rect 3860 870 4050 880
rect 4570 870 4610 880
rect 5340 870 5350 880
rect 5380 870 5390 880
rect 5420 870 5430 880
rect 5440 870 5450 880
rect 5470 870 5480 880
rect 6480 870 6570 880
rect 6820 870 6830 880
rect 6860 870 6890 880
rect 7290 870 7380 880
rect 7990 870 8140 880
rect 8430 870 8640 880
rect 8680 870 8710 880
rect 9100 870 9110 880
rect 9470 870 9480 880
rect 9520 870 9530 880
rect 9550 870 9590 880
rect 690 860 760 870
rect 1270 860 1360 870
rect 2040 860 2680 870
rect 3870 860 4050 870
rect 4240 860 4260 870
rect 4560 860 4570 870
rect 4860 860 4870 870
rect 6470 860 6570 870
rect 6820 860 6840 870
rect 6860 860 6890 870
rect 7290 860 7380 870
rect 7990 860 8140 870
rect 8450 860 8640 870
rect 9180 860 9190 870
rect 9520 860 9530 870
rect 9550 860 9560 870
rect 9820 860 9830 870
rect 670 850 760 860
rect 1260 850 1340 860
rect 2050 850 2450 860
rect 2470 850 2530 860
rect 2540 850 2550 860
rect 2560 850 2660 860
rect 3870 850 4050 860
rect 4240 850 4270 860
rect 4560 850 4570 860
rect 6480 850 6570 860
rect 6830 850 6840 860
rect 6860 850 6890 860
rect 7290 850 7380 860
rect 7990 850 8140 860
rect 8460 850 8640 860
rect 9800 850 9830 860
rect 670 840 760 850
rect 1250 840 1330 850
rect 2040 840 2430 850
rect 2490 840 2520 850
rect 2570 840 2650 850
rect 3890 840 4050 850
rect 4250 840 4260 850
rect 4270 840 4280 850
rect 6480 840 6580 850
rect 6830 840 6840 850
rect 6860 840 6890 850
rect 7290 840 7370 850
rect 7990 840 8140 850
rect 8480 840 8520 850
rect 8530 840 8630 850
rect 9450 840 9460 850
rect 9780 840 9800 850
rect 9850 840 9890 850
rect 680 830 760 840
rect 1240 830 1330 840
rect 2040 830 2420 840
rect 2490 830 2540 840
rect 2580 830 2640 840
rect 3890 830 3970 840
rect 4010 830 4050 840
rect 4250 830 4260 840
rect 4280 830 4290 840
rect 4330 830 4340 840
rect 4570 830 4580 840
rect 6480 830 6580 840
rect 6830 830 6840 840
rect 6860 830 6890 840
rect 7290 830 7370 840
rect 7990 830 8140 840
rect 8480 830 8520 840
rect 8530 830 8630 840
rect 9190 830 9200 840
rect 9780 830 9800 840
rect 9850 830 9880 840
rect 690 820 760 830
rect 1220 820 1310 830
rect 2040 820 2370 830
rect 2380 820 2420 830
rect 2470 820 2480 830
rect 2500 820 2520 830
rect 2570 820 2620 830
rect 3910 820 3960 830
rect 4020 820 4050 830
rect 4290 820 4300 830
rect 4320 820 4340 830
rect 6500 820 6580 830
rect 6860 820 6890 830
rect 7280 820 7370 830
rect 7990 820 8140 830
rect 8540 820 8620 830
rect 9440 820 9450 830
rect 9830 820 9880 830
rect 9910 820 9920 830
rect 660 810 670 820
rect 680 810 760 820
rect 1210 810 1310 820
rect 2050 810 2370 820
rect 2390 810 2410 820
rect 2450 810 2460 820
rect 2470 810 2500 820
rect 2560 810 2600 820
rect 3910 810 3950 820
rect 4020 810 4040 820
rect 4270 810 4280 820
rect 4300 810 4340 820
rect 4890 810 4900 820
rect 6500 810 6580 820
rect 6860 810 6890 820
rect 7280 810 7370 820
rect 7990 810 8140 820
rect 8550 810 8620 820
rect 9290 810 9300 820
rect 9810 810 9820 820
rect 9850 810 9860 820
rect 9880 810 9910 820
rect 9920 810 9940 820
rect 670 800 750 810
rect 1190 800 1260 810
rect 2060 800 2390 810
rect 2430 800 2470 810
rect 2560 800 2580 810
rect 3930 800 3960 810
rect 4020 800 4040 810
rect 4280 800 4290 810
rect 4310 800 4350 810
rect 6500 800 6580 810
rect 6860 800 6890 810
rect 7280 800 7370 810
rect 8000 800 8130 810
rect 8610 800 8630 810
rect 9290 800 9320 810
rect 9880 800 9890 810
rect 9900 800 9910 810
rect 9930 800 9950 810
rect 650 790 660 800
rect 670 790 740 800
rect 1180 790 1240 800
rect 2060 790 2360 800
rect 2370 790 2380 800
rect 2420 790 2470 800
rect 2550 790 2560 800
rect 3940 790 3960 800
rect 4020 790 4030 800
rect 4290 790 4300 800
rect 4320 790 4350 800
rect 6510 790 6590 800
rect 6870 790 6890 800
rect 7280 790 7370 800
rect 8000 790 8140 800
rect 9290 790 9320 800
rect 9940 790 9950 800
rect 650 780 740 790
rect 1160 780 1240 790
rect 2070 780 2360 790
rect 2430 780 2470 790
rect 3960 780 3980 790
rect 4010 780 4030 790
rect 4300 780 4310 790
rect 4330 780 4350 790
rect 4900 780 4910 790
rect 6520 780 6590 790
rect 6870 780 6900 790
rect 7280 780 7360 790
rect 8000 780 8140 790
rect 9200 780 9210 790
rect 9300 780 9330 790
rect 650 770 660 780
rect 670 770 730 780
rect 1160 770 1240 780
rect 2070 770 2340 780
rect 2430 770 2460 780
rect 2520 770 2530 780
rect 3680 770 3700 780
rect 3980 770 3990 780
rect 4000 770 4030 780
rect 4310 770 4320 780
rect 6510 770 6520 780
rect 6530 770 6590 780
rect 6840 770 6850 780
rect 6870 770 6900 780
rect 7280 770 7360 780
rect 8000 770 8130 780
rect 9240 770 9250 780
rect 9410 770 9420 780
rect 9610 770 9620 780
rect 9840 770 9850 780
rect 670 760 720 770
rect 1140 760 1240 770
rect 2070 760 2320 770
rect 2330 760 2340 770
rect 2430 760 2460 770
rect 2500 760 2510 770
rect 3690 760 3710 770
rect 3760 760 3770 770
rect 3790 760 3800 770
rect 3810 760 3840 770
rect 3990 760 4030 770
rect 4320 760 4330 770
rect 6530 760 6590 770
rect 6840 760 6850 770
rect 6870 760 6900 770
rect 7280 760 7360 770
rect 8010 760 8140 770
rect 9240 760 9260 770
rect 9360 760 9370 770
rect 9460 760 9510 770
rect 9610 760 9630 770
rect 640 750 650 760
rect 660 750 720 760
rect 1130 750 1250 760
rect 2070 750 2310 760
rect 2440 750 2450 760
rect 2480 750 2490 760
rect 3570 750 3600 760
rect 3660 750 3710 760
rect 3870 750 3880 760
rect 4020 750 4040 760
rect 4330 750 4340 760
rect 4530 750 4540 760
rect 4800 750 4810 760
rect 6530 750 6590 760
rect 6840 750 6850 760
rect 6870 750 6900 760
rect 7280 750 7360 760
rect 8010 750 8130 760
rect 9240 750 9250 760
rect 9400 750 9410 760
rect 9480 750 9490 760
rect 9620 750 9630 760
rect 660 740 720 750
rect 1110 740 1240 750
rect 2080 740 2290 750
rect 2470 740 2480 750
rect 3530 740 3560 750
rect 3890 740 3900 750
rect 4000 740 4010 750
rect 4020 740 4060 750
rect 4340 740 4350 750
rect 4530 740 4540 750
rect 4790 740 4810 750
rect 6530 740 6600 750
rect 6840 740 6850 750
rect 6870 740 6900 750
rect 7280 740 7360 750
rect 8010 740 8130 750
rect 9220 740 9230 750
rect 9350 740 9360 750
rect 9390 740 9400 750
rect 9450 740 9480 750
rect 660 730 710 740
rect 1100 730 1220 740
rect 2080 730 2270 740
rect 2450 730 2460 740
rect 3510 730 3520 740
rect 3900 730 3910 740
rect 4010 730 4080 740
rect 4110 730 4130 740
rect 4140 730 4160 740
rect 4170 730 4180 740
rect 4520 730 4540 740
rect 4780 730 4810 740
rect 4910 730 4920 740
rect 6540 730 6600 740
rect 6840 730 6850 740
rect 6870 730 6910 740
rect 7270 730 7360 740
rect 8010 730 8130 740
rect 9120 730 9140 740
rect 9290 730 9310 740
rect 9450 730 9460 740
rect 9680 730 9690 740
rect 9720 730 9730 740
rect 630 720 640 730
rect 660 720 710 730
rect 1090 720 1220 730
rect 2090 720 2180 730
rect 2220 720 2240 730
rect 3420 720 3490 730
rect 4020 720 4220 730
rect 4770 720 4780 730
rect 4910 720 4920 730
rect 6540 720 6610 730
rect 6840 720 6850 730
rect 6880 720 6910 730
rect 7270 720 7360 730
rect 8020 720 8130 730
rect 9210 720 9300 730
rect 9670 720 9690 730
rect 650 710 700 720
rect 1090 710 1210 720
rect 2090 710 2190 720
rect 2200 710 2210 720
rect 2230 710 2240 720
rect 2390 710 2410 720
rect 3390 710 3410 720
rect 3920 710 3930 720
rect 4020 710 4230 720
rect 4730 710 4770 720
rect 4790 710 4820 720
rect 6550 710 6620 720
rect 6840 710 6850 720
rect 6880 710 6920 720
rect 7270 710 7350 720
rect 8020 710 8130 720
rect 9100 710 9110 720
rect 9220 710 9260 720
rect 9380 710 9390 720
rect 9510 710 9520 720
rect 9530 710 9560 720
rect 620 700 630 710
rect 650 700 700 710
rect 1080 700 1210 710
rect 2100 700 2200 710
rect 2380 700 2390 710
rect 2400 700 2410 710
rect 3380 700 3390 710
rect 4020 700 4160 710
rect 4170 700 4210 710
rect 4710 700 4750 710
rect 4790 700 4830 710
rect 4910 700 4920 710
rect 6550 700 6620 710
rect 6840 700 6860 710
rect 6880 700 6920 710
rect 7260 700 7350 710
rect 8020 700 8130 710
rect 9210 700 9220 710
rect 640 690 690 700
rect 1070 690 1210 700
rect 2100 690 2220 700
rect 2320 690 2330 700
rect 2360 690 2370 700
rect 2380 690 2390 700
rect 4040 690 4130 700
rect 4180 690 4200 700
rect 4800 690 4840 700
rect 4890 690 4920 700
rect 6560 690 6630 700
rect 6850 690 6860 700
rect 6880 690 6920 700
rect 7240 690 7350 700
rect 8020 690 8130 700
rect 9100 690 9110 700
rect 640 680 690 690
rect 1060 680 1210 690
rect 2110 680 2260 690
rect 2300 680 2330 690
rect 2350 680 2360 690
rect 3340 680 3350 690
rect 4050 680 4110 690
rect 4180 680 4190 690
rect 4810 680 4850 690
rect 4880 680 4920 690
rect 6560 680 6640 690
rect 6850 680 6860 690
rect 6880 680 6940 690
rect 7250 680 7340 690
rect 8030 680 8130 690
rect 9680 680 9690 690
rect 9700 680 9710 690
rect 610 670 690 680
rect 1060 670 1210 680
rect 2110 670 2250 680
rect 2300 670 2330 680
rect 2340 670 2360 680
rect 4050 670 4100 680
rect 4170 670 4180 680
rect 4810 670 4890 680
rect 6560 670 6640 680
rect 6850 670 6860 680
rect 6890 670 6940 680
rect 7240 670 7340 680
rect 8040 670 8130 680
rect 9310 670 9320 680
rect 9610 670 9630 680
rect 9680 670 9690 680
rect 9710 670 9720 680
rect 610 660 690 670
rect 1040 660 1210 670
rect 2120 660 2260 670
rect 2280 660 2290 670
rect 2300 660 2310 670
rect 2330 660 2340 670
rect 4060 660 4100 670
rect 4160 660 4170 670
rect 4820 660 4850 670
rect 4860 660 4870 670
rect 6570 660 6650 670
rect 6850 660 6860 670
rect 6890 660 6940 670
rect 7230 660 7340 670
rect 8040 660 8130 670
rect 9220 660 9230 670
rect 9630 660 9640 670
rect 9690 660 9700 670
rect 610 650 690 660
rect 1050 650 1200 660
rect 2120 650 2270 660
rect 2280 650 2320 660
rect 4070 650 4090 660
rect 4130 650 4160 660
rect 4560 650 4570 660
rect 4700 650 4710 660
rect 4850 650 4860 660
rect 4920 650 4930 660
rect 6580 650 6660 660
rect 6850 650 6860 660
rect 6890 650 6940 660
rect 7230 650 7340 660
rect 8050 650 8120 660
rect 9160 650 9220 660
rect 9340 650 9350 660
rect 9640 650 9650 660
rect 9680 650 9700 660
rect 650 640 670 650
rect 680 640 690 650
rect 1010 640 1030 650
rect 1050 640 1170 650
rect 2120 640 2310 650
rect 3280 640 3290 650
rect 4110 640 4130 650
rect 4560 640 4570 650
rect 4690 640 4710 650
rect 4840 640 4850 650
rect 6590 640 6660 650
rect 6850 640 6860 650
rect 6890 640 6950 650
rect 6960 640 6970 650
rect 7220 640 7330 650
rect 8060 640 8120 650
rect 9140 640 9180 650
rect 9640 640 9660 650
rect 9670 640 9690 650
rect 9720 640 9740 650
rect 9940 640 9960 650
rect 710 630 760 640
rect 980 630 1100 640
rect 2120 630 2290 640
rect 4080 630 4090 640
rect 4110 630 4120 640
rect 4550 630 4570 640
rect 4680 630 4710 640
rect 4820 630 4830 640
rect 6590 630 6680 640
rect 6860 630 6870 640
rect 6890 630 6960 640
rect 7210 630 7330 640
rect 8060 630 8120 640
rect 9150 630 9200 640
rect 9290 630 9300 640
rect 9330 630 9340 640
rect 9640 630 9690 640
rect 9910 630 9920 640
rect 9940 630 9960 640
rect 500 620 610 630
rect 700 620 770 630
rect 960 620 1090 630
rect 2130 620 2270 630
rect 3250 620 3260 630
rect 4050 620 4110 630
rect 4550 620 4560 630
rect 4670 620 4710 630
rect 4800 620 4820 630
rect 6590 620 6680 630
rect 6860 620 6870 630
rect 6900 620 6960 630
rect 7220 620 7320 630
rect 8070 620 8110 630
rect 9150 620 9200 630
rect 9210 620 9220 630
rect 9590 620 9610 630
rect 9620 620 9630 630
rect 9660 620 9690 630
rect 9940 620 9950 630
rect 470 610 630 620
rect 700 610 770 620
rect 930 610 940 620
rect 950 610 1060 620
rect 2140 610 2260 620
rect 3160 610 3170 620
rect 3210 610 3240 620
rect 4040 610 4050 620
rect 4670 610 4710 620
rect 4790 610 4800 620
rect 4930 610 4940 620
rect 6610 610 6690 620
rect 6860 610 6870 620
rect 6900 610 6970 620
rect 7220 610 7310 620
rect 8090 610 8110 620
rect 9150 610 9200 620
rect 9620 610 9660 620
rect 9670 610 9690 620
rect 9960 610 9990 620
rect 430 600 540 610
rect 560 600 630 610
rect 700 600 770 610
rect 930 600 1060 610
rect 2150 600 2240 610
rect 3140 600 3160 610
rect 3170 600 3220 610
rect 4040 600 4050 610
rect 4540 600 4550 610
rect 4560 600 4570 610
rect 4670 600 4710 610
rect 4780 600 4800 610
rect 6610 600 6700 610
rect 6860 600 6870 610
rect 6910 600 6980 610
rect 7210 600 7310 610
rect 8100 600 8110 610
rect 9160 600 9170 610
rect 9180 600 9200 610
rect 9230 600 9240 610
rect 9310 600 9320 610
rect 9690 600 9700 610
rect 410 590 460 600
rect 580 590 640 600
rect 710 590 770 600
rect 910 590 920 600
rect 930 590 1060 600
rect 2150 590 2210 600
rect 3130 590 3140 600
rect 4050 590 4060 600
rect 4080 590 4090 600
rect 4530 590 4540 600
rect 4560 590 4570 600
rect 4660 590 4710 600
rect 4770 590 4790 600
rect 6620 590 6710 600
rect 6870 590 6880 600
rect 6910 590 6990 600
rect 7200 590 7300 600
rect 9110 590 9120 600
rect 9140 590 9220 600
rect 9230 590 9240 600
rect 9670 590 9680 600
rect 9700 590 9730 600
rect 9910 590 9930 600
rect 9980 590 9990 600
rect 380 580 430 590
rect 600 580 650 590
rect 720 580 730 590
rect 740 580 750 590
rect 910 580 1050 590
rect 1400 580 1420 590
rect 2160 580 2180 590
rect 3120 580 3130 590
rect 4060 580 4070 590
rect 4080 580 4090 590
rect 4510 580 4530 590
rect 4560 580 4570 590
rect 4660 580 4690 590
rect 4770 580 4790 590
rect 4880 580 4890 590
rect 6640 580 6710 590
rect 6870 580 6880 590
rect 6910 580 6990 590
rect 7180 580 7190 590
rect 7200 580 7300 590
rect 9090 580 9100 590
rect 9120 580 9130 590
rect 9200 580 9220 590
rect 9300 580 9310 590
rect 9620 580 9640 590
rect 9670 580 9700 590
rect 360 570 390 580
rect 590 570 650 580
rect 910 570 1050 580
rect 1310 570 1320 580
rect 1330 570 1340 580
rect 1380 570 1430 580
rect 2170 570 2190 580
rect 3110 570 3120 580
rect 4070 570 4080 580
rect 4370 570 4390 580
rect 4460 570 4530 580
rect 4560 570 4570 580
rect 4650 570 4690 580
rect 4760 570 4800 580
rect 4870 570 4890 580
rect 6640 570 6710 580
rect 6870 570 6880 580
rect 6910 570 7020 580
rect 7160 570 7190 580
rect 7200 570 7310 580
rect 9090 570 9100 580
rect 9630 570 9660 580
rect 9960 570 9970 580
rect 340 560 370 570
rect 600 560 650 570
rect 920 560 1050 570
rect 1280 560 1440 570
rect 3040 560 3110 570
rect 4350 560 4460 570
rect 4470 560 4510 570
rect 4640 560 4670 570
rect 4770 560 4800 570
rect 4860 560 4900 570
rect 4940 560 4950 570
rect 6650 560 6720 570
rect 6870 560 6880 570
rect 6910 560 7030 570
rect 7160 560 7300 570
rect 9180 560 9190 570
rect 9230 560 9240 570
rect 9290 560 9300 570
rect 9650 560 9660 570
rect 9780 560 9790 570
rect 9930 560 9940 570
rect 9950 560 9960 570
rect 330 550 360 560
rect 550 550 560 560
rect 580 550 650 560
rect 930 550 1050 560
rect 1260 550 1400 560
rect 1440 550 1450 560
rect 3010 550 3030 560
rect 3080 550 3100 560
rect 4330 550 4430 560
rect 4460 550 4480 560
rect 4550 550 4570 560
rect 4630 550 4670 560
rect 4770 550 4810 560
rect 4840 550 4900 560
rect 6660 550 6730 560
rect 6880 550 6890 560
rect 6910 550 7030 560
rect 7140 550 7310 560
rect 9190 550 9230 560
rect 330 540 360 550
rect 540 540 650 550
rect 930 540 1050 550
rect 1250 540 1390 550
rect 1440 540 1470 550
rect 3000 540 3010 550
rect 4250 540 4470 550
rect 4550 540 4580 550
rect 4600 540 4660 550
rect 4770 540 4800 550
rect 4840 540 4900 550
rect 6660 540 6740 550
rect 6880 540 6890 550
rect 6930 540 7030 550
rect 7130 540 7300 550
rect 9190 540 9220 550
rect 9280 540 9290 550
rect 9980 540 9990 550
rect 340 530 350 540
rect 530 530 640 540
rect 940 530 1050 540
rect 1240 530 1310 540
rect 1330 530 1370 540
rect 1440 530 1480 540
rect 2980 530 2990 540
rect 4240 530 4450 540
rect 4550 530 4650 540
rect 4770 530 4790 540
rect 4850 530 4900 540
rect 6660 530 6750 540
rect 6880 530 6890 540
rect 6920 530 7030 540
rect 7120 530 7300 540
rect 9210 530 9220 540
rect 9230 530 9240 540
rect 340 520 370 530
rect 510 520 630 530
rect 950 520 1040 530
rect 1230 520 1260 530
rect 1460 520 1490 530
rect 2970 520 2980 530
rect 4220 520 4360 530
rect 4560 520 4640 530
rect 4770 520 4790 530
rect 4860 520 4900 530
rect 6660 520 6750 530
rect 6880 520 6890 530
rect 6940 520 7080 530
rect 7130 520 7300 530
rect 9210 520 9230 530
rect 9990 520 9990 530
rect 350 510 370 520
rect 490 510 580 520
rect 990 510 1030 520
rect 1220 510 1260 520
rect 1490 510 1500 520
rect 2950 510 2970 520
rect 4220 510 4280 520
rect 4610 510 4630 520
rect 4760 510 4790 520
rect 4870 510 4900 520
rect 4950 510 4960 520
rect 6660 510 6750 520
rect 6890 510 6900 520
rect 6940 510 7110 520
rect 7120 510 7290 520
rect 9190 510 9220 520
rect 9920 510 9930 520
rect 9990 510 9990 520
rect 200 500 250 510
rect 360 500 380 510
rect 470 500 530 510
rect 1200 500 1250 510
rect 1490 500 1500 510
rect 2910 500 2940 510
rect 4210 500 4260 510
rect 4770 500 4790 510
rect 4870 500 4900 510
rect 6660 500 6770 510
rect 6880 500 6900 510
rect 6940 500 7280 510
rect 9190 500 9220 510
rect 180 490 290 500
rect 370 490 390 500
rect 460 490 520 500
rect 1190 490 1200 500
rect 1480 490 1490 500
rect 2870 490 2900 500
rect 4200 490 4260 500
rect 4770 490 4790 500
rect 4860 490 4900 500
rect 6670 490 6760 500
rect 6890 490 6900 500
rect 6940 490 7280 500
rect 9140 490 9210 500
rect 9250 490 9260 500
rect 9860 490 9890 500
rect 9900 490 9910 500
rect 160 480 310 490
rect 380 480 400 490
rect 440 480 500 490
rect 1170 480 1180 490
rect 1480 480 1490 490
rect 1510 480 1530 490
rect 2850 480 2870 490
rect 4190 480 4250 490
rect 4760 480 4800 490
rect 4860 480 4900 490
rect 6690 480 6770 490
rect 6900 480 6910 490
rect 6950 480 7280 490
rect 9130 480 9210 490
rect 9880 480 9900 490
rect 150 470 320 480
rect 390 470 490 480
rect 1160 470 1170 480
rect 1480 470 1520 480
rect 1530 470 1540 480
rect 2810 470 2840 480
rect 4180 470 4240 480
rect 4760 470 4790 480
rect 4860 470 4910 480
rect 6700 470 6790 480
rect 6810 470 6830 480
rect 6890 470 6910 480
rect 6940 470 7280 480
rect 9130 470 9190 480
rect 9880 470 9900 480
rect 9930 470 9940 480
rect 140 460 330 470
rect 390 460 470 470
rect 1150 460 1160 470
rect 1480 460 1510 470
rect 2140 460 2150 470
rect 2780 460 2800 470
rect 4180 460 4230 470
rect 4760 460 4790 470
rect 4870 460 4910 470
rect 6690 460 6800 470
rect 6810 460 6840 470
rect 6900 460 6940 470
rect 6950 460 7280 470
rect 9130 460 9180 470
rect 9190 460 9200 470
rect 9240 460 9250 470
rect 9300 460 9320 470
rect 9910 460 9930 470
rect 130 450 160 460
rect 240 450 340 460
rect 400 450 470 460
rect 1140 450 1150 460
rect 1470 450 1510 460
rect 2730 450 2740 460
rect 4170 450 4220 460
rect 4760 450 4780 460
rect 4880 450 4920 460
rect 6700 450 6870 460
rect 6900 450 7270 460
rect 9070 450 9100 460
rect 9110 450 9170 460
rect 9230 450 9240 460
rect 9290 450 9320 460
rect 9370 450 9410 460
rect 120 440 140 450
rect 270 440 350 450
rect 420 440 460 450
rect 1470 440 1510 450
rect 1540 440 1550 450
rect 2020 440 2030 450
rect 4170 440 4210 450
rect 4750 440 4780 450
rect 4880 440 4920 450
rect 4960 440 4970 450
rect 6700 440 6870 450
rect 6890 440 7260 450
rect 9060 440 9090 450
rect 9120 440 9130 450
rect 9160 440 9170 450
rect 9180 440 9190 450
rect 9220 440 9230 450
rect 9320 440 9340 450
rect 9860 440 9880 450
rect 110 430 120 440
rect 280 430 350 440
rect 420 430 460 440
rect 1470 430 1510 440
rect 1860 430 1870 440
rect 4160 430 4210 440
rect 4740 430 4770 440
rect 4890 430 4910 440
rect 6720 430 6860 440
rect 6880 430 7250 440
rect 9010 430 9020 440
rect 9060 430 9080 440
rect 9150 430 9160 440
rect 9280 430 9290 440
rect 9330 430 9350 440
rect 100 420 110 430
rect 280 420 370 430
rect 430 420 460 430
rect 1120 420 1130 430
rect 1470 420 1500 430
rect 1690 420 1710 430
rect 1830 420 1860 430
rect 2580 420 2600 430
rect 4160 420 4200 430
rect 4740 420 4770 430
rect 4900 420 4910 430
rect 6720 420 7240 430
rect 9020 420 9030 430
rect 9060 420 9080 430
rect 9140 420 9160 430
rect 9210 420 9220 430
rect 9300 420 9380 430
rect 90 410 100 420
rect 290 410 370 420
rect 430 410 470 420
rect 1110 410 1120 420
rect 1470 410 1500 420
rect 2340 410 2350 420
rect 4150 410 4190 420
rect 4740 410 4760 420
rect 6730 410 7240 420
rect 9030 410 9040 420
rect 9140 410 9160 420
rect 9290 410 9300 420
rect 9320 410 9340 420
rect 9390 410 9400 420
rect 90 400 100 410
rect 300 400 380 410
rect 440 400 480 410
rect 1470 400 1500 410
rect 2420 400 2460 410
rect 4150 400 4190 410
rect 4730 400 4760 410
rect 6730 400 7240 410
rect 9270 400 9290 410
rect 9310 400 9330 410
rect 9390 400 9400 410
rect 9980 400 9990 410
rect 80 390 90 400
rect 300 390 390 400
rect 450 390 470 400
rect 1100 390 1110 400
rect 1470 390 1500 400
rect 4140 390 4190 400
rect 4730 390 4760 400
rect 6740 390 7230 400
rect 9130 390 9140 400
rect 9150 390 9160 400
rect 9260 390 9320 400
rect 9380 390 9410 400
rect 9990 390 9990 400
rect 70 380 80 390
rect 300 380 390 390
rect 450 380 470 390
rect 1090 380 1100 390
rect 1230 380 1250 390
rect 1470 380 1490 390
rect 4140 380 4190 390
rect 4730 380 4750 390
rect 6760 380 7220 390
rect 9120 380 9130 390
rect 9190 380 9200 390
rect 9250 380 9260 390
rect 9280 380 9320 390
rect 9410 380 9420 390
rect 300 370 390 380
rect 450 370 480 380
rect 1230 370 1240 380
rect 1250 370 1260 380
rect 1470 370 1490 380
rect 4140 370 4190 380
rect 4730 370 4760 380
rect 4920 370 4930 380
rect 6770 370 7220 380
rect 9110 370 9120 380
rect 9140 370 9150 380
rect 9700 370 9710 380
rect 60 360 70 370
rect 290 360 380 370
rect 450 360 470 370
rect 1220 360 1230 370
rect 1470 360 1480 370
rect 4140 360 4190 370
rect 4300 360 4320 370
rect 4340 360 4350 370
rect 4740 360 4760 370
rect 4910 360 4940 370
rect 6780 360 7220 370
rect 9110 360 9120 370
rect 9240 360 9250 370
rect 9310 360 9320 370
rect 290 350 380 360
rect 450 350 460 360
rect 1070 350 1080 360
rect 4130 350 4190 360
rect 4280 350 4350 360
rect 4740 350 4760 360
rect 4900 350 4960 360
rect 6780 350 7210 360
rect 9130 350 9140 360
rect 9170 350 9180 360
rect 9230 350 9240 360
rect 9430 350 9440 360
rect 50 340 60 350
rect 280 340 380 350
rect 1060 340 1070 350
rect 4120 340 4180 350
rect 4280 340 4360 350
rect 4740 340 4770 350
rect 4900 340 4980 350
rect 6790 340 7200 350
rect 9100 340 9110 350
rect 9220 340 9230 350
rect 9940 340 9970 350
rect 9990 340 9990 350
rect 40 330 50 340
rect 100 330 110 340
rect 270 330 390 340
rect 530 330 690 340
rect 4110 330 4170 340
rect 4220 330 4230 340
rect 4260 330 4360 340
rect 4750 330 4770 340
rect 4820 330 4830 340
rect 4850 330 4860 340
rect 4880 330 4960 340
rect 4970 330 4980 340
rect 6800 330 7210 340
rect 9120 330 9130 340
rect 9500 330 9510 340
rect 9980 330 9990 340
rect 40 320 50 330
rect 100 320 120 330
rect 260 320 390 330
rect 500 320 700 330
rect 4090 320 4220 330
rect 4250 320 4370 330
rect 4750 320 4800 330
rect 4810 320 4960 330
rect 4970 320 4980 330
rect 6820 320 7170 330
rect 9150 320 9160 330
rect 9210 320 9220 330
rect 9410 320 9420 330
rect 9490 320 9530 330
rect 30 310 40 320
rect 70 310 130 320
rect 240 310 400 320
rect 480 310 720 320
rect 1040 310 1050 320
rect 4080 310 4220 320
rect 4240 310 4390 320
rect 4410 310 4420 320
rect 4430 310 4460 320
rect 4500 310 4530 320
rect 4750 310 4950 320
rect 4970 310 4980 320
rect 6840 310 7120 320
rect 9080 310 9090 320
rect 9150 310 9160 320
rect 9410 310 9420 320
rect 30 300 40 310
rect 70 300 140 310
rect 230 300 400 310
rect 470 300 790 310
rect 4070 300 4140 310
rect 4150 300 4180 310
rect 4240 300 4460 310
rect 4490 300 4530 310
rect 4740 300 4960 310
rect 4970 300 4980 310
rect 6860 300 7110 310
rect 9140 300 9150 310
rect 9420 300 9430 310
rect 9720 300 9740 310
rect 9750 300 9760 310
rect 70 290 150 300
rect 210 290 400 300
rect 460 290 510 300
rect 550 290 820 300
rect 4070 290 4120 300
rect 4230 290 4470 300
rect 4490 290 4530 300
rect 4710 290 4950 300
rect 4960 290 4970 300
rect 6890 290 7050 300
rect 7080 290 7090 300
rect 7100 290 7110 300
rect 9430 290 9440 300
rect 9500 290 9520 300
rect 9560 290 9580 300
rect 9690 290 9700 300
rect 9720 290 9750 300
rect 9810 290 9820 300
rect 60 280 400 290
rect 450 280 520 290
rect 560 280 650 290
rect 680 280 850 290
rect 4070 280 4120 290
rect 4220 280 4470 290
rect 4480 280 4530 290
rect 4680 280 4950 290
rect 6900 280 6920 290
rect 6930 280 6970 290
rect 7000 280 7030 290
rect 7050 280 7060 290
rect 9060 280 9070 290
rect 9200 280 9210 290
rect 9440 280 9450 290
rect 9500 280 9520 290
rect 9550 280 9580 290
rect 9620 280 9640 290
rect 9810 280 9820 290
rect 20 270 30 280
rect 50 270 400 280
rect 450 270 520 280
rect 560 270 640 280
rect 680 270 860 280
rect 1030 270 1040 280
rect 4070 270 4110 280
rect 4210 270 4220 280
rect 4230 270 4530 280
rect 4670 270 4950 280
rect 6990 270 7010 280
rect 7050 270 7070 280
rect 9190 270 9200 280
rect 9310 270 9320 280
rect 9450 270 9470 280
rect 9500 270 9530 280
rect 9560 270 9570 280
rect 9580 270 9590 280
rect 9810 270 9820 280
rect 9990 270 9990 280
rect 20 260 400 270
rect 440 260 520 270
rect 550 260 640 270
rect 680 260 870 270
rect 1230 260 1240 270
rect 4080 260 4110 270
rect 4200 260 4540 270
rect 4660 260 4940 270
rect 6990 260 7010 270
rect 7050 260 7060 270
rect 9050 260 9060 270
rect 9190 260 9200 270
rect 9300 260 9310 270
rect 9440 260 9480 270
rect 9520 260 9540 270
rect 9550 260 9580 270
rect 9790 260 9800 270
rect 9820 260 9840 270
rect 9980 260 9990 270
rect 20 250 130 260
rect 190 250 390 260
rect 440 250 520 260
rect 550 250 630 260
rect 680 250 870 260
rect 4090 250 4110 260
rect 4190 250 4540 260
rect 4550 250 4570 260
rect 4600 250 4610 260
rect 4660 250 4940 260
rect 8900 250 8930 260
rect 9040 250 9050 260
rect 9190 250 9200 260
rect 9280 250 9300 260
rect 9460 250 9480 260
rect 9530 250 9550 260
rect 9590 250 9600 260
rect 9820 250 9850 260
rect 9990 250 9990 260
rect 20 240 120 250
rect 200 240 380 250
rect 440 240 520 250
rect 550 240 630 250
rect 680 240 870 250
rect 1020 240 1030 250
rect 1220 240 1230 250
rect 4090 240 4110 250
rect 4180 240 4540 250
rect 4550 240 4560 250
rect 4600 240 4620 250
rect 4660 240 4840 250
rect 4850 240 4950 250
rect 8890 240 8950 250
rect 9180 240 9190 250
rect 9290 240 9300 250
rect 9330 240 9340 250
rect 9380 240 9390 250
rect 9400 240 9410 250
rect 9440 240 9450 250
rect 9490 240 9500 250
rect 9590 240 9610 250
rect 9810 240 9820 250
rect 20 230 120 240
rect 210 230 380 240
rect 430 230 530 240
rect 540 230 630 240
rect 680 230 870 240
rect 1020 230 1030 240
rect 1220 230 1230 240
rect 4100 230 4110 240
rect 4170 230 4210 240
rect 4220 230 4530 240
rect 4550 230 4570 240
rect 4590 230 4620 240
rect 4660 230 4840 240
rect 4870 230 4880 240
rect 4890 230 4950 240
rect 8880 230 8970 240
rect 9030 230 9040 240
rect 9160 230 9170 240
rect 9300 230 9330 240
rect 9420 230 9430 240
rect 9450 230 9460 240
rect 9470 230 9510 240
rect 9780 230 9790 240
rect 10 220 90 230
rect 210 220 370 230
rect 430 220 530 230
rect 540 220 620 230
rect 680 220 870 230
rect 1020 220 1030 230
rect 4100 220 4130 230
rect 4160 220 4200 230
rect 4220 220 4230 230
rect 4240 220 4540 230
rect 4550 220 4560 230
rect 4590 220 4630 230
rect 4650 220 4850 230
rect 4890 220 4940 230
rect 4990 220 5000 230
rect 8890 220 8960 230
rect 9300 220 9330 230
rect 9400 220 9410 230
rect 9430 220 9500 230
rect 9510 220 9520 230
rect 9780 220 9790 230
rect 9850 220 9860 230
rect 10 210 60 220
rect 210 210 360 220
rect 430 210 520 220
rect 540 210 620 220
rect 680 210 880 220
rect 1020 210 1030 220
rect 4110 210 4130 220
rect 4160 210 4180 220
rect 4250 210 4330 220
rect 4350 210 4560 220
rect 4590 210 4630 220
rect 4650 210 4850 220
rect 4880 210 4940 220
rect 8890 210 8970 220
rect 9020 210 9030 220
rect 9090 210 9100 220
rect 9310 210 9320 220
rect 9350 210 9360 220
rect 9400 210 9410 220
rect 9930 210 9940 220
rect 9950 210 9960 220
rect 10 200 60 210
rect 220 200 340 210
rect 430 200 610 210
rect 680 200 860 210
rect 4120 200 4150 210
rect 4250 200 4320 210
rect 4380 200 4520 210
rect 4540 200 4560 210
rect 4590 200 4630 210
rect 4640 200 4920 210
rect 4930 200 4950 210
rect 8870 200 8880 210
rect 8910 200 8930 210
rect 8940 200 8960 210
rect 9150 200 9160 210
rect 9300 200 9310 210
rect 9680 200 9690 210
rect 9780 200 9800 210
rect 9940 200 9960 210
rect 10 190 70 200
rect 220 190 330 200
rect 450 190 610 200
rect 690 190 860 200
rect 4130 190 4150 200
rect 4250 190 4290 200
rect 4400 190 4420 200
rect 4440 190 4490 200
rect 4540 190 4560 200
rect 4580 190 4930 200
rect 8860 190 8870 200
rect 8910 190 8920 200
rect 9040 190 9050 200
rect 9180 190 9190 200
rect 9680 190 9700 200
rect 9740 190 9760 200
rect 9790 190 9800 200
rect 9930 190 9950 200
rect 10 180 80 190
rect 220 180 320 190
rect 470 180 600 190
rect 690 180 840 190
rect 4140 180 4160 190
rect 4540 180 4560 190
rect 4580 180 4930 190
rect 8880 180 8890 190
rect 8900 180 8910 190
rect 9130 180 9140 190
rect 9300 180 9310 190
rect 9690 180 9700 190
rect 9730 180 9740 190
rect 9840 180 9850 190
rect 9860 180 9870 190
rect 9890 180 9910 190
rect 9960 180 9970 190
rect 10 170 100 180
rect 230 170 250 180
rect 260 170 310 180
rect 490 170 580 180
rect 700 170 830 180
rect 4150 170 4160 180
rect 4540 170 4550 180
rect 4580 170 4940 180
rect 8860 170 8890 180
rect 9070 170 9080 180
rect 9160 170 9190 180
rect 9710 170 9720 180
rect 9840 170 9850 180
rect 9950 170 9960 180
rect 10 160 110 170
rect 250 160 280 170
rect 510 160 550 170
rect 710 160 810 170
rect 1010 160 1020 170
rect 4160 160 4170 170
rect 4540 160 4550 170
rect 4580 160 4820 170
rect 4900 160 4940 170
rect 5000 160 5010 170
rect 8850 160 8860 170
rect 9000 160 9010 170
rect 9180 160 9190 170
rect 9330 160 9340 170
rect 9550 160 9560 170
rect 9690 160 9710 170
rect 0 150 110 160
rect 250 150 260 160
rect 720 150 780 160
rect 4170 150 4180 160
rect 4580 150 4820 160
rect 4920 150 4980 160
rect 8870 150 8880 160
rect 9010 150 9020 160
rect 9160 150 9170 160
rect 9550 150 9570 160
rect 9600 150 9610 160
rect 9700 150 9710 160
rect 9950 150 9970 160
rect 0 140 110 150
rect 4180 140 4190 150
rect 4570 140 4810 150
rect 4940 140 4980 150
rect 9130 140 9140 150
rect 9340 140 9350 150
rect 9560 140 9570 150
rect 9580 140 9610 150
rect 9620 140 9630 150
rect 9650 140 9660 150
rect 9950 140 9990 150
rect 0 130 110 140
rect 4570 130 4610 140
rect 4630 130 4700 140
rect 4730 130 4800 140
rect 4960 130 4980 140
rect 5010 130 5020 140
rect 8830 130 8840 140
rect 9100 130 9110 140
rect 9600 130 9610 140
rect 9970 130 9980 140
rect 0 120 100 130
rect 1010 120 1020 130
rect 4570 120 4600 130
rect 4630 120 4690 130
rect 4740 120 4800 130
rect 4970 120 4980 130
rect 9100 120 9110 130
rect 9710 120 9720 130
rect 9980 120 9990 130
rect 0 110 100 120
rect 1010 110 1020 120
rect 4570 110 4590 120
rect 4630 110 4680 120
rect 4740 110 4780 120
rect 4960 110 4970 120
rect 8930 110 8940 120
rect 9140 110 9150 120
rect 9380 110 9400 120
rect 9410 110 9420 120
rect 9860 110 9880 120
rect 9920 110 9940 120
rect 0 100 100 110
rect 4230 100 4240 110
rect 4560 100 4580 110
rect 4640 100 4660 110
rect 4750 100 4770 110
rect 4950 100 4970 110
rect 8830 100 8840 110
rect 8930 100 8940 110
rect 9090 100 9100 110
rect 9140 100 9150 110
rect 9410 100 9430 110
rect 9490 100 9500 110
rect 9570 100 9580 110
rect 9640 100 9650 110
rect 9860 100 9870 110
rect 9880 100 9890 110
rect 9950 100 9960 110
rect 0 90 90 100
rect 4240 90 4250 100
rect 4950 90 4970 100
rect 8800 90 8810 100
rect 9180 90 9190 100
rect 9430 90 9440 100
rect 9870 90 9890 100
rect 9900 90 9920 100
rect 9950 90 9970 100
rect 0 80 100 90
rect 1020 80 1030 90
rect 4250 80 4260 90
rect 4940 80 4970 90
rect 8930 80 8940 90
rect 9590 80 9600 90
rect 9900 80 9910 90
rect 9950 80 9970 90
rect 20 70 100 80
rect 1020 70 1030 80
rect 4940 70 4980 80
rect 8900 70 8930 80
rect 9010 70 9020 80
rect 9060 70 9070 80
rect 9080 70 9090 80
rect 9140 70 9150 80
rect 9550 70 9560 80
rect 9660 70 9680 80
rect 9920 70 9930 80
rect 9940 70 9960 80
rect 20 60 100 70
rect 1020 60 1030 70
rect 4280 60 4290 70
rect 4940 60 4980 70
rect 8770 60 8780 70
rect 8930 60 8940 70
rect 9030 60 9060 70
rect 9070 60 9090 70
rect 9150 60 9160 70
rect 9470 60 9480 70
rect 9540 60 9560 70
rect 9580 60 9590 70
rect 9710 60 9720 70
rect 9740 60 9750 70
rect 9950 60 9960 70
rect 20 50 100 60
rect 1020 50 1030 60
rect 4300 50 4310 60
rect 4940 50 4980 60
rect 5040 50 5050 60
rect 8900 50 8940 60
rect 9070 50 9080 60
rect 9090 50 9100 60
rect 9290 50 9300 60
rect 9560 50 9570 60
rect 9580 50 9590 60
rect 9610 50 9640 60
rect 9660 50 9670 60
rect 9740 50 9750 60
rect 9930 50 9940 60
rect 9950 50 9960 60
rect 20 40 100 50
rect 1020 40 1030 50
rect 4310 40 4330 50
rect 4940 40 4980 50
rect 8920 40 8930 50
rect 9010 40 9020 50
rect 9590 40 9630 50
rect 9670 40 9680 50
rect 9740 40 9750 50
rect 9930 40 9940 50
rect 9970 40 9990 50
rect 20 30 100 40
rect 4330 30 4340 40
rect 4950 30 4980 40
rect 9020 30 9030 40
rect 9080 30 9090 40
rect 9600 30 9610 40
rect 9620 30 9630 40
rect 9670 30 9690 40
rect 9930 30 9940 40
rect 9980 30 9990 40
rect 20 20 100 30
rect 1290 20 1310 30
rect 4340 20 4350 30
rect 4940 20 4980 30
rect 8920 20 8930 30
rect 9030 20 9040 30
rect 9100 20 9110 30
rect 9160 20 9170 30
rect 9500 20 9520 30
rect 9580 20 9590 30
rect 9610 20 9630 30
rect 9660 20 9670 30
rect 9710 20 9720 30
rect 9770 20 9780 30
rect 9930 20 9940 30
rect 10 10 90 20
rect 1280 10 1290 20
rect 1310 10 1320 20
rect 4350 10 4360 20
rect 4930 10 4980 20
rect 5050 10 5060 20
rect 8610 10 8630 20
rect 8720 10 8730 20
rect 9110 10 9120 20
rect 9590 10 9600 20
rect 9630 10 9640 20
rect 9660 10 9670 20
rect 9710 10 9720 20
rect 9780 10 9790 20
rect 9940 10 9950 20
rect 9960 10 9980 20
rect 0 0 90 10
rect 1010 0 1020 10
rect 1280 0 1290 10
rect 1310 0 1320 10
rect 4660 0 4710 10
rect 4910 0 4980 10
rect 8600 0 8610 10
rect 8670 0 8680 10
rect 8790 0 8800 10
rect 9020 0 9030 10
rect 9110 0 9120 10
rect 9600 0 9610 10
rect 9640 0 9670 10
rect 9720 0 9740 10
rect 9980 0 9990 10
<< metal4 >>
rect 0 7490 2160 7500
rect 3340 7490 3560 7500
rect 3810 7490 5020 7500
rect 5110 7490 9530 7500
rect 0 7480 2150 7490
rect 3340 7480 3560 7490
rect 3820 7480 5030 7490
rect 5120 7480 9540 7490
rect 0 7470 2140 7480
rect 3340 7470 3560 7480
rect 3680 7470 3730 7480
rect 3820 7470 5040 7480
rect 5130 7470 9500 7480
rect 9510 7470 9540 7480
rect 0 7460 2120 7470
rect 3330 7460 3560 7470
rect 3670 7460 3760 7470
rect 3830 7460 5070 7470
rect 5130 7460 9500 7470
rect 9510 7460 9540 7470
rect 0 7450 2120 7460
rect 3330 7450 3560 7460
rect 3670 7450 3780 7460
rect 3830 7450 5060 7460
rect 5140 7450 9500 7460
rect 9510 7450 9540 7460
rect 0 7440 2100 7450
rect 3330 7440 3560 7450
rect 3660 7440 3790 7450
rect 3840 7440 5060 7450
rect 5070 7440 5080 7450
rect 5140 7440 9540 7450
rect 0 7430 2100 7440
rect 3330 7430 3570 7440
rect 3660 7430 3800 7440
rect 3850 7430 5090 7440
rect 5140 7430 9540 7440
rect 0 7420 2090 7430
rect 3330 7420 3570 7430
rect 3660 7420 3810 7430
rect 3850 7420 5080 7430
rect 5090 7420 5100 7430
rect 5150 7420 9540 7430
rect 0 7410 2080 7420
rect 3330 7410 3580 7420
rect 3650 7410 3810 7420
rect 3850 7410 5080 7420
rect 5090 7410 5110 7420
rect 5170 7410 9540 7420
rect 0 7400 2070 7410
rect 3340 7400 3590 7410
rect 3650 7400 3780 7410
rect 3790 7400 3820 7410
rect 3860 7400 5090 7410
rect 5100 7400 5120 7410
rect 5170 7400 9540 7410
rect 0 7390 2070 7400
rect 3340 7390 3600 7400
rect 3640 7390 3830 7400
rect 3860 7390 5120 7400
rect 5180 7390 9540 7400
rect 0 7380 2060 7390
rect 3340 7380 3620 7390
rect 3640 7380 3840 7390
rect 3870 7380 5120 7390
rect 5150 7380 5160 7390
rect 5180 7380 9500 7390
rect 9510 7380 9540 7390
rect 0 7370 2050 7380
rect 3340 7370 3840 7380
rect 3880 7370 5170 7380
rect 5180 7370 9500 7380
rect 9510 7370 9540 7380
rect 0 7360 2040 7370
rect 3350 7360 3850 7370
rect 3880 7360 5160 7370
rect 5180 7360 9540 7370
rect 0 7350 2030 7360
rect 3360 7350 3850 7360
rect 3880 7350 5160 7360
rect 5170 7350 5190 7360
rect 5200 7350 9550 7360
rect 0 7340 2020 7350
rect 3360 7340 3860 7350
rect 3890 7340 5140 7350
rect 5150 7340 9550 7350
rect 0 7330 2010 7340
rect 3370 7330 3860 7340
rect 3890 7330 5190 7340
rect 5210 7330 9510 7340
rect 9520 7330 9550 7340
rect 0 7320 2010 7330
rect 3360 7320 3840 7330
rect 3850 7320 3870 7330
rect 3890 7320 9510 7330
rect 9520 7320 9550 7330
rect 9850 7320 9870 7330
rect 0 7310 2000 7320
rect 3370 7310 3380 7320
rect 3390 7310 3870 7320
rect 3900 7310 5200 7320
rect 5230 7310 9510 7320
rect 9520 7310 9550 7320
rect 9850 7310 9880 7320
rect 0 7300 2000 7310
rect 3370 7300 3380 7310
rect 3390 7300 3400 7310
rect 3410 7300 3820 7310
rect 3830 7300 3870 7310
rect 3900 7300 5210 7310
rect 5230 7300 9550 7310
rect 9860 7300 9880 7310
rect 0 7290 1990 7300
rect 3370 7290 3400 7300
rect 3410 7290 3820 7300
rect 3860 7290 3880 7300
rect 3910 7290 5210 7300
rect 5220 7290 5230 7300
rect 5250 7290 9550 7300
rect 9850 7290 9880 7300
rect 0 7280 1990 7290
rect 3370 7280 3380 7290
rect 3390 7280 3400 7290
rect 3420 7280 3830 7290
rect 3860 7280 3880 7290
rect 3910 7280 5200 7290
rect 5210 7280 5230 7290
rect 5240 7280 9550 7290
rect 9860 7280 9880 7290
rect 0 7270 1980 7280
rect 3370 7270 3380 7280
rect 3390 7270 3400 7280
rect 3430 7270 3830 7280
rect 3870 7270 3880 7280
rect 3920 7270 9300 7280
rect 9330 7270 9550 7280
rect 9860 7270 9880 7280
rect 0 7260 1980 7270
rect 3390 7260 3400 7270
rect 3440 7260 3830 7270
rect 3870 7260 3890 7270
rect 3910 7260 6550 7270
rect 6590 7260 9290 7270
rect 9340 7260 9550 7270
rect 9860 7260 9880 7270
rect 0 7250 1980 7260
rect 3390 7250 3400 7260
rect 3440 7250 3820 7260
rect 3870 7250 3890 7260
rect 3920 7250 6540 7260
rect 6600 7250 9260 7260
rect 9350 7250 9550 7260
rect 9860 7250 9880 7260
rect 0 7240 1970 7250
rect 3380 7240 3390 7250
rect 3440 7240 3830 7250
rect 3870 7240 3880 7250
rect 3920 7240 6540 7250
rect 6600 7240 9260 7250
rect 9370 7240 9550 7250
rect 9860 7240 9880 7250
rect 0 7230 1960 7240
rect 3390 7230 3410 7240
rect 3440 7230 3830 7240
rect 3930 7230 6480 7240
rect 6490 7230 6500 7240
rect 6510 7230 6530 7240
rect 6590 7230 8970 7240
rect 8990 7230 9260 7240
rect 9370 7230 9560 7240
rect 0 7220 1960 7230
rect 3390 7220 3400 7230
rect 3450 7220 3830 7230
rect 3880 7220 3890 7230
rect 3930 7220 6490 7230
rect 6580 7220 8970 7230
rect 9030 7220 9300 7230
rect 9360 7220 9570 7230
rect 0 7210 1950 7220
rect 3410 7210 3420 7220
rect 3450 7210 3830 7220
rect 3930 7210 6490 7220
rect 6560 7210 8970 7220
rect 9010 7210 9020 7220
rect 9030 7210 9310 7220
rect 9360 7210 9570 7220
rect 0 7200 1940 7210
rect 3400 7200 3410 7210
rect 3450 7200 3830 7210
rect 3940 7200 6500 7210
rect 6560 7200 6600 7210
rect 6650 7200 8970 7210
rect 9020 7200 9040 7210
rect 9060 7200 9320 7210
rect 9370 7200 9570 7210
rect 0 7190 1930 7200
rect 3450 7190 3810 7200
rect 3940 7190 6500 7200
rect 6560 7190 6580 7200
rect 6650 7190 8980 7200
rect 9010 7190 9330 7200
rect 9370 7190 9580 7200
rect 0 7180 1930 7190
rect 3410 7180 3420 7190
rect 3450 7180 3740 7190
rect 3750 7180 3810 7190
rect 3940 7180 6510 7190
rect 6560 7180 6580 7190
rect 6660 7180 6690 7190
rect 6710 7180 9330 7190
rect 9380 7180 9580 7190
rect 0 7170 1930 7180
rect 3410 7170 3440 7180
rect 3450 7170 3730 7180
rect 3750 7170 3810 7180
rect 3950 7170 6510 7180
rect 6560 7170 6570 7180
rect 6720 7170 9030 7180
rect 9050 7170 9350 7180
rect 9380 7170 9580 7180
rect 0 7160 1930 7170
rect 3360 7160 3390 7170
rect 3400 7160 3730 7170
rect 3750 7160 3810 7170
rect 3950 7160 5280 7170
rect 5300 7160 6520 7170
rect 6720 7160 9580 7170
rect 0 7150 1920 7160
rect 3350 7150 3500 7160
rect 3530 7150 3690 7160
rect 3700 7150 3730 7160
rect 3750 7150 3800 7160
rect 3810 7150 3820 7160
rect 3950 7150 5290 7160
rect 5300 7150 6530 7160
rect 6720 7150 8940 7160
rect 8950 7150 9570 7160
rect 0 7140 1910 7150
rect 3370 7140 3490 7150
rect 3540 7140 3680 7150
rect 3700 7140 3730 7150
rect 3750 7140 3790 7150
rect 3810 7140 3820 7150
rect 3950 7140 6460 7150
rect 6470 7140 6530 7150
rect 6720 7140 8860 7150
rect 8880 7140 8930 7150
rect 8940 7140 9570 7150
rect 0 7130 1910 7140
rect 3400 7130 3490 7140
rect 3540 7130 3660 7140
rect 3710 7130 3730 7140
rect 3750 7130 3780 7140
rect 3810 7130 3820 7140
rect 3950 7130 6540 7140
rect 6720 7130 8860 7140
rect 8880 7130 8930 7140
rect 8940 7130 9570 7140
rect 0 7120 1910 7130
rect 3460 7120 3510 7130
rect 3550 7120 3650 7130
rect 3710 7120 3730 7130
rect 3750 7120 3770 7130
rect 3950 7120 6540 7130
rect 6710 7120 9560 7130
rect 0 7110 1910 7120
rect 3470 7110 3520 7120
rect 3550 7110 3630 7120
rect 3720 7110 3730 7120
rect 3750 7110 3760 7120
rect 3950 7110 6540 7120
rect 6700 7110 8960 7120
rect 8990 7110 9380 7120
rect 9390 7110 9570 7120
rect 0 7100 1900 7110
rect 3480 7100 3490 7110
rect 3500 7100 3520 7110
rect 3560 7100 3630 7110
rect 3960 7100 6550 7110
rect 6700 7100 9380 7110
rect 9400 7100 9500 7110
rect 9530 7100 9570 7110
rect 0 7090 1900 7100
rect 3490 7090 3500 7100
rect 3510 7090 3520 7100
rect 3570 7090 3630 7100
rect 3970 7090 6560 7100
rect 6690 7090 9390 7100
rect 9410 7090 9490 7100
rect 9530 7090 9570 7100
rect 0 7080 1900 7090
rect 3500 7080 3530 7090
rect 3580 7080 3630 7090
rect 3970 7080 6550 7090
rect 6680 7080 8950 7090
rect 8970 7080 9400 7090
rect 9420 7080 9510 7090
rect 9520 7080 9570 7090
rect 0 7070 1900 7080
rect 3510 7070 3540 7080
rect 3580 7070 3620 7080
rect 3970 7070 6550 7080
rect 6680 7070 8960 7080
rect 8970 7070 9570 7080
rect 0 7060 1900 7070
rect 3520 7060 3550 7070
rect 3590 7060 3620 7070
rect 3970 7060 6540 7070
rect 6670 7060 8870 7070
rect 8890 7060 9490 7070
rect 9500 7060 9570 7070
rect 0 7050 1890 7060
rect 3520 7050 3580 7060
rect 3590 7050 3630 7060
rect 3730 7050 3740 7060
rect 3800 7050 3810 7060
rect 3980 7050 6550 7060
rect 6670 7050 8860 7060
rect 8890 7050 9530 7060
rect 9540 7050 9570 7060
rect 0 7040 1890 7050
rect 3540 7040 3630 7050
rect 3790 7040 3810 7050
rect 3970 7040 6530 7050
rect 6560 7040 6570 7050
rect 6680 7040 6710 7050
rect 6720 7040 9570 7050
rect 0 7030 1890 7040
rect 3560 7030 3630 7040
rect 3750 7030 3760 7040
rect 3780 7030 3810 7040
rect 3980 7030 6520 7040
rect 6550 7030 6570 7040
rect 6690 7030 6700 7040
rect 6720 7030 9570 7040
rect 0 7020 1880 7030
rect 1940 7020 1950 7030
rect 3570 7020 3630 7030
rect 3780 7020 3790 7030
rect 3800 7020 3810 7030
rect 3990 7020 6510 7030
rect 6550 7020 6580 7030
rect 6620 7020 6660 7030
rect 6720 7020 9580 7030
rect 0 7010 1880 7020
rect 1930 7010 1940 7020
rect 3590 7010 3600 7020
rect 3620 7010 3640 7020
rect 3760 7010 3800 7020
rect 3990 7010 6500 7020
rect 6540 7010 6570 7020
rect 6620 7010 6700 7020
rect 6720 7010 8940 7020
rect 8960 7010 9580 7020
rect 0 7000 1880 7010
rect 1920 7000 1940 7010
rect 3610 7000 3650 7010
rect 3740 7000 3750 7010
rect 3770 7000 3800 7010
rect 3990 7000 6320 7010
rect 6330 7000 6500 7010
rect 6530 7000 6570 7010
rect 6600 7000 8950 7010
rect 8960 7000 9580 7010
rect 0 6990 1880 7000
rect 1920 6990 1930 7000
rect 3620 6990 3670 7000
rect 3750 6990 3810 7000
rect 3990 6990 6500 7000
rect 6520 6990 6580 7000
rect 6600 6990 9580 7000
rect 0 6980 1940 6990
rect 3640 6980 3690 6990
rect 3740 6980 3810 6990
rect 4000 6980 6500 6990
rect 6510 6980 6580 6990
rect 6590 6980 9580 6990
rect 0 6970 1960 6980
rect 3650 6970 3680 6980
rect 3700 6970 3800 6980
rect 3820 6970 3830 6980
rect 4000 6970 9580 6980
rect 0 6960 1940 6970
rect 1960 6960 1970 6970
rect 3670 6960 3710 6970
rect 3720 6960 3730 6970
rect 3750 6960 3800 6970
rect 3990 6960 8880 6970
rect 8890 6960 9580 6970
rect 0 6950 1930 6960
rect 3290 6950 3300 6960
rect 3710 6950 3810 6960
rect 3990 6950 8610 6960
rect 8630 6950 8910 6960
rect 8920 6950 9580 6960
rect 0 6940 1910 6950
rect 1920 6940 1930 6950
rect 3800 6940 3810 6950
rect 3990 6940 5470 6950
rect 5480 6940 8600 6950
rect 8630 6940 8850 6950
rect 8880 6940 8920 6950
rect 8930 6940 9590 6950
rect 0 6930 1900 6940
rect 3350 6930 3360 6940
rect 3980 6930 8560 6940
rect 8570 6930 8580 6940
rect 8610 6930 8620 6940
rect 8650 6930 8850 6940
rect 8860 6930 8910 6940
rect 8920 6930 9590 6940
rect 0 6920 1890 6930
rect 3350 6920 3390 6930
rect 3980 6920 5480 6930
rect 5500 6920 8440 6930
rect 8450 6920 8550 6930
rect 8560 6920 8570 6930
rect 8590 6920 8620 6930
rect 8640 6920 9590 6930
rect 0 6910 1880 6920
rect 3360 6910 3410 6920
rect 3850 6910 3860 6920
rect 3990 6910 5490 6920
rect 5510 6910 9590 6920
rect 0 6900 1870 6910
rect 3380 6900 3440 6910
rect 3990 6900 5490 6910
rect 5520 6900 8550 6910
rect 8560 6900 9590 6910
rect 0 6890 1870 6900
rect 3380 6890 3460 6900
rect 4000 6890 5500 6900
rect 5520 6890 8550 6900
rect 8560 6890 9070 6900
rect 9080 6890 9590 6900
rect 0 6880 1870 6890
rect 3380 6880 3480 6890
rect 4000 6880 5500 6890
rect 5510 6880 8480 6890
rect 8490 6880 9060 6890
rect 9100 6880 9580 6890
rect 0 6870 1870 6880
rect 3400 6870 3510 6880
rect 4000 6870 5510 6880
rect 5520 6870 5530 6880
rect 5540 6870 8480 6880
rect 8490 6870 8690 6880
rect 8710 6870 9060 6880
rect 9080 6870 9580 6880
rect 0 6860 1910 6870
rect 3400 6860 3520 6870
rect 3990 6860 5520 6870
rect 5530 6860 8470 6870
rect 8500 6860 8600 6870
rect 8610 6860 8700 6870
rect 8710 6860 8760 6870
rect 8770 6860 8790 6870
rect 8810 6860 9040 6870
rect 9050 6860 9580 6870
rect 0 6850 1870 6860
rect 2670 6850 2680 6860
rect 3420 6850 3540 6860
rect 3990 6850 5530 6860
rect 5560 6850 6770 6860
rect 6790 6850 8590 6860
rect 8620 6850 9040 6860
rect 9050 6850 9520 6860
rect 9540 6850 9590 6860
rect 0 6840 1880 6850
rect 2690 6840 2700 6850
rect 3430 6840 3560 6850
rect 3990 6840 5530 6850
rect 5570 6840 8710 6850
rect 8720 6840 9010 6850
rect 9050 6840 9590 6850
rect 0 6830 1880 6840
rect 2730 6830 2760 6840
rect 3300 6830 3330 6840
rect 3430 6830 3580 6840
rect 3970 6830 5540 6840
rect 5590 6830 8720 6840
rect 8730 6830 9030 6840
rect 9050 6830 9590 6840
rect 0 6820 1880 6830
rect 2780 6820 2790 6830
rect 3290 6820 3360 6830
rect 3370 6820 3380 6830
rect 3430 6820 3600 6830
rect 3970 6820 5550 6830
rect 5560 6820 5570 6830
rect 5600 6820 9030 6830
rect 9040 6820 9590 6830
rect 0 6810 1840 6820
rect 1850 6810 1870 6820
rect 2800 6810 2840 6820
rect 3290 6810 3410 6820
rect 3460 6810 3480 6820
rect 3490 6810 3620 6820
rect 3960 6810 5560 6820
rect 5620 6810 9590 6820
rect 0 6800 1850 6810
rect 2880 6800 2890 6810
rect 3290 6800 3430 6810
rect 3480 6800 3630 6810
rect 3960 6800 5570 6810
rect 5610 6800 9590 6810
rect 0 6790 1870 6800
rect 2940 6790 2980 6800
rect 3300 6790 3460 6800
rect 3480 6790 3490 6800
rect 3500 6790 3650 6800
rect 3960 6790 5570 6800
rect 5600 6790 9590 6800
rect 0 6780 1860 6790
rect 1870 6780 1880 6790
rect 3000 6780 3040 6790
rect 3350 6780 3660 6790
rect 3960 6780 5580 6790
rect 5590 6780 9590 6790
rect 0 6770 1860 6780
rect 1970 6770 1990 6780
rect 3070 6770 3080 6780
rect 3090 6770 3150 6780
rect 3380 6770 3680 6780
rect 3960 6770 9590 6780
rect 0 6760 1870 6770
rect 1970 6760 1980 6770
rect 3130 6760 3210 6770
rect 3400 6760 3690 6770
rect 3960 6760 5630 6770
rect 5650 6760 9570 6770
rect 9580 6760 9600 6770
rect 0 6750 1870 6760
rect 1970 6750 1980 6760
rect 3190 6750 3300 6760
rect 3370 6750 3380 6760
rect 3410 6750 3710 6760
rect 3960 6750 5630 6760
rect 5650 6750 9550 6760
rect 9580 6750 9600 6760
rect 0 6740 1860 6750
rect 3250 6740 3350 6750
rect 3360 6740 3380 6750
rect 3400 6740 3410 6750
rect 3420 6740 3720 6750
rect 3960 6740 5620 6750
rect 5640 6740 5650 6750
rect 5660 6740 9550 6750
rect 9580 6740 9590 6750
rect 0 6730 1850 6740
rect 3310 6730 3420 6740
rect 3450 6730 3740 6740
rect 3970 6730 9540 6740
rect 9570 6730 9590 6740
rect 0 6720 1850 6730
rect 3350 6720 3460 6730
rect 3480 6720 3750 6730
rect 3970 6720 8980 6730
rect 8990 6720 9540 6730
rect 9570 6720 9590 6730
rect 0 6710 1830 6720
rect 2390 6710 2430 6720
rect 3390 6710 3480 6720
rect 3510 6710 3760 6720
rect 3970 6710 9530 6720
rect 9570 6710 9590 6720
rect 0 6700 1840 6710
rect 1850 6700 1870 6710
rect 2330 6700 2340 6710
rect 2350 6700 2450 6710
rect 3430 6700 3770 6710
rect 3970 6700 9530 6710
rect 9580 6700 9590 6710
rect 0 6690 1810 6700
rect 1840 6690 1850 6700
rect 2310 6690 2480 6700
rect 3470 6690 3790 6700
rect 3970 6690 9530 6700
rect 9580 6690 9600 6700
rect 0 6680 1790 6690
rect 2280 6680 2480 6690
rect 3490 6680 3800 6690
rect 3970 6680 9520 6690
rect 9580 6680 9600 6690
rect 9980 6680 9990 6690
rect 0 6670 1770 6680
rect 1780 6670 1800 6680
rect 1810 6670 1820 6680
rect 2270 6670 2480 6680
rect 3540 6670 3810 6680
rect 3980 6670 8930 6680
rect 8940 6670 9510 6680
rect 9580 6670 9600 6680
rect 9960 6670 9990 6680
rect 0 6660 1750 6670
rect 1760 6660 1860 6670
rect 2270 6660 2480 6670
rect 3550 6660 3820 6670
rect 3980 6660 8930 6670
rect 8940 6660 9500 6670
rect 9570 6660 9600 6670
rect 9920 6660 9990 6670
rect 0 6650 1850 6660
rect 2270 6650 2490 6660
rect 3570 6650 3840 6660
rect 3980 6650 8570 6660
rect 8580 6650 9500 6660
rect 9570 6650 9600 6660
rect 9890 6650 9990 6660
rect 0 6640 1710 6650
rect 1730 6640 1800 6650
rect 2260 6640 2510 6650
rect 3600 6640 3850 6650
rect 3990 6640 9490 6650
rect 9560 6640 9610 6650
rect 9860 6640 9990 6650
rect 0 6630 1750 6640
rect 2250 6630 2520 6640
rect 3620 6630 3860 6640
rect 3990 6630 9480 6640
rect 9550 6630 9610 6640
rect 9830 6630 9990 6640
rect 0 6620 1660 6630
rect 2250 6620 2540 6630
rect 3650 6620 3870 6630
rect 3990 6620 8510 6630
rect 8520 6620 9480 6630
rect 9540 6620 9610 6630
rect 9800 6620 9990 6630
rect 0 6610 1610 6620
rect 1670 6610 1720 6620
rect 1740 6610 1750 6620
rect 2240 6610 2540 6620
rect 3680 6610 3880 6620
rect 3990 6610 8500 6620
rect 8510 6610 9480 6620
rect 9560 6610 9610 6620
rect 9770 6610 9990 6620
rect 0 6600 1590 6610
rect 1640 6600 1750 6610
rect 2240 6600 2540 6610
rect 3690 6600 3890 6610
rect 3990 6600 6040 6610
rect 6050 6600 6070 6610
rect 6090 6600 8760 6610
rect 8780 6600 9480 6610
rect 9580 6600 9610 6610
rect 9730 6600 9990 6610
rect 0 6590 1580 6600
rect 1630 6590 1640 6600
rect 1670 6590 1740 6600
rect 2240 6590 2550 6600
rect 3730 6590 3900 6600
rect 3990 6590 6070 6600
rect 6090 6590 6220 6600
rect 6260 6590 6270 6600
rect 6300 6590 8760 6600
rect 8770 6590 9480 6600
rect 9590 6590 9610 6600
rect 9690 6590 9990 6600
rect 0 6580 1340 6590
rect 1350 6580 1470 6590
rect 1480 6580 1550 6590
rect 1650 6580 1750 6590
rect 2230 6580 2540 6590
rect 3740 6580 3910 6590
rect 4000 6580 5940 6590
rect 5950 6580 6060 6590
rect 6110 6580 6120 6590
rect 6130 6580 6210 6590
rect 6260 6580 6270 6590
rect 6320 6580 6340 6590
rect 6350 6580 8540 6590
rect 8570 6580 8690 6590
rect 8700 6580 8870 6590
rect 8890 6580 9480 6590
rect 9530 6580 9560 6590
rect 9680 6580 9990 6590
rect 0 6570 1350 6580
rect 1360 6570 1530 6580
rect 1640 6570 1760 6580
rect 2090 6570 2110 6580
rect 2210 6570 2540 6580
rect 3760 6570 3920 6580
rect 4010 6570 5940 6580
rect 5960 6570 6010 6580
rect 6020 6570 6050 6580
rect 6130 6570 6210 6580
rect 6360 6570 6380 6580
rect 6390 6570 8550 6580
rect 8560 6570 8600 6580
rect 8610 6570 8750 6580
rect 8760 6570 8870 6580
rect 8880 6570 9490 6580
rect 9530 6570 9570 6580
rect 9680 6570 9990 6580
rect 0 6560 1350 6570
rect 1380 6560 1490 6570
rect 1630 6560 1760 6570
rect 2090 6560 2150 6570
rect 2160 6560 2550 6570
rect 3770 6560 3920 6570
rect 4010 6560 5940 6570
rect 5970 6560 6000 6570
rect 6040 6560 6050 6570
rect 6070 6560 6090 6570
rect 6140 6560 6170 6570
rect 6410 6560 6430 6570
rect 6460 6560 6560 6570
rect 6580 6560 8750 6570
rect 8760 6560 9490 6570
rect 9520 6560 9580 6570
rect 9590 6560 9640 6570
rect 9680 6560 9990 6570
rect 0 6550 1350 6560
rect 1390 6550 1480 6560
rect 1750 6550 1770 6560
rect 2060 6550 2560 6560
rect 3790 6550 3930 6560
rect 4010 6550 5950 6560
rect 5980 6550 6000 6560
rect 6080 6550 6090 6560
rect 6130 6550 6140 6560
rect 6470 6550 6510 6560
rect 6600 6550 9490 6560
rect 9520 6550 9990 6560
rect 0 6540 1350 6550
rect 1400 6540 1450 6550
rect 1760 6540 1770 6550
rect 2060 6540 2570 6550
rect 3800 6540 3940 6550
rect 4020 6540 5950 6550
rect 5990 6540 6010 6550
rect 6080 6540 6100 6550
rect 6470 6540 6480 6550
rect 6610 6540 8020 6550
rect 8040 6540 8730 6550
rect 8750 6540 9500 6550
rect 9510 6540 9990 6550
rect 0 6530 1370 6540
rect 1760 6530 1770 6540
rect 2090 6530 2570 6540
rect 3830 6530 3950 6540
rect 4010 6530 5810 6540
rect 5820 6530 5960 6540
rect 6010 6530 6020 6540
rect 6090 6530 6110 6540
rect 6600 6530 6620 6540
rect 6670 6530 8720 6540
rect 8740 6530 9550 6540
rect 9560 6530 9990 6540
rect 0 6520 1330 6530
rect 2060 6520 2070 6530
rect 2090 6520 2220 6530
rect 2260 6520 2560 6530
rect 3850 6520 3950 6530
rect 4020 6520 5810 6530
rect 5830 6520 5840 6530
rect 5880 6520 5970 6530
rect 6090 6520 6120 6530
rect 6670 6520 8710 6530
rect 8740 6520 9420 6530
rect 9430 6520 9970 6530
rect 0 6510 1300 6520
rect 2090 6510 2230 6520
rect 2280 6510 2530 6520
rect 3870 6510 3960 6520
rect 4020 6510 5820 6520
rect 5840 6510 5850 6520
rect 5890 6510 5970 6520
rect 6090 6510 6100 6520
rect 6660 6510 8710 6520
rect 8730 6510 9190 6520
rect 9200 6510 9410 6520
rect 9440 6510 9940 6520
rect 0 6500 1270 6510
rect 1290 6500 1300 6510
rect 2100 6500 2240 6510
rect 2280 6500 2410 6510
rect 2440 6500 2490 6510
rect 3890 6500 3970 6510
rect 4030 6500 5800 6510
rect 5840 6500 5870 6510
rect 5890 6500 5940 6510
rect 5960 6500 5980 6510
rect 6660 6500 8020 6510
rect 8050 6500 8700 6510
rect 8720 6500 9410 6510
rect 9420 6500 9910 6510
rect 0 6490 1260 6500
rect 2120 6490 2250 6500
rect 2280 6490 2400 6500
rect 3900 6490 3980 6500
rect 4020 6490 5800 6500
rect 5860 6490 5930 6500
rect 6690 6490 8020 6500
rect 8050 6490 8690 6500
rect 8720 6490 9880 6500
rect 0 6480 1250 6490
rect 2140 6480 2260 6490
rect 2280 6480 2400 6490
rect 3920 6480 3980 6490
rect 4030 6480 5740 6490
rect 5750 6480 5760 6490
rect 5770 6480 5790 6490
rect 5800 6480 5810 6490
rect 5880 6480 5930 6490
rect 5990 6480 6000 6490
rect 6720 6480 8030 6490
rect 8050 6480 8690 6490
rect 8710 6480 9680 6490
rect 9690 6480 9850 6490
rect 0 6470 1240 6480
rect 2160 6470 2270 6480
rect 2290 6470 2400 6480
rect 3930 6470 3990 6480
rect 4030 6470 5770 6480
rect 5910 6470 5950 6480
rect 5960 6470 6010 6480
rect 6730 6470 8030 6480
rect 8040 6470 8680 6480
rect 8700 6470 9800 6480
rect 0 6460 1230 6470
rect 2170 6460 2200 6470
rect 2210 6460 2270 6470
rect 2290 6460 2390 6470
rect 2530 6460 2560 6470
rect 3950 6460 4000 6470
rect 4040 6460 5780 6470
rect 5820 6460 5840 6470
rect 5910 6460 6020 6470
rect 6730 6460 8680 6470
rect 8700 6460 9760 6470
rect 0 6450 1240 6460
rect 2170 6450 2220 6460
rect 2310 6450 2390 6460
rect 2520 6450 2560 6460
rect 3960 6450 4010 6460
rect 4040 6450 5720 6460
rect 5730 6450 5870 6460
rect 5910 6450 5950 6460
rect 6000 6450 6030 6460
rect 6750 6450 8670 6460
rect 8690 6450 9680 6460
rect 0 6440 1240 6450
rect 2160 6440 2250 6450
rect 2320 6440 2380 6450
rect 2520 6440 2540 6450
rect 3970 6440 4030 6450
rect 4040 6440 5680 6450
rect 5700 6440 5720 6450
rect 5790 6440 5810 6450
rect 5840 6440 5870 6450
rect 6000 6440 6030 6450
rect 6780 6440 8670 6450
rect 8680 6440 9680 6450
rect 0 6430 1220 6440
rect 1300 6430 1320 6440
rect 1330 6430 1350 6440
rect 1670 6430 1690 6440
rect 2150 6430 2280 6440
rect 2340 6430 2370 6440
rect 3990 6430 5680 6440
rect 6790 6430 8660 6440
rect 8680 6430 9580 6440
rect 9600 6430 9670 6440
rect 0 6420 1220 6430
rect 1300 6420 1320 6430
rect 1670 6420 1690 6430
rect 2140 6420 2310 6430
rect 2350 6420 2370 6430
rect 4000 6420 5690 6430
rect 6800 6420 8650 6430
rect 8670 6420 9580 6430
rect 9600 6420 9640 6430
rect 0 6410 1220 6420
rect 1230 6410 1250 6420
rect 1670 6410 1690 6420
rect 1750 6410 1800 6420
rect 2120 6410 2350 6420
rect 4020 6410 5690 6420
rect 5900 6410 5980 6420
rect 6810 6410 8650 6420
rect 8670 6410 9590 6420
rect 9600 6410 9630 6420
rect 0 6400 1200 6410
rect 1210 6400 1220 6410
rect 1650 6400 1820 6410
rect 2080 6400 2090 6410
rect 2110 6400 2380 6410
rect 4030 6400 5720 6410
rect 5840 6400 5990 6410
rect 6000 6400 6010 6410
rect 6830 6400 8640 6410
rect 8660 6400 9630 6410
rect 0 6390 1200 6400
rect 1220 6390 1230 6400
rect 1250 6390 1260 6400
rect 1300 6390 1330 6400
rect 1640 6390 1780 6400
rect 1810 6390 1830 6400
rect 2080 6390 2090 6400
rect 2100 6390 2390 6400
rect 4050 6390 5670 6400
rect 5700 6390 5870 6400
rect 6830 6390 8640 6400
rect 8660 6390 9630 6400
rect 0 6380 1230 6390
rect 1250 6380 1260 6390
rect 1340 6380 1400 6390
rect 1640 6380 1680 6390
rect 1700 6380 1730 6390
rect 1900 6380 1930 6390
rect 2090 6380 2390 6390
rect 4060 6380 5660 6390
rect 5720 6380 5840 6390
rect 6830 6380 8630 6390
rect 8650 6380 9630 6390
rect 0 6370 1210 6380
rect 1250 6370 1340 6380
rect 1360 6370 1390 6380
rect 1630 6370 1670 6380
rect 1890 6370 1950 6380
rect 2060 6370 2400 6380
rect 4070 6370 5650 6380
rect 5670 6370 5700 6380
rect 6820 6370 7500 6380
rect 7510 6370 8630 6380
rect 8650 6370 9610 6380
rect 0 6360 1220 6370
rect 1260 6360 1390 6370
rect 1620 6360 1670 6370
rect 1880 6360 1970 6370
rect 2020 6360 2400 6370
rect 4090 6360 5660 6370
rect 6290 6360 6300 6370
rect 6830 6360 8620 6370
rect 8640 6360 9480 6370
rect 9490 6360 9610 6370
rect 0 6350 1230 6360
rect 1270 6350 1400 6360
rect 1620 6350 1660 6360
rect 1880 6350 1970 6360
rect 2020 6350 2400 6360
rect 4100 6350 5660 6360
rect 5980 6350 6030 6360
rect 6270 6350 6340 6360
rect 6840 6350 8050 6360
rect 8060 6350 8620 6360
rect 8630 6350 9450 6360
rect 9490 6350 9630 6360
rect 0 6340 1240 6350
rect 1280 6340 1370 6350
rect 1380 6340 1400 6350
rect 1610 6340 1640 6350
rect 1850 6340 1970 6350
rect 2020 6340 2400 6350
rect 4110 6340 5570 6350
rect 5900 6340 6050 6350
rect 6080 6340 6350 6350
rect 6840 6340 8050 6350
rect 8070 6340 8610 6350
rect 8630 6340 9420 6350
rect 9430 6340 9450 6350
rect 9500 6340 9630 6350
rect 0 6330 1210 6340
rect 1220 6330 1260 6340
rect 1290 6330 1390 6340
rect 1610 6330 1630 6340
rect 1870 6330 1900 6340
rect 1910 6330 1970 6340
rect 2020 6330 2380 6340
rect 2460 6330 2470 6340
rect 4120 6330 5480 6340
rect 5690 6330 5700 6340
rect 5860 6330 6360 6340
rect 6850 6330 7590 6340
rect 7600 6330 8050 6340
rect 8060 6330 8610 6340
rect 8620 6330 9380 6340
rect 9420 6330 9460 6340
rect 9500 6330 9630 6340
rect 0 6320 1220 6330
rect 1250 6320 1270 6330
rect 1300 6320 1390 6330
rect 1900 6320 1970 6330
rect 2020 6320 2390 6330
rect 2460 6320 2470 6330
rect 4130 6320 5430 6330
rect 5850 6320 6370 6330
rect 6860 6320 7590 6330
rect 7610 6320 8600 6330
rect 8620 6320 9350 6330
rect 9380 6320 9400 6330
rect 9420 6320 9460 6330
rect 9510 6320 9640 6330
rect 0 6310 1200 6320
rect 1310 6310 1390 6320
rect 1890 6310 2010 6320
rect 2020 6310 2390 6320
rect 2460 6310 2470 6320
rect 4140 6310 5400 6320
rect 5840 6310 6400 6320
rect 6860 6310 7590 6320
rect 7610 6310 8600 6320
rect 8610 6310 9320 6320
rect 9380 6310 9390 6320
rect 9420 6310 9460 6320
rect 9510 6310 9590 6320
rect 9600 6310 9640 6320
rect 0 6300 1200 6310
rect 1240 6300 1250 6310
rect 1320 6300 1390 6310
rect 1880 6300 2400 6310
rect 4160 6300 5380 6310
rect 5840 6300 6420 6310
rect 6870 6300 7590 6310
rect 7610 6300 8590 6310
rect 8610 6300 9290 6310
rect 9370 6300 9400 6310
rect 9420 6300 9470 6310
rect 9510 6300 9590 6310
rect 9600 6300 9630 6310
rect 0 6290 1210 6300
rect 1290 6290 1300 6300
rect 1320 6290 1390 6300
rect 1860 6290 2400 6300
rect 2450 6290 2460 6300
rect 4170 6290 5360 6300
rect 5820 6290 6450 6300
rect 6840 6290 8580 6300
rect 8600 6290 9280 6300
rect 9350 6290 9400 6300
rect 9430 6290 9470 6300
rect 9500 6290 9590 6300
rect 9620 6290 9630 6300
rect 0 6280 1210 6290
rect 1330 6280 1390 6290
rect 1860 6280 2400 6290
rect 2450 6280 2460 6290
rect 4180 6280 5360 6290
rect 5710 6280 6460 6290
rect 6840 6280 7390 6290
rect 7400 6280 8580 6290
rect 8590 6280 9280 6290
rect 9330 6280 9400 6290
rect 9430 6280 9470 6290
rect 9510 6280 9640 6290
rect 0 6270 1200 6280
rect 1290 6270 1310 6280
rect 1330 6270 1390 6280
rect 1850 6270 2400 6280
rect 2450 6270 2460 6280
rect 4190 6270 5360 6280
rect 5690 6270 6460 6280
rect 6840 6270 8070 6280
rect 8080 6270 8570 6280
rect 8590 6270 9270 6280
rect 9330 6270 9400 6280
rect 9430 6270 9470 6280
rect 9520 6270 9640 6280
rect 0 6260 1200 6270
rect 1300 6260 1320 6270
rect 1340 6260 1390 6270
rect 1830 6260 2390 6270
rect 2450 6260 2460 6270
rect 4200 6260 5340 6270
rect 5680 6260 6470 6270
rect 6850 6260 7430 6270
rect 7450 6260 8070 6270
rect 8080 6260 8570 6270
rect 8590 6260 9270 6270
rect 9340 6260 9400 6270
rect 9430 6260 9480 6270
rect 9530 6260 9560 6270
rect 9620 6260 9640 6270
rect 9880 6260 9900 6270
rect 9960 6260 9980 6270
rect 0 6250 1200 6260
rect 1340 6250 1360 6260
rect 1370 6250 1390 6260
rect 1820 6250 2400 6260
rect 2450 6250 2460 6260
rect 4210 6250 5320 6260
rect 5650 6250 6480 6260
rect 6860 6250 7430 6260
rect 7440 6250 8070 6260
rect 8080 6250 8570 6260
rect 8590 6250 9260 6260
rect 9320 6250 9400 6260
rect 9440 6250 9480 6260
rect 9620 6250 9640 6260
rect 9880 6250 9900 6260
rect 9950 6250 9990 6260
rect 0 6240 1180 6250
rect 1390 6240 1400 6250
rect 1810 6240 2400 6250
rect 4220 6240 5310 6250
rect 5630 6240 6510 6250
rect 6870 6240 7620 6250
rect 7630 6240 8070 6250
rect 8090 6240 9250 6250
rect 9310 6240 9410 6250
rect 9440 6240 9490 6250
rect 9620 6240 9640 6250
rect 9820 6240 9870 6250
rect 9890 6240 9940 6250
rect 9950 6240 9990 6250
rect 0 6230 1180 6240
rect 1810 6230 2400 6240
rect 4230 6230 5300 6240
rect 5620 6230 6520 6240
rect 6880 6230 7450 6240
rect 7470 6230 8070 6240
rect 8080 6230 9250 6240
rect 9300 6230 9370 6240
rect 9380 6230 9410 6240
rect 9450 6230 9470 6240
rect 9820 6230 9940 6240
rect 9980 6230 9990 6240
rect 0 6220 1180 6230
rect 1800 6220 2400 6230
rect 4230 6220 5300 6230
rect 5600 6220 6540 6230
rect 6890 6220 8070 6230
rect 8080 6220 9240 6230
rect 9300 6220 9360 6230
rect 9380 6220 9410 6230
rect 9610 6220 9630 6230
rect 9650 6220 9660 6230
rect 9810 6220 9920 6230
rect 9940 6220 9980 6230
rect 9990 6220 9990 6230
rect 0 6210 1170 6220
rect 1800 6210 2400 6220
rect 4240 6210 5290 6220
rect 5590 6210 6550 6220
rect 6900 6210 8070 6220
rect 8090 6210 9240 6220
rect 9320 6210 9350 6220
rect 9610 6210 9630 6220
rect 9650 6210 9660 6220
rect 9810 6210 9900 6220
rect 9960 6210 9990 6220
rect 0 6200 1180 6210
rect 1790 6200 2400 6210
rect 4250 6200 5280 6210
rect 5570 6200 6550 6210
rect 6910 6200 7630 6210
rect 7650 6200 8070 6210
rect 8100 6200 9230 6210
rect 9290 6200 9300 6210
rect 9360 6200 9370 6210
rect 9610 6200 9670 6210
rect 9810 6200 9910 6210
rect 9930 6200 9940 6210
rect 9950 6200 9990 6210
rect 0 6190 1170 6200
rect 1790 6190 2400 6200
rect 4250 6190 5270 6200
rect 5300 6190 5310 6200
rect 5550 6190 6560 6200
rect 6920 6190 7630 6200
rect 7650 6190 9230 6200
rect 9280 6190 9300 6200
rect 9620 6190 9670 6200
rect 9820 6190 9990 6200
rect 0 6180 1170 6190
rect 1790 6180 2370 6190
rect 4260 6180 5260 6190
rect 5290 6180 5300 6190
rect 5540 6180 6570 6190
rect 6940 6180 7650 6190
rect 7660 6180 9210 6190
rect 9240 6180 9250 6190
rect 9280 6180 9290 6190
rect 9620 6180 9680 6190
rect 9820 6180 9940 6190
rect 9950 6180 9990 6190
rect 0 6170 1170 6180
rect 1220 6170 1240 6180
rect 1790 6170 2370 6180
rect 4270 6170 5250 6180
rect 5280 6170 5290 6180
rect 5510 6170 6610 6180
rect 6960 6170 7480 6180
rect 7500 6170 7650 6180
rect 7670 6170 9210 6180
rect 9260 6170 9280 6180
rect 9620 6170 9680 6180
rect 9830 6170 9930 6180
rect 9950 6170 9990 6180
rect 0 6160 1170 6170
rect 1180 6160 1210 6170
rect 1230 6160 1240 6170
rect 1790 6160 2380 6170
rect 4280 6160 5260 6170
rect 5270 6160 5280 6170
rect 5490 6160 6620 6170
rect 6960 6160 7480 6170
rect 7490 6160 7590 6170
rect 7610 6160 7650 6170
rect 7670 6160 9210 6170
rect 9230 6160 9240 6170
rect 9620 6160 9640 6170
rect 9830 6160 9940 6170
rect 9950 6160 9990 6170
rect 0 6150 1150 6160
rect 1160 6150 1170 6160
rect 1180 6150 1210 6160
rect 1230 6150 1240 6160
rect 1300 6150 1310 6160
rect 1780 6150 2380 6160
rect 4290 6150 5250 6160
rect 5260 6150 5280 6160
rect 5470 6150 5480 6160
rect 5490 6150 6630 6160
rect 6970 6150 7620 6160
rect 7630 6150 7650 6160
rect 7670 6150 7980 6160
rect 7990 6150 8110 6160
rect 8120 6150 9220 6160
rect 9830 6150 9940 6160
rect 9960 6150 9990 6160
rect 0 6140 1130 6150
rect 1170 6140 1210 6150
rect 1790 6140 2410 6150
rect 4290 6140 5240 6150
rect 5250 6140 5270 6150
rect 5470 6140 6640 6150
rect 6980 6140 7630 6150
rect 7670 6140 7910 6150
rect 7930 6140 8080 6150
rect 8120 6140 8510 6150
rect 8520 6140 9200 6150
rect 9840 6140 9940 6150
rect 9960 6140 9990 6150
rect 0 6130 1120 6140
rect 1160 6130 1220 6140
rect 1230 6130 1240 6140
rect 1690 6130 1720 6140
rect 1800 6130 2420 6140
rect 4300 6130 5220 6140
rect 5240 6130 5260 6140
rect 5470 6130 6630 6140
rect 6980 6130 7540 6140
rect 7580 6130 8510 6140
rect 8570 6130 9180 6140
rect 9840 6130 9920 6140
rect 9930 6130 9950 6140
rect 9970 6130 9990 6140
rect 0 6120 1110 6130
rect 1150 6120 1180 6130
rect 1190 6120 1210 6130
rect 1230 6120 1240 6130
rect 1680 6120 1730 6130
rect 1800 6120 2420 6130
rect 4300 6120 5220 6130
rect 5240 6120 5250 6130
rect 5450 6120 5460 6130
rect 5470 6120 6660 6130
rect 6990 6120 7550 6130
rect 7580 6120 7690 6130
rect 7700 6120 8510 6130
rect 8540 6120 9150 6130
rect 9850 6120 9900 6130
rect 9930 6120 9950 6130
rect 9970 6120 9990 6130
rect 0 6110 1170 6120
rect 1180 6110 1210 6120
rect 1240 6110 1250 6120
rect 1680 6110 1730 6120
rect 1810 6110 2430 6120
rect 4310 6110 5210 6120
rect 5230 6110 5250 6120
rect 5450 6110 6660 6120
rect 6990 6110 7520 6120
rect 7540 6110 7550 6120
rect 7560 6110 7680 6120
rect 7700 6110 8510 6120
rect 8540 6110 9120 6120
rect 9860 6110 9880 6120
rect 9920 6110 9950 6120
rect 9980 6110 9990 6120
rect 0 6100 1120 6110
rect 1180 6100 1190 6110
rect 1200 6100 1220 6110
rect 1240 6100 1250 6110
rect 1680 6100 1730 6110
rect 1810 6100 2430 6110
rect 3920 6100 3940 6110
rect 4310 6100 5200 6110
rect 5230 6100 5250 6110
rect 5430 6100 6670 6110
rect 6990 6100 7520 6110
rect 7550 6100 7680 6110
rect 7700 6100 8510 6110
rect 8540 6100 9090 6110
rect 9920 6100 9950 6110
rect 9980 6100 9990 6110
rect 0 6090 1120 6100
rect 1170 6090 1180 6100
rect 1210 6090 1230 6100
rect 1260 6090 1270 6100
rect 1690 6090 1740 6100
rect 1810 6090 2440 6100
rect 3900 6090 3950 6100
rect 4320 6090 5220 6100
rect 5230 6090 5240 6100
rect 5430 6090 6670 6100
rect 6990 6090 7540 6100
rect 7550 6090 9070 6100
rect 9390 6090 9470 6100
rect 9860 6090 9870 6100
rect 9980 6090 9990 6100
rect 0 6080 1110 6090
rect 1210 6080 1230 6090
rect 1700 6080 1740 6090
rect 1820 6080 2440 6090
rect 3890 6080 3960 6090
rect 4320 6080 5210 6090
rect 5230 6080 5240 6090
rect 5410 6080 6680 6090
rect 6990 6080 7610 6090
rect 7620 6080 9030 6090
rect 9360 6080 9480 6090
rect 9860 6080 9880 6090
rect 9970 6080 9990 6090
rect 0 6070 1110 6080
rect 1220 6070 1230 6080
rect 1820 6070 2440 6080
rect 3870 6070 3970 6080
rect 4330 6070 5200 6080
rect 5220 6070 5230 6080
rect 5410 6070 6680 6080
rect 7000 6070 7530 6080
rect 7540 6070 9000 6080
rect 9350 6070 9480 6080
rect 9860 6070 9890 6080
rect 9960 6070 9990 6080
rect 0 6060 810 6070
rect 820 6060 1010 6070
rect 1040 6060 1060 6070
rect 1110 6060 1150 6070
rect 1820 6060 2450 6070
rect 3850 6060 3980 6070
rect 4330 6060 5190 6070
rect 5210 6060 5230 6070
rect 5400 6060 6690 6070
rect 7000 6060 8960 6070
rect 9340 6060 9400 6070
rect 9450 6060 9490 6070
rect 9870 6060 9900 6070
rect 9950 6060 9990 6070
rect 0 6050 800 6060
rect 840 6050 850 6060
rect 860 6050 1060 6060
rect 1740 6050 1790 6060
rect 1820 6050 2450 6060
rect 3840 6050 3980 6060
rect 4340 6050 5180 6060
rect 5210 6050 5220 6060
rect 5400 6050 6700 6060
rect 6990 6050 7590 6060
rect 7600 6050 8930 6060
rect 9260 6050 9300 6060
rect 9350 6050 9390 6060
rect 9450 6050 9490 6060
rect 9870 6050 9930 6060
rect 9940 6050 9990 6060
rect 0 6040 780 6050
rect 860 6040 910 6050
rect 940 6040 1040 6050
rect 1070 6040 1100 6050
rect 1110 6040 1130 6050
rect 1740 6040 2460 6050
rect 3790 6040 3800 6050
rect 3820 6040 3990 6050
rect 4340 6040 5180 6050
rect 5200 6040 5210 6050
rect 5400 6040 6700 6050
rect 7000 6040 7510 6050
rect 7530 6040 7590 6050
rect 7600 6040 8910 6050
rect 9230 6040 9300 6050
rect 9350 6040 9390 6050
rect 9450 6040 9490 6050
rect 9870 6040 9930 6050
rect 9940 6040 9990 6050
rect 0 6030 770 6040
rect 1020 6030 1030 6040
rect 1060 6030 1080 6040
rect 1100 6030 1120 6040
rect 1750 6030 2470 6040
rect 3790 6030 4000 6040
rect 4340 6030 5200 6040
rect 5390 6030 6710 6040
rect 7000 6030 7500 6040
rect 7510 6030 7580 6040
rect 7590 6030 7630 6040
rect 7640 6030 8850 6040
rect 9190 6030 9300 6040
rect 9350 6030 9390 6040
rect 9440 6030 9480 6040
rect 9870 6030 9920 6040
rect 9940 6030 9990 6040
rect 0 6020 770 6030
rect 810 6020 820 6030
rect 1020 6020 1060 6030
rect 1100 6020 1110 6030
rect 1750 6020 2470 6030
rect 3790 6020 4010 6030
rect 4350 6020 5190 6030
rect 5390 6020 6720 6030
rect 7010 6020 8420 6030
rect 8440 6020 8820 6030
rect 9180 6020 9270 6030
rect 9350 6020 9390 6030
rect 9420 6020 9480 6030
rect 9870 6020 9910 6030
rect 9940 6020 9990 6030
rect 0 6010 760 6020
rect 790 6010 810 6020
rect 1060 6010 1090 6020
rect 1100 6010 1110 6020
rect 1750 6010 2480 6020
rect 3800 6010 4030 6020
rect 4350 6010 5180 6020
rect 5390 6010 6720 6020
rect 7010 6010 7400 6020
rect 7420 6010 7490 6020
rect 7500 6010 8420 6020
rect 8440 6010 8790 6020
rect 9180 6010 9240 6020
rect 9360 6010 9470 6020
rect 9880 6010 9900 6020
rect 9940 6010 9990 6020
rect 0 6000 750 6010
rect 780 6000 790 6010
rect 1030 6000 1070 6010
rect 1090 6000 1110 6010
rect 1770 6000 2490 6010
rect 3810 6000 3940 6010
rect 3950 6000 3960 6010
rect 3970 6000 4010 6010
rect 4020 6000 4040 6010
rect 4350 6000 5180 6010
rect 5390 6000 6720 6010
rect 7010 6000 7400 6010
rect 7420 6000 7490 6010
rect 7510 6000 7600 6010
rect 7610 6000 8420 6010
rect 8430 6000 8760 6010
rect 9110 6000 9140 6010
rect 9180 6000 9230 6010
rect 9360 6000 9450 6010
rect 9900 6000 9920 6010
rect 9950 6000 9990 6010
rect 0 5990 750 6000
rect 780 5990 790 6000
rect 970 5990 990 6000
rect 1010 5990 1050 6000
rect 1090 5990 1110 6000
rect 1810 5990 2490 6000
rect 3830 5990 4010 6000
rect 4020 5990 4060 6000
rect 4350 5990 5160 6000
rect 5380 5990 6720 6000
rect 7010 5990 7390 6000
rect 7410 5990 7470 6000
rect 7510 5990 7590 6000
rect 7610 5990 8410 6000
rect 8420 5990 8730 6000
rect 9100 5990 9140 6000
rect 9190 5990 9230 6000
rect 9360 5990 9450 6000
rect 9920 5990 9930 6000
rect 9960 5990 9990 6000
rect 0 5980 740 5990
rect 780 5980 790 5990
rect 990 5980 1100 5990
rect 1810 5980 2500 5990
rect 3780 5980 3820 5990
rect 3840 5980 4010 5990
rect 4020 5980 4070 5990
rect 4350 5980 5150 5990
rect 5380 5980 6730 5990
rect 7010 5980 7400 5990
rect 7410 5980 7470 5990
rect 7490 5980 7530 5990
rect 7550 5980 7590 5990
rect 7600 5980 7690 5990
rect 7720 5980 8330 5990
rect 8350 5980 8400 5990
rect 8420 5980 8700 5990
rect 9040 5980 9070 5990
rect 9100 5980 9150 5990
rect 9190 5980 9230 5990
rect 9360 5980 9470 5990
rect 9920 5980 9940 5990
rect 9950 5980 9960 5990
rect 9970 5980 9990 5990
rect 0 5970 740 5980
rect 770 5970 780 5980
rect 880 5970 900 5980
rect 1000 5970 1090 5980
rect 1160 5970 1180 5980
rect 1820 5970 2510 5980
rect 3780 5970 3840 5980
rect 3860 5970 3920 5980
rect 3930 5970 4090 5980
rect 4350 5970 5150 5980
rect 5370 5970 6730 5980
rect 7010 5970 7450 5980
rect 7470 5970 7500 5980
rect 7520 5970 7530 5980
rect 7550 5970 7580 5980
rect 7590 5970 7660 5980
rect 7690 5970 7720 5980
rect 7730 5970 8330 5980
rect 8350 5970 8400 5980
rect 8410 5970 8660 5980
rect 9030 5970 9080 5980
rect 9100 5970 9150 5980
rect 9190 5970 9230 5980
rect 9270 5970 9300 5980
rect 9370 5970 9410 5980
rect 9430 5970 9480 5980
rect 9890 5970 9990 5980
rect 0 5960 740 5970
rect 870 5960 910 5970
rect 1820 5960 1990 5970
rect 2010 5960 2490 5970
rect 2510 5960 2520 5970
rect 3780 5960 3850 5970
rect 3870 5960 3930 5970
rect 3950 5960 4100 5970
rect 4350 5960 4500 5970
rect 4530 5960 5150 5970
rect 5370 5960 6730 5970
rect 7000 5960 7280 5970
rect 7300 5960 7430 5970
rect 7460 5960 7510 5970
rect 7520 5960 7530 5970
rect 7550 5960 7650 5970
rect 7660 5960 7670 5970
rect 7680 5960 7700 5970
rect 7730 5960 8330 5970
rect 8350 5960 8360 5970
rect 8370 5960 8390 5970
rect 8410 5960 8620 5970
rect 8970 5960 9000 5970
rect 9030 5960 9090 5970
rect 9110 5960 9150 5970
rect 9200 5960 9310 5970
rect 9370 5960 9410 5970
rect 9440 5960 9490 5970
rect 9900 5960 9930 5970
rect 0 5950 730 5960
rect 860 5950 910 5960
rect 1820 5950 1990 5960
rect 2000 5950 2480 5960
rect 3770 5950 3860 5960
rect 3880 5950 4120 5960
rect 4350 5950 5160 5960
rect 5360 5950 6730 5960
rect 7000 5950 7530 5960
rect 7550 5950 7670 5960
rect 7680 5950 7700 5960
rect 7710 5950 8310 5960
rect 8350 5950 8360 5960
rect 8370 5950 8390 5960
rect 8400 5950 8590 5960
rect 8970 5950 9010 5960
rect 9030 5950 9090 5960
rect 9110 5950 9150 5960
rect 9200 5950 9300 5960
rect 9370 5950 9410 5960
rect 9450 5950 9500 5960
rect 9980 5950 9990 5960
rect 0 5940 720 5950
rect 860 5940 920 5950
rect 1810 5940 2480 5950
rect 3770 5940 3870 5950
rect 3890 5940 4140 5950
rect 4350 5940 5150 5950
rect 5360 5940 6730 5950
rect 7010 5940 7320 5950
rect 7330 5940 7490 5950
rect 7550 5940 8380 5950
rect 8400 5940 8560 5950
rect 8970 5940 9010 5950
rect 9030 5940 9100 5950
rect 9110 5940 9150 5950
rect 9200 5940 9280 5950
rect 9380 5940 9420 5950
rect 9460 5940 9510 5950
rect 9910 5940 9990 5950
rect 0 5930 700 5940
rect 850 5930 930 5940
rect 1790 5930 2470 5940
rect 3770 5930 3880 5940
rect 3900 5930 3940 5940
rect 3950 5930 4160 5940
rect 4340 5930 5150 5940
rect 5360 5930 6740 5940
rect 7010 5930 7310 5940
rect 7350 5930 8120 5940
rect 8150 5930 8370 5940
rect 8390 5930 8540 5940
rect 8860 5930 8900 5940
rect 8970 5930 9020 5940
rect 9030 5930 9150 5940
rect 9200 5930 9250 5940
rect 9380 5930 9420 5940
rect 9470 5930 9510 5940
rect 9900 5930 9960 5940
rect 9970 5930 9990 5940
rect 0 5920 700 5930
rect 840 5920 940 5930
rect 1780 5920 2460 5930
rect 3760 5920 3840 5930
rect 3860 5920 3890 5930
rect 3910 5920 4170 5930
rect 4340 5920 5140 5930
rect 5360 5920 6740 5930
rect 7010 5920 7310 5930
rect 7320 5920 7340 5930
rect 7360 5920 8090 5930
rect 8150 5920 8370 5930
rect 8380 5920 8510 5930
rect 8840 5920 8920 5930
rect 8980 5920 9020 5930
rect 9030 5920 9150 5930
rect 9210 5920 9250 5930
rect 9380 5920 9420 5930
rect 9900 5920 9960 5930
rect 9970 5920 9990 5930
rect 0 5910 680 5920
rect 830 5910 940 5920
rect 1760 5910 2390 5920
rect 2410 5910 2450 5920
rect 3770 5910 3840 5920
rect 3860 5910 3900 5920
rect 3920 5910 4200 5920
rect 4330 5910 5130 5920
rect 5360 5910 6750 5920
rect 7010 5910 8090 5920
rect 8150 5910 8370 5920
rect 8380 5910 8470 5920
rect 8820 5910 8930 5920
rect 8980 5910 9020 5920
rect 9030 5910 9150 5920
rect 9210 5910 9250 5920
rect 9380 5910 9420 5920
rect 9910 5910 9990 5920
rect 0 5900 670 5910
rect 830 5900 920 5910
rect 1760 5900 1830 5910
rect 1860 5900 2360 5910
rect 3770 5900 3860 5910
rect 3870 5900 3910 5910
rect 3930 5900 4010 5910
rect 4020 5900 4210 5910
rect 4310 5900 5120 5910
rect 5350 5900 6760 5910
rect 7010 5900 7300 5910
rect 7320 5900 8090 5910
rect 8150 5900 8250 5910
rect 8260 5900 8350 5910
rect 8370 5900 8440 5910
rect 8810 5900 8940 5910
rect 8980 5900 9070 5910
rect 9080 5900 9160 5910
rect 9210 5900 9250 5910
rect 9390 5900 9420 5910
rect 9910 5900 9990 5910
rect 0 5890 650 5900
rect 830 5890 920 5900
rect 1860 5890 2350 5900
rect 3780 5890 3920 5900
rect 3930 5890 4010 5900
rect 4020 5890 4230 5900
rect 4290 5890 5120 5900
rect 5350 5890 6760 5900
rect 7020 5890 7290 5900
rect 7330 5890 7360 5900
rect 7390 5890 8090 5900
rect 8160 5890 8350 5900
rect 8360 5890 8410 5900
rect 8730 5890 8750 5900
rect 8810 5890 8850 5900
rect 8900 5890 8940 5900
rect 8990 5890 9070 5900
rect 9080 5890 9160 5900
rect 9210 5890 9260 5900
rect 9290 5890 9340 5900
rect 9910 5890 9990 5900
rect 0 5880 640 5890
rect 820 5880 930 5890
rect 1870 5880 2340 5890
rect 3760 5880 3880 5890
rect 3890 5880 3920 5890
rect 3940 5880 4010 5890
rect 4030 5880 5120 5890
rect 5350 5880 6760 5890
rect 7020 5880 7300 5890
rect 7330 5880 7350 5890
rect 7370 5880 7380 5890
rect 7390 5880 8030 5890
rect 8040 5880 8090 5890
rect 8160 5880 8370 5890
rect 8700 5880 8760 5890
rect 8800 5880 8840 5890
rect 8910 5880 8950 5890
rect 8990 5880 9070 5890
rect 9090 5880 9160 5890
rect 9220 5880 9340 5890
rect 9920 5880 9990 5890
rect 0 5870 390 5880
rect 400 5870 640 5880
rect 800 5870 870 5880
rect 880 5870 940 5880
rect 1870 5870 2330 5880
rect 3760 5870 3890 5880
rect 3900 5870 3930 5880
rect 3940 5870 4020 5880
rect 4030 5870 5110 5880
rect 5350 5870 6760 5880
rect 7020 5870 7330 5880
rect 7340 5870 7350 5880
rect 7360 5870 7380 5880
rect 7390 5870 7930 5880
rect 7950 5870 8030 5880
rect 8040 5870 8090 5880
rect 8160 5870 8340 5880
rect 8670 5870 8750 5880
rect 8800 5870 8840 5880
rect 8910 5870 8950 5880
rect 8990 5870 9070 5880
rect 9100 5870 9160 5880
rect 9220 5870 9330 5880
rect 9920 5870 9990 5880
rect 0 5860 370 5870
rect 380 5860 590 5870
rect 600 5860 650 5870
rect 900 5860 960 5870
rect 1870 5860 2300 5870
rect 3760 5860 3770 5870
rect 3780 5860 3820 5870
rect 3860 5860 3880 5870
rect 3890 5860 3930 5870
rect 3950 5860 5110 5870
rect 5350 5860 6770 5870
rect 7020 5860 7370 5870
rect 7400 5860 7910 5870
rect 7980 5860 7990 5870
rect 8010 5860 8090 5870
rect 8160 5860 8310 5870
rect 8630 5860 8730 5870
rect 8800 5860 8840 5870
rect 8910 5860 8950 5870
rect 9000 5860 9070 5870
rect 9100 5860 9160 5870
rect 9220 5860 9300 5870
rect 9930 5860 9990 5870
rect 0 5850 340 5860
rect 380 5850 590 5860
rect 610 5850 630 5860
rect 890 5850 960 5860
rect 1870 5850 2290 5860
rect 3770 5850 3800 5860
rect 3810 5850 3820 5860
rect 3840 5850 3860 5860
rect 3880 5850 3940 5860
rect 3950 5850 5110 5860
rect 5350 5850 6770 5860
rect 7020 5850 7880 5860
rect 7970 5850 8000 5860
rect 8010 5850 8090 5860
rect 8160 5850 8260 5860
rect 8620 5850 8710 5860
rect 8800 5850 8840 5860
rect 8920 5850 8950 5860
rect 9000 5850 9070 5860
rect 9110 5850 9160 5860
rect 9230 5850 9270 5860
rect 9930 5850 9990 5860
rect 0 5840 580 5850
rect 930 5840 970 5850
rect 1880 5840 2280 5850
rect 3760 5840 3790 5850
rect 3830 5840 3860 5850
rect 3870 5840 3940 5850
rect 3960 5840 5100 5850
rect 5350 5840 6770 5850
rect 7020 5840 7870 5850
rect 7970 5840 8090 5850
rect 8160 5840 8240 5850
rect 8620 5840 8710 5850
rect 8800 5840 8840 5850
rect 8920 5840 8960 5850
rect 9010 5840 9070 5850
rect 9110 5840 9170 5850
rect 9920 5840 9970 5850
rect 0 5830 580 5840
rect 1880 5830 2270 5840
rect 2460 5830 2490 5840
rect 3770 5830 3790 5840
rect 3870 5830 3940 5840
rect 3960 5830 4590 5840
rect 4610 5830 5100 5840
rect 5350 5830 6780 5840
rect 7000 5830 7010 5840
rect 7020 5830 7880 5840
rect 7980 5830 8090 5840
rect 8130 5830 8220 5840
rect 8680 5830 8720 5840
rect 8810 5830 8840 5840
rect 8920 5830 8960 5840
rect 9010 5830 9070 5840
rect 9120 5830 9160 5840
rect 9930 5830 9960 5840
rect 9990 5830 9990 5840
rect 0 5820 570 5830
rect 1880 5820 2270 5830
rect 2430 5820 2490 5830
rect 3150 5820 3170 5830
rect 3750 5820 3760 5830
rect 3770 5820 3800 5830
rect 3880 5820 3940 5830
rect 3970 5820 4570 5830
rect 4610 5820 5100 5830
rect 5350 5820 6780 5830
rect 7000 5820 7890 5830
rect 8000 5820 8100 5830
rect 8110 5820 8200 5830
rect 8680 5820 8720 5830
rect 8810 5820 8850 5830
rect 8920 5820 8960 5830
rect 9010 5820 9070 5830
rect 9130 5820 9160 5830
rect 9970 5820 9990 5830
rect 0 5810 560 5820
rect 750 5810 810 5820
rect 1890 5810 2250 5820
rect 2420 5810 2490 5820
rect 3130 5810 3170 5820
rect 3780 5810 3800 5820
rect 3850 5810 3860 5820
rect 3870 5810 3940 5820
rect 3970 5810 4570 5820
rect 4620 5810 5100 5820
rect 5350 5810 6790 5820
rect 7000 5810 7860 5820
rect 7870 5810 7880 5820
rect 8010 5810 8160 5820
rect 8680 5810 8720 5820
rect 8810 5810 8850 5820
rect 8930 5810 8960 5820
rect 9020 5810 9060 5820
rect 9960 5810 9990 5820
rect 0 5800 550 5810
rect 630 5800 650 5810
rect 740 5800 800 5810
rect 850 5800 880 5810
rect 1890 5800 2250 5810
rect 2420 5800 2490 5810
rect 3110 5800 3160 5810
rect 3850 5800 3900 5810
rect 3910 5800 3950 5810
rect 3970 5800 4580 5810
rect 4620 5800 5090 5810
rect 5350 5800 6790 5810
rect 7010 5800 7830 5810
rect 7850 5800 7870 5810
rect 7930 5800 7940 5810
rect 8020 5800 8120 5810
rect 8690 5800 8720 5810
rect 8810 5800 8850 5810
rect 8920 5800 8960 5810
rect 9020 5800 9060 5810
rect 9950 5800 9990 5810
rect 0 5790 550 5800
rect 740 5790 800 5800
rect 830 5790 880 5800
rect 1890 5790 1900 5800
rect 1930 5790 2240 5800
rect 2410 5790 2480 5800
rect 3080 5790 3160 5800
rect 3930 5790 3960 5800
rect 3970 5790 4050 5800
rect 4070 5790 4580 5800
rect 4620 5790 5090 5800
rect 5340 5790 6790 5800
rect 7010 5790 7750 5800
rect 7790 5790 7870 5800
rect 7920 5790 7940 5800
rect 8000 5790 8100 5800
rect 8690 5790 8730 5800
rect 8820 5790 8860 5800
rect 8920 5790 8960 5800
rect 9030 5790 9060 5800
rect 9940 5790 9990 5800
rect 0 5780 550 5790
rect 720 5780 790 5790
rect 820 5780 880 5790
rect 1950 5780 2230 5790
rect 2390 5780 2470 5790
rect 2480 5780 2490 5790
rect 3110 5780 3170 5790
rect 3890 5780 3900 5790
rect 3930 5780 3960 5790
rect 3980 5780 4060 5790
rect 4080 5780 4480 5790
rect 4490 5780 4560 5790
rect 4620 5780 5090 5790
rect 5340 5780 6800 5790
rect 7010 5780 7740 5790
rect 7790 5780 8050 5790
rect 8390 5780 8420 5790
rect 8690 5780 8730 5790
rect 8820 5780 8860 5790
rect 8910 5780 8950 5790
rect 9940 5780 9990 5790
rect 0 5770 550 5780
rect 610 5770 630 5780
rect 720 5770 780 5780
rect 830 5770 840 5780
rect 1950 5770 2220 5780
rect 2350 5770 2370 5780
rect 2400 5770 2470 5780
rect 3120 5770 3180 5780
rect 3880 5770 3960 5780
rect 3980 5770 4070 5780
rect 4080 5770 4560 5780
rect 4610 5770 4680 5780
rect 4720 5770 4740 5780
rect 4750 5770 5090 5780
rect 5340 5770 6800 5780
rect 7010 5770 7750 5780
rect 7770 5770 8010 5780
rect 8390 5770 8420 5780
rect 8690 5770 8730 5780
rect 8820 5770 8950 5780
rect 9950 5770 9990 5780
rect 0 5760 540 5770
rect 580 5760 640 5770
rect 710 5760 770 5770
rect 830 5760 840 5770
rect 1960 5760 2210 5770
rect 2350 5760 2370 5770
rect 2390 5760 2400 5770
rect 2410 5760 2450 5770
rect 3050 5760 3100 5770
rect 3120 5760 3180 5770
rect 3900 5760 3920 5770
rect 3930 5760 3950 5770
rect 3960 5760 3970 5770
rect 3980 5760 4090 5770
rect 4100 5760 4510 5770
rect 4520 5760 4540 5770
rect 4600 5760 4680 5770
rect 4710 5760 4740 5770
rect 4750 5760 5090 5770
rect 5340 5760 6790 5770
rect 7010 5760 7980 5770
rect 8390 5760 8420 5770
rect 8700 5760 8730 5770
rect 8830 5760 8940 5770
rect 9950 5760 9990 5770
rect 0 5750 540 5760
rect 580 5750 640 5760
rect 710 5750 770 5760
rect 820 5750 850 5760
rect 1960 5750 2210 5760
rect 2340 5750 2350 5760
rect 3040 5750 3180 5760
rect 3930 5750 3970 5760
rect 3990 5750 4500 5760
rect 4520 5750 4550 5760
rect 4560 5750 4580 5760
rect 4600 5750 4640 5760
rect 4650 5750 4670 5760
rect 4680 5750 4750 5760
rect 4770 5750 5080 5760
rect 5330 5750 6790 5760
rect 7000 5750 7920 5760
rect 8390 5750 8420 5760
rect 8700 5750 8730 5760
rect 8850 5750 8920 5760
rect 9950 5750 9990 5760
rect 0 5740 530 5750
rect 540 5740 610 5750
rect 750 5740 770 5750
rect 830 5740 860 5750
rect 1960 5740 2200 5750
rect 2320 5740 2340 5750
rect 3030 5740 3180 5750
rect 3930 5740 3950 5750
rect 4000 5740 4350 5750
rect 4370 5740 4500 5750
rect 4560 5740 4590 5750
rect 4600 5740 4750 5750
rect 4770 5740 5080 5750
rect 5330 5740 6800 5750
rect 7000 5740 7920 5750
rect 8250 5740 8270 5750
rect 8390 5740 8430 5750
rect 8700 5740 8740 5750
rect 8880 5740 8890 5750
rect 9960 5740 9990 5750
rect 0 5730 590 5740
rect 1960 5730 2200 5740
rect 2330 5730 2340 5740
rect 3010 5730 3180 5740
rect 3950 5730 3960 5740
rect 4010 5730 4350 5740
rect 4360 5730 4520 5740
rect 4530 5730 4580 5740
rect 4600 5730 5080 5740
rect 5320 5730 6810 5740
rect 6990 5730 7850 5740
rect 7870 5730 7890 5740
rect 8250 5730 8280 5740
rect 8390 5730 8430 5740
rect 8700 5730 8740 5740
rect 9960 5730 9990 5740
rect 0 5720 560 5730
rect 700 5720 730 5730
rect 1960 5720 2200 5730
rect 2330 5720 2350 5730
rect 3000 5720 3030 5730
rect 3050 5720 3180 5730
rect 3780 5720 3810 5730
rect 4020 5720 4290 5730
rect 4300 5720 4340 5730
rect 4350 5720 4380 5730
rect 4410 5720 4520 5730
rect 4530 5720 4590 5730
rect 4610 5720 5080 5730
rect 5320 5720 6810 5730
rect 6990 5720 7790 5730
rect 8190 5720 8210 5730
rect 8250 5720 8280 5730
rect 8400 5720 8430 5730
rect 8700 5720 8740 5730
rect 9960 5720 9990 5730
rect 0 5710 490 5720
rect 550 5710 630 5720
rect 670 5710 780 5720
rect 1950 5710 2190 5720
rect 2310 5710 2350 5720
rect 3010 5710 3020 5720
rect 3040 5710 3190 5720
rect 3800 5710 3820 5720
rect 4010 5710 4280 5720
rect 4310 5710 4400 5720
rect 4410 5710 4560 5720
rect 4660 5710 4760 5720
rect 4770 5710 5070 5720
rect 5320 5710 6820 5720
rect 6990 5710 7610 5720
rect 7640 5710 7750 5720
rect 8180 5710 8220 5720
rect 8250 5710 8280 5720
rect 8400 5710 8430 5720
rect 8710 5710 8750 5720
rect 9960 5710 9990 5720
rect 0 5700 460 5710
rect 510 5700 630 5710
rect 670 5700 790 5710
rect 1960 5700 2190 5710
rect 2300 5700 2330 5710
rect 3030 5700 3180 5710
rect 4010 5700 4040 5710
rect 4060 5700 4230 5710
rect 4250 5700 4290 5710
rect 4300 5700 4320 5710
rect 4340 5700 4550 5710
rect 4580 5700 4600 5710
rect 4630 5700 4640 5710
rect 4660 5700 4710 5710
rect 4730 5700 4760 5710
rect 4790 5700 5070 5710
rect 5310 5700 6820 5710
rect 6990 5700 7730 5710
rect 8120 5700 8140 5710
rect 8180 5700 8220 5710
rect 8250 5700 8290 5710
rect 8400 5700 8440 5710
rect 8710 5700 8740 5710
rect 9970 5700 9990 5710
rect 0 5690 550 5700
rect 560 5690 630 5700
rect 670 5690 800 5700
rect 1960 5690 1970 5700
rect 1980 5690 2190 5700
rect 2290 5690 2330 5700
rect 2840 5690 2880 5700
rect 2900 5690 2920 5700
rect 3020 5690 3180 5700
rect 4010 5690 4260 5700
rect 4280 5690 4320 5700
rect 4340 5690 4550 5700
rect 4570 5690 4600 5700
rect 4630 5690 4680 5700
rect 4760 5690 4770 5700
rect 4800 5690 5070 5700
rect 5310 5690 6820 5700
rect 6990 5690 7700 5700
rect 8120 5690 8150 5700
rect 8190 5690 8220 5700
rect 8250 5690 8290 5700
rect 8400 5690 8440 5700
rect 0 5680 550 5690
rect 560 5680 620 5690
rect 650 5680 790 5690
rect 1090 5680 1100 5690
rect 1990 5680 2180 5690
rect 2290 5680 2320 5690
rect 2840 5680 2920 5690
rect 3020 5680 3180 5690
rect 3800 5680 3810 5690
rect 4000 5680 4190 5690
rect 4200 5680 4250 5690
rect 4270 5680 4300 5690
rect 4310 5680 4570 5690
rect 4640 5680 4710 5690
rect 4760 5680 4790 5690
rect 4800 5680 5070 5690
rect 5300 5680 6820 5690
rect 7000 5680 7670 5690
rect 7710 5680 7720 5690
rect 8120 5680 8150 5690
rect 8190 5680 8220 5690
rect 8250 5680 8290 5690
rect 8410 5680 8440 5690
rect 0 5670 540 5680
rect 550 5670 630 5680
rect 650 5670 790 5680
rect 1980 5670 2180 5680
rect 2280 5670 2300 5680
rect 2380 5670 2390 5680
rect 2820 5670 2910 5680
rect 2950 5670 2960 5680
rect 3010 5670 3150 5680
rect 3170 5670 3180 5680
rect 4000 5670 4180 5680
rect 4200 5670 4290 5680
rect 4310 5670 4360 5680
rect 4370 5670 4410 5680
rect 4420 5670 4580 5680
rect 4600 5670 4610 5680
rect 4630 5670 4710 5680
rect 4720 5670 4740 5680
rect 4770 5670 5070 5680
rect 5300 5670 6830 5680
rect 6990 5670 7650 5680
rect 7660 5670 7690 5680
rect 8030 5670 8060 5680
rect 8120 5670 8150 5680
rect 8190 5670 8230 5680
rect 8260 5670 8290 5680
rect 8410 5670 8440 5680
rect 0 5660 620 5670
rect 650 5660 780 5670
rect 1980 5660 2170 5670
rect 2280 5660 2300 5670
rect 2380 5660 2390 5670
rect 2820 5660 2910 5670
rect 2960 5660 2970 5670
rect 3010 5660 3150 5670
rect 3190 5660 3200 5670
rect 3740 5660 3760 5670
rect 3900 5660 3910 5670
rect 3990 5660 4220 5670
rect 4240 5660 4280 5670
rect 4320 5660 4350 5670
rect 4360 5660 4390 5670
rect 4420 5660 4580 5670
rect 4600 5660 4750 5670
rect 4780 5660 5070 5670
rect 5300 5660 6830 5670
rect 6990 5660 7660 5670
rect 8030 5660 8060 5670
rect 8120 5660 8160 5670
rect 8190 5660 8230 5670
rect 8260 5660 8290 5670
rect 8410 5660 8450 5670
rect 0 5650 610 5660
rect 660 5650 760 5660
rect 1980 5650 2170 5660
rect 2270 5650 2290 5660
rect 2360 5650 2420 5660
rect 2820 5650 2970 5660
rect 3010 5650 3160 5660
rect 3700 5650 3710 5660
rect 3800 5650 3810 5660
rect 3880 5650 3900 5660
rect 3990 5650 4210 5660
rect 4240 5650 4280 5660
rect 4300 5650 4330 5660
rect 4340 5650 4400 5660
rect 4410 5650 4580 5660
rect 4600 5650 4720 5660
rect 4780 5650 5070 5660
rect 5100 5650 5130 5660
rect 5300 5650 5710 5660
rect 5730 5650 6830 5660
rect 6960 5650 6980 5660
rect 7000 5650 7580 5660
rect 7600 5650 7630 5660
rect 8030 5650 8070 5660
rect 8120 5650 8160 5660
rect 8190 5650 8230 5660
rect 8260 5650 8290 5660
rect 8410 5650 8450 5660
rect 8480 5650 8530 5660
rect 0 5640 530 5650
rect 570 5640 610 5650
rect 660 5640 760 5650
rect 1970 5640 2160 5650
rect 2270 5640 2290 5650
rect 2350 5640 2400 5650
rect 2820 5640 2980 5650
rect 3010 5640 3170 5650
rect 3790 5640 3800 5650
rect 3880 5640 3900 5650
rect 3940 5640 4210 5650
rect 4240 5640 4270 5650
rect 4280 5640 4330 5650
rect 4340 5640 4730 5650
rect 4750 5640 5070 5650
rect 5100 5640 5120 5650
rect 5290 5640 5600 5650
rect 5770 5640 6840 5650
rect 6980 5640 7570 5650
rect 8030 5640 8070 5650
rect 8120 5640 8160 5650
rect 8190 5640 8230 5650
rect 8260 5640 8300 5650
rect 8410 5640 8530 5650
rect 9990 5640 9990 5650
rect 0 5630 520 5640
rect 660 5630 750 5640
rect 1970 5630 2110 5640
rect 2140 5630 2150 5640
rect 2260 5630 2290 5640
rect 2350 5630 2440 5640
rect 2830 5630 3170 5640
rect 3720 5630 3730 5640
rect 3820 5630 3840 5640
rect 3870 5630 3900 5640
rect 3920 5630 4090 5640
rect 4100 5630 4200 5640
rect 4230 5630 4260 5640
rect 4290 5630 5080 5640
rect 5100 5630 5120 5640
rect 5290 5630 5550 5640
rect 5790 5630 5840 5640
rect 5860 5630 6840 5640
rect 6990 5630 7510 5640
rect 8030 5630 8070 5640
rect 8130 5630 8160 5640
rect 8200 5630 8230 5640
rect 8260 5630 8300 5640
rect 8410 5630 8520 5640
rect 9990 5630 9990 5640
rect 0 5620 520 5630
rect 660 5620 730 5630
rect 2000 5620 2030 5630
rect 2050 5620 2090 5630
rect 2260 5620 2280 5630
rect 2350 5620 2420 5630
rect 2850 5620 3170 5630
rect 3800 5620 3810 5630
rect 3820 5620 3840 5630
rect 3860 5620 3900 5630
rect 3910 5620 4090 5630
rect 4100 5620 4190 5630
rect 4230 5620 4260 5630
rect 4290 5620 5080 5630
rect 5100 5620 5110 5630
rect 5290 5620 5540 5630
rect 5870 5620 5940 5630
rect 5950 5620 6850 5630
rect 6990 5620 7460 5630
rect 7480 5620 7490 5630
rect 8040 5620 8070 5630
rect 8120 5620 8170 5630
rect 8200 5620 8230 5630
rect 8270 5620 8300 5630
rect 8420 5620 8500 5630
rect 9990 5620 9990 5630
rect 0 5610 520 5620
rect 670 5610 720 5620
rect 2010 5610 2020 5620
rect 2060 5610 2110 5620
rect 2260 5610 2270 5620
rect 2350 5610 2420 5620
rect 2880 5610 3160 5620
rect 3800 5610 4120 5620
rect 4130 5610 4190 5620
rect 4220 5610 5070 5620
rect 5090 5610 5110 5620
rect 5290 5610 5510 5620
rect 5880 5610 5890 5620
rect 5960 5610 5990 5620
rect 6060 5610 6200 5620
rect 6270 5610 6280 5620
rect 6290 5610 6320 5620
rect 6430 5610 6440 5620
rect 6450 5610 6850 5620
rect 6980 5610 7440 5620
rect 7820 5610 7900 5620
rect 8040 5610 8070 5620
rect 8080 5610 8170 5620
rect 8200 5610 8240 5620
rect 8270 5610 8300 5620
rect 8360 5610 8390 5620
rect 8420 5610 8460 5620
rect 0 5600 510 5610
rect 670 5600 700 5610
rect 2030 5600 2040 5610
rect 2050 5600 2110 5610
rect 2350 5600 2410 5610
rect 2890 5600 2910 5610
rect 2940 5600 3170 5610
rect 3800 5600 4190 5610
rect 4210 5600 4260 5610
rect 4290 5600 5110 5610
rect 5290 5600 5480 5610
rect 5490 5600 5500 5610
rect 6070 5600 6170 5610
rect 6530 5600 6860 5610
rect 6980 5600 7430 5610
rect 7800 5600 7910 5610
rect 8040 5600 8170 5610
rect 8200 5600 8240 5610
rect 8270 5600 8310 5610
rect 8330 5600 8390 5610
rect 0 5590 510 5600
rect 560 5590 570 5600
rect 620 5590 630 5600
rect 680 5590 690 5600
rect 2050 5590 2080 5600
rect 2090 5590 2110 5600
rect 2350 5590 2380 5600
rect 2390 5590 2400 5600
rect 2940 5590 3160 5600
rect 3670 5590 3700 5600
rect 3780 5590 3870 5600
rect 3880 5590 4100 5600
rect 4110 5590 4150 5600
rect 4170 5590 4180 5600
rect 4210 5590 4310 5600
rect 4330 5590 5100 5600
rect 5280 5590 5470 5600
rect 6090 5590 6150 5600
rect 6610 5590 6860 5600
rect 6980 5590 7300 5600
rect 7320 5590 7420 5600
rect 7790 5590 7920 5600
rect 8040 5590 8170 5600
rect 8210 5590 8240 5600
rect 8280 5590 8390 5600
rect 8990 5590 9070 5600
rect 0 5580 510 5590
rect 620 5580 630 5590
rect 2090 5580 2100 5590
rect 2340 5580 2380 5590
rect 2950 5580 3160 5590
rect 3680 5580 3700 5590
rect 3780 5580 3820 5590
rect 3830 5580 3860 5590
rect 3870 5580 4110 5590
rect 4130 5580 4150 5590
rect 4210 5580 4240 5590
rect 4250 5580 4290 5590
rect 4320 5580 5090 5590
rect 5280 5580 5460 5590
rect 6090 5580 6110 5590
rect 6120 5580 6130 5590
rect 6620 5580 6870 5590
rect 6980 5580 7300 5590
rect 7320 5580 7400 5590
rect 7730 5580 7750 5590
rect 7790 5580 7840 5590
rect 7880 5580 7920 5590
rect 8040 5580 8100 5590
rect 8140 5580 8180 5590
rect 8210 5580 8250 5590
rect 8280 5580 8370 5590
rect 8970 5580 9080 5590
rect 0 5570 510 5580
rect 610 5570 630 5580
rect 2100 5570 2110 5580
rect 2340 5570 2380 5580
rect 2960 5570 3160 5580
rect 3440 5570 3450 5580
rect 3780 5570 3810 5580
rect 3820 5570 3850 5580
rect 3870 5570 4100 5580
rect 4120 5570 4160 5580
rect 4220 5570 4240 5580
rect 4280 5570 5090 5580
rect 5280 5570 5460 5580
rect 6620 5570 6870 5580
rect 6980 5570 7290 5580
rect 7320 5570 7360 5580
rect 7690 5570 7760 5580
rect 7790 5570 7830 5580
rect 7880 5570 7920 5580
rect 8050 5570 8080 5580
rect 8140 5570 8180 5580
rect 8210 5570 8250 5580
rect 8280 5570 8330 5580
rect 8970 5570 9090 5580
rect 0 5560 510 5570
rect 610 5560 650 5570
rect 2340 5560 2360 5570
rect 2980 5560 3170 5570
rect 3450 5560 3460 5570
rect 3780 5560 3840 5570
rect 3850 5560 4100 5570
rect 4120 5560 4160 5570
rect 4170 5560 4190 5570
rect 4300 5560 4490 5570
rect 4500 5560 5090 5570
rect 5280 5560 5450 5570
rect 6670 5560 6880 5570
rect 6970 5560 7300 5570
rect 7310 5560 7360 5570
rect 7670 5560 7760 5570
rect 7790 5560 7830 5570
rect 7890 5560 7930 5570
rect 8050 5560 8080 5570
rect 8140 5560 8180 5570
rect 8210 5560 8250 5570
rect 8960 5560 9010 5570
rect 9050 5560 9090 5570
rect 0 5550 500 5560
rect 610 5550 650 5560
rect 2100 5550 2110 5560
rect 2350 5550 2370 5560
rect 2990 5550 3170 5560
rect 3460 5550 3480 5560
rect 3730 5550 3740 5560
rect 3750 5550 3760 5560
rect 3800 5550 3830 5560
rect 3840 5550 3910 5560
rect 3920 5550 4100 5560
rect 4170 5550 4190 5560
rect 4270 5550 4280 5560
rect 4300 5550 4330 5560
rect 4350 5550 4370 5560
rect 4380 5550 4480 5560
rect 4500 5550 5090 5560
rect 5270 5550 5450 5560
rect 6670 5550 6880 5560
rect 6970 5550 7260 5560
rect 7300 5550 7320 5560
rect 7330 5550 7370 5560
rect 7660 5550 7740 5560
rect 7800 5550 7830 5560
rect 7890 5550 7930 5560
rect 8050 5550 8090 5560
rect 8140 5550 8180 5560
rect 8220 5550 8240 5560
rect 8870 5550 8900 5560
rect 8960 5550 9000 5560
rect 0 5540 510 5550
rect 610 5540 620 5550
rect 630 5540 650 5550
rect 2990 5540 3160 5550
rect 3470 5540 3490 5550
rect 3680 5540 3710 5550
rect 3730 5540 3740 5550
rect 3790 5540 3810 5550
rect 3830 5540 4100 5550
rect 4160 5540 4190 5550
rect 4210 5540 4230 5550
rect 4250 5540 4280 5550
rect 4300 5540 4330 5550
rect 4340 5540 4350 5550
rect 4370 5540 5090 5550
rect 5270 5540 5430 5550
rect 6080 5540 6090 5550
rect 6670 5540 6880 5550
rect 6960 5540 7260 5550
rect 7280 5540 7300 5550
rect 7330 5540 7370 5550
rect 7650 5540 7710 5550
rect 7800 5540 7830 5550
rect 7890 5540 7930 5550
rect 8050 5540 8090 5550
rect 8150 5540 8180 5550
rect 8870 5540 8900 5550
rect 8950 5540 8990 5550
rect 0 5530 500 5540
rect 630 5530 640 5540
rect 3030 5530 3160 5540
rect 3490 5530 3500 5540
rect 3670 5530 3710 5540
rect 3740 5530 3760 5540
rect 3780 5530 3800 5540
rect 3810 5530 4110 5540
rect 4160 5530 4180 5540
rect 4210 5530 4260 5540
rect 4270 5530 4290 5540
rect 4310 5530 4350 5540
rect 4360 5530 5090 5540
rect 5270 5530 5420 5540
rect 6680 5530 6880 5540
rect 6980 5530 7290 5540
rect 7340 5530 7370 5540
rect 7560 5530 7600 5540
rect 7660 5530 7700 5540
rect 7800 5530 7840 5540
rect 7890 5530 7930 5540
rect 8060 5530 8090 5540
rect 8150 5530 8180 5540
rect 8870 5530 8910 5540
rect 8950 5530 8990 5540
rect 0 5520 500 5530
rect 600 5520 610 5530
rect 940 5520 960 5530
rect 3050 5520 3160 5530
rect 3670 5520 3710 5530
rect 3740 5520 3750 5530
rect 3760 5520 3790 5530
rect 3800 5520 4130 5530
rect 4220 5520 4250 5530
rect 4280 5520 4350 5530
rect 4370 5520 5110 5530
rect 5270 5520 5410 5530
rect 6050 5520 6100 5530
rect 6710 5520 6880 5530
rect 6970 5520 7290 5530
rect 7340 5520 7350 5530
rect 7360 5520 7370 5530
rect 7530 5520 7620 5530
rect 7660 5520 7700 5530
rect 7800 5520 7840 5530
rect 7890 5520 7930 5530
rect 8060 5520 8090 5530
rect 8770 5520 8810 5530
rect 8870 5520 8910 5530
rect 8950 5520 8990 5530
rect 0 5510 460 5520
rect 600 5510 610 5520
rect 3060 5510 3160 5520
rect 3660 5510 3710 5520
rect 3740 5510 3770 5520
rect 3790 5510 4130 5520
rect 4260 5510 4300 5520
rect 4330 5510 4360 5520
rect 4370 5510 5100 5520
rect 5260 5510 5410 5520
rect 6050 5510 6110 5520
rect 6730 5510 6890 5520
rect 6970 5510 7250 5520
rect 7270 5510 7350 5520
rect 7360 5510 7380 5520
rect 7510 5510 7630 5520
rect 7660 5510 7700 5520
rect 7810 5510 7840 5520
rect 7900 5510 7930 5520
rect 8060 5510 8090 5520
rect 8760 5510 8820 5520
rect 8870 5510 8910 5520
rect 8960 5510 8990 5520
rect 9080 5510 9110 5520
rect 0 5500 350 5510
rect 600 5500 610 5510
rect 3060 5500 3150 5510
rect 3670 5500 3700 5510
rect 3730 5500 3740 5510
rect 3770 5500 4090 5510
rect 4120 5500 4140 5510
rect 4180 5500 4200 5510
rect 4210 5500 4230 5510
rect 4240 5500 4300 5510
rect 4330 5500 4360 5510
rect 4390 5500 4430 5510
rect 4460 5500 5100 5510
rect 5260 5500 5410 5510
rect 6040 5500 6120 5510
rect 6730 5500 6890 5510
rect 6970 5500 7230 5510
rect 7280 5500 7380 5510
rect 7510 5500 7630 5510
rect 7660 5500 7700 5510
rect 7730 5500 7740 5510
rect 7810 5500 7840 5510
rect 7900 5500 7940 5510
rect 8060 5500 8090 5510
rect 8690 5500 8720 5510
rect 8760 5500 8830 5510
rect 8870 5500 8910 5510
rect 8960 5500 9000 5510
rect 9050 5500 9110 5510
rect 0 5490 370 5500
rect 3070 5490 3140 5500
rect 3690 5490 3710 5500
rect 3750 5490 4090 5500
rect 4100 5490 4110 5500
rect 4150 5490 4190 5500
rect 4200 5490 4220 5500
rect 4250 5490 4360 5500
rect 4380 5490 4430 5500
rect 4460 5490 5100 5500
rect 5260 5490 5410 5500
rect 6020 5490 6120 5500
rect 6730 5490 6900 5500
rect 6960 5490 7220 5500
rect 7280 5490 7300 5500
rect 7340 5490 7380 5500
rect 7510 5490 7550 5500
rect 7590 5490 7630 5500
rect 7660 5490 7750 5500
rect 7810 5490 7850 5500
rect 7890 5490 7940 5500
rect 8690 5490 8730 5500
rect 8770 5490 8840 5500
rect 8880 5490 8920 5500
rect 8960 5490 9000 5500
rect 9050 5490 9120 5500
rect 0 5480 400 5490
rect 950 5480 960 5490
rect 3080 5480 3130 5490
rect 3660 5480 4000 5490
rect 4010 5480 4080 5490
rect 4140 5480 4180 5490
rect 4190 5480 4430 5490
rect 4470 5480 4500 5490
rect 4510 5480 5100 5490
rect 5260 5480 5410 5490
rect 6000 5480 6010 5490
rect 6020 5480 6120 5490
rect 6730 5480 6900 5490
rect 6970 5480 7230 5490
rect 7340 5480 7380 5490
rect 7510 5480 7550 5490
rect 7600 5480 7630 5490
rect 7660 5480 7750 5490
rect 7810 5480 7850 5490
rect 7890 5480 7930 5490
rect 8620 5480 8650 5490
rect 8690 5480 8730 5490
rect 8770 5480 8850 5490
rect 8880 5480 8920 5490
rect 8960 5480 9000 5490
rect 9050 5480 9120 5490
rect 0 5470 430 5480
rect 3080 5470 3110 5480
rect 3660 5470 4050 5480
rect 4070 5470 4080 5480
rect 4130 5470 4160 5480
rect 4190 5470 4250 5480
rect 4260 5470 4270 5480
rect 4320 5470 4440 5480
rect 4470 5470 4610 5480
rect 4620 5470 5090 5480
rect 5250 5470 5400 5480
rect 6000 5470 6120 5480
rect 6730 5470 6900 5480
rect 6970 5470 7230 5480
rect 7240 5470 7250 5480
rect 7340 5470 7380 5480
rect 7510 5470 7550 5480
rect 7590 5470 7630 5480
rect 7670 5470 7740 5480
rect 7810 5470 7850 5480
rect 7880 5470 7930 5480
rect 8620 5470 8660 5480
rect 8700 5470 8730 5480
rect 8770 5470 8860 5480
rect 8880 5470 8920 5480
rect 8970 5470 9000 5480
rect 9080 5470 9120 5480
rect 0 5460 440 5470
rect 3600 5460 4080 5470
rect 4120 5460 4150 5470
rect 4160 5460 4180 5470
rect 4190 5460 4270 5470
rect 4380 5460 4450 5470
rect 4460 5460 4490 5470
rect 4520 5460 4530 5470
rect 4550 5460 4570 5470
rect 4590 5460 4620 5470
rect 4630 5460 4700 5470
rect 4720 5460 5080 5470
rect 5250 5460 5400 5470
rect 5990 5460 6130 5470
rect 6740 5460 6900 5470
rect 6960 5460 7230 5470
rect 7290 5460 7300 5470
rect 7340 5460 7370 5470
rect 7510 5460 7550 5470
rect 7570 5460 7620 5470
rect 7670 5460 7710 5470
rect 7820 5460 7920 5470
rect 8620 5460 8660 5470
rect 8700 5460 8730 5470
rect 8770 5460 8870 5470
rect 8890 5460 8920 5470
rect 8970 5460 9010 5470
rect 9080 5460 9120 5470
rect 0 5450 440 5460
rect 540 5450 580 5460
rect 3600 5450 4080 5460
rect 4150 5450 4270 5460
rect 4290 5450 4300 5460
rect 4340 5450 4350 5460
rect 4380 5450 4480 5460
rect 4520 5450 4580 5460
rect 4590 5450 4660 5460
rect 4750 5450 5100 5460
rect 5250 5450 5400 5460
rect 5990 5450 6130 5460
rect 6730 5450 6900 5460
rect 6960 5450 7200 5460
rect 7210 5450 7220 5460
rect 7290 5450 7300 5460
rect 7350 5450 7360 5460
rect 7520 5450 7610 5460
rect 7670 5450 7710 5460
rect 7820 5450 7910 5460
rect 8520 5450 8560 5460
rect 8620 5450 8660 5460
rect 8700 5450 8740 5460
rect 8780 5450 8810 5460
rect 8830 5450 8870 5460
rect 8890 5450 8930 5460
rect 8970 5450 9010 5460
rect 9080 5450 9120 5460
rect 0 5440 440 5450
rect 530 5440 580 5450
rect 3590 5440 4070 5450
rect 4080 5440 4100 5450
rect 4120 5440 4270 5450
rect 4310 5440 4320 5450
rect 4340 5440 4350 5450
rect 4360 5440 4370 5450
rect 4420 5440 4470 5450
rect 4520 5440 4550 5450
rect 4590 5440 4620 5450
rect 4630 5440 4650 5450
rect 4660 5440 4670 5450
rect 4700 5440 4710 5450
rect 4730 5440 5100 5450
rect 5250 5440 5400 5450
rect 5990 5440 6130 5450
rect 6730 5440 6900 5450
rect 6950 5440 7190 5450
rect 7290 5440 7300 5450
rect 7520 5440 7600 5450
rect 7670 5440 7710 5450
rect 7820 5440 7900 5450
rect 8520 5440 8570 5450
rect 8630 5440 8660 5450
rect 8700 5440 8740 5450
rect 8780 5440 8820 5450
rect 8830 5440 8880 5450
rect 8890 5440 8930 5450
rect 8970 5440 9020 5450
rect 9070 5440 9110 5450
rect 0 5430 440 5440
rect 520 5430 570 5440
rect 3590 5430 4100 5440
rect 4110 5430 4330 5440
rect 4340 5430 4400 5440
rect 4410 5430 4460 5440
rect 4520 5430 4550 5440
rect 4580 5430 4600 5440
rect 4630 5430 4700 5440
rect 4720 5430 4740 5440
rect 4760 5430 5080 5440
rect 5240 5430 5400 5440
rect 5980 5430 6130 5440
rect 6730 5430 6900 5440
rect 6950 5430 7180 5440
rect 7290 5430 7300 5440
rect 7520 5430 7600 5440
rect 7680 5430 7710 5440
rect 7750 5430 7790 5440
rect 7820 5430 7870 5440
rect 8520 5430 8580 5440
rect 8630 5430 8670 5440
rect 8700 5430 8740 5440
rect 8780 5430 8820 5440
rect 8840 5430 8930 5440
rect 8980 5430 9110 5440
rect 0 5420 440 5430
rect 510 5420 570 5430
rect 3590 5420 4090 5430
rect 4110 5420 4320 5430
rect 4350 5420 4470 5430
rect 4550 5420 4570 5430
rect 4590 5420 4610 5430
rect 4630 5420 4670 5430
rect 4710 5420 4730 5430
rect 4780 5420 5090 5430
rect 5240 5420 5420 5430
rect 5980 5420 6130 5430
rect 6730 5420 6900 5430
rect 6960 5420 7180 5430
rect 7210 5420 7230 5430
rect 7290 5420 7300 5430
rect 7520 5420 7610 5430
rect 7680 5420 7790 5430
rect 8410 5420 8460 5430
rect 8520 5420 8590 5430
rect 8630 5420 8670 5430
rect 8710 5420 8750 5430
rect 8780 5420 8820 5430
rect 8850 5420 8930 5430
rect 8990 5420 9100 5430
rect 9560 5420 9580 5430
rect 0 5410 440 5420
rect 500 5410 560 5420
rect 3590 5410 4090 5420
rect 4100 5410 4310 5420
rect 4340 5410 4400 5420
rect 4410 5410 4460 5420
rect 4470 5410 4480 5420
rect 4520 5410 4570 5420
rect 4600 5410 4630 5420
rect 4660 5410 4680 5420
rect 4770 5410 5080 5420
rect 5240 5410 5410 5420
rect 5970 5410 6130 5420
rect 6720 5410 6900 5420
rect 6970 5410 7180 5420
rect 7200 5410 7240 5420
rect 7290 5410 7300 5420
rect 7520 5410 7560 5420
rect 7570 5410 7620 5420
rect 7680 5410 7790 5420
rect 8380 5410 8480 5420
rect 8520 5410 8600 5420
rect 8630 5410 8670 5420
rect 8710 5410 8750 5420
rect 8790 5410 8830 5420
rect 8860 5410 8940 5420
rect 8990 5410 9080 5420
rect 9550 5410 9580 5420
rect 0 5400 410 5410
rect 500 5400 560 5410
rect 3590 5400 4090 5410
rect 4100 5400 4230 5410
rect 4240 5400 4460 5410
rect 4470 5400 4500 5410
rect 4540 5400 4560 5410
rect 4580 5400 4590 5410
rect 4610 5400 4620 5410
rect 4750 5400 5090 5410
rect 5240 5400 5400 5410
rect 5970 5400 6130 5410
rect 6720 5400 6900 5410
rect 6970 5400 7190 5410
rect 7200 5400 7240 5410
rect 7290 5400 7300 5410
rect 7530 5400 7560 5410
rect 7580 5400 7630 5410
rect 7680 5400 7770 5410
rect 8360 5400 8480 5410
rect 8530 5400 8610 5410
rect 8640 5400 8670 5410
rect 8710 5400 8750 5410
rect 8790 5400 8830 5410
rect 8870 5400 8940 5410
rect 9010 5400 9060 5410
rect 9480 5400 9510 5410
rect 9550 5400 9580 5410
rect 0 5390 400 5400
rect 520 5390 560 5400
rect 3580 5390 4090 5400
rect 4100 5390 4220 5400
rect 4240 5390 4410 5400
rect 4440 5390 4450 5400
rect 4460 5390 4500 5400
rect 4520 5390 4530 5400
rect 4540 5390 4560 5400
rect 4590 5390 4600 5400
rect 4630 5390 4650 5400
rect 4750 5390 5080 5400
rect 5240 5390 5380 5400
rect 5970 5390 6130 5400
rect 6720 5390 6900 5400
rect 6930 5390 7190 5400
rect 7210 5390 7240 5400
rect 7290 5390 7300 5400
rect 7530 5390 7560 5400
rect 7590 5390 7640 5400
rect 7690 5390 7730 5400
rect 8350 5390 8420 5400
rect 8440 5390 8490 5400
rect 8530 5390 8620 5400
rect 8640 5390 8680 5400
rect 8710 5390 8750 5400
rect 8790 5390 8830 5400
rect 8880 5390 8940 5400
rect 9490 5390 9520 5400
rect 9550 5390 9580 5400
rect 0 5380 380 5390
rect 500 5380 540 5390
rect 3580 5380 3800 5390
rect 3810 5380 4080 5390
rect 4100 5380 4470 5390
rect 4480 5380 4490 5390
rect 4510 5380 4530 5390
rect 4540 5380 4560 5390
rect 4620 5380 4640 5390
rect 4650 5380 4680 5390
rect 4710 5380 5080 5390
rect 5240 5380 5370 5390
rect 5970 5380 6130 5390
rect 6730 5380 6910 5390
rect 6940 5380 7200 5390
rect 7210 5380 7240 5390
rect 7530 5380 7570 5390
rect 7600 5380 7650 5390
rect 8350 5380 8390 5390
rect 8450 5380 8490 5390
rect 8530 5380 8570 5390
rect 8580 5380 8630 5390
rect 8640 5380 8680 5390
rect 8720 5380 8760 5390
rect 8800 5380 8830 5390
rect 8890 5380 8940 5390
rect 9410 5380 9440 5390
rect 9490 5380 9530 5390
rect 9550 5380 9580 5390
rect 0 5370 360 5380
rect 450 5370 490 5380
rect 3580 5370 3800 5380
rect 3820 5370 4080 5380
rect 4100 5370 4180 5380
rect 4190 5370 4460 5380
rect 4490 5370 4530 5380
rect 4540 5370 4560 5380
rect 4590 5370 4620 5380
rect 4630 5370 4660 5380
rect 4700 5370 5080 5380
rect 5240 5370 5380 5380
rect 5970 5370 6130 5380
rect 6740 5370 6910 5380
rect 6950 5370 7220 5380
rect 7280 5370 7290 5380
rect 7530 5370 7570 5380
rect 7610 5370 7650 5380
rect 8240 5370 8270 5380
rect 8350 5370 8390 5380
rect 8460 5370 8490 5380
rect 8530 5370 8570 5380
rect 8590 5370 8640 5380
rect 8650 5370 8680 5380
rect 8720 5370 8760 5380
rect 8800 5370 8840 5380
rect 8900 5370 8940 5380
rect 9410 5370 9440 5380
rect 9500 5370 9570 5380
rect 0 5360 330 5370
rect 3570 5360 4080 5370
rect 4100 5360 4170 5370
rect 4190 5360 4440 5370
rect 4460 5360 4520 5370
rect 4540 5360 4650 5370
rect 4700 5360 5080 5370
rect 5240 5360 5380 5370
rect 5970 5360 6140 5370
rect 6760 5360 6910 5370
rect 6950 5360 7220 5370
rect 7280 5360 7290 5370
rect 7530 5360 7570 5370
rect 7620 5360 7630 5370
rect 8230 5360 8280 5370
rect 8360 5360 8390 5370
rect 8450 5360 8490 5370
rect 8530 5360 8570 5370
rect 8600 5360 8680 5370
rect 8720 5360 8760 5370
rect 8800 5360 8840 5370
rect 9410 5360 9440 5370
rect 9510 5360 9570 5370
rect 0 5350 300 5360
rect 3570 5350 3880 5360
rect 3890 5350 4080 5360
rect 4120 5350 4160 5360
rect 4190 5350 4470 5360
rect 4490 5350 4510 5360
rect 4520 5350 4640 5360
rect 4690 5350 4720 5360
rect 4730 5350 5090 5360
rect 5230 5350 5370 5360
rect 5970 5350 6140 5360
rect 6760 5350 6910 5360
rect 6950 5350 7250 5360
rect 7270 5350 7290 5360
rect 7530 5350 7570 5360
rect 8230 5350 8280 5360
rect 8360 5350 8400 5360
rect 8440 5350 8490 5360
rect 8540 5350 8580 5360
rect 8610 5350 8690 5360
rect 8730 5350 8760 5360
rect 8800 5350 8840 5360
rect 9290 5350 9360 5360
rect 9420 5350 9450 5360
rect 9520 5350 9570 5360
rect 0 5340 260 5350
rect 3570 5340 4080 5350
rect 4140 5340 4490 5350
rect 4510 5340 4570 5350
rect 4580 5340 4620 5350
rect 4700 5340 4720 5350
rect 4730 5340 5080 5350
rect 5230 5340 5360 5350
rect 5520 5340 5570 5350
rect 5960 5340 6150 5350
rect 6750 5340 6910 5350
rect 6940 5340 7250 5350
rect 7270 5340 7280 5350
rect 7540 5340 7560 5350
rect 8140 5340 8160 5350
rect 8230 5340 8290 5350
rect 8360 5340 8400 5350
rect 8410 5340 8480 5350
rect 8540 5340 8580 5350
rect 8620 5340 8690 5350
rect 8730 5340 8770 5350
rect 8810 5340 8830 5350
rect 9280 5340 9370 5350
rect 9420 5340 9450 5350
rect 9530 5340 9570 5350
rect 0 5330 250 5340
rect 3560 5330 4100 5340
rect 4140 5330 4450 5340
rect 4460 5330 4490 5340
rect 4510 5330 4560 5340
rect 4690 5330 4720 5340
rect 4730 5330 4750 5340
rect 4780 5330 5080 5340
rect 5230 5330 5350 5340
rect 5410 5330 5460 5340
rect 5510 5330 5600 5340
rect 5940 5330 6150 5340
rect 6760 5330 6910 5340
rect 6940 5330 7280 5340
rect 8130 5330 8170 5340
rect 8230 5330 8290 5340
rect 8360 5330 8470 5340
rect 8540 5330 8580 5340
rect 8620 5330 8690 5340
rect 8730 5330 8770 5340
rect 9270 5330 9320 5340
rect 9350 5330 9370 5340
rect 9420 5330 9450 5340
rect 9530 5330 9580 5340
rect 0 5320 240 5330
rect 3560 5320 4110 5330
rect 4140 5320 4500 5330
rect 4520 5320 4580 5330
rect 4600 5320 4630 5330
rect 4680 5320 4710 5330
rect 4730 5320 4750 5330
rect 4760 5320 5090 5330
rect 5230 5320 5460 5330
rect 5500 5320 5640 5330
rect 5940 5320 6150 5330
rect 6780 5320 6910 5330
rect 6950 5320 7270 5330
rect 8070 5320 8100 5330
rect 8130 5320 8170 5330
rect 8230 5320 8300 5330
rect 8370 5320 8460 5330
rect 8550 5320 8580 5330
rect 8630 5320 8690 5330
rect 8730 5320 8760 5330
rect 9270 5320 9300 5330
rect 9430 5320 9450 5330
rect 9530 5320 9590 5330
rect 0 5310 230 5320
rect 3550 5310 4110 5320
rect 4130 5310 4570 5320
rect 4610 5310 4640 5320
rect 4680 5310 4700 5320
rect 4730 5310 4760 5320
rect 4770 5310 5080 5320
rect 5230 5310 5670 5320
rect 5930 5310 6150 5320
rect 6800 5310 6920 5320
rect 6940 5310 7260 5320
rect 8060 5310 8110 5320
rect 8130 5310 8170 5320
rect 8230 5310 8310 5320
rect 8370 5310 8470 5320
rect 8550 5310 8580 5320
rect 8640 5310 8690 5320
rect 9260 5310 9300 5320
rect 9430 5310 9460 5320
rect 9530 5310 9600 5320
rect 0 5300 210 5310
rect 3550 5300 4600 5310
rect 4620 5300 4660 5310
rect 4720 5300 5090 5310
rect 5110 5300 5120 5310
rect 5230 5300 5680 5310
rect 5930 5300 6160 5310
rect 6810 5300 6910 5310
rect 6930 5300 7230 5310
rect 7240 5300 7260 5310
rect 8010 5300 8030 5310
rect 8060 5300 8120 5310
rect 8130 5300 8170 5310
rect 8230 5300 8310 5310
rect 8370 5300 8410 5310
rect 8430 5300 8470 5310
rect 8550 5300 8590 5310
rect 8650 5300 8690 5310
rect 9130 5300 9150 5310
rect 9270 5300 9300 5310
rect 9430 5300 9460 5310
rect 9530 5300 9560 5310
rect 9570 5300 9610 5310
rect 0 5290 200 5300
rect 3540 5290 4690 5300
rect 4710 5290 4740 5300
rect 4750 5290 5080 5300
rect 5230 5290 5590 5300
rect 5650 5290 5660 5300
rect 5920 5290 6160 5300
rect 6550 5290 6590 5300
rect 6800 5290 7250 5300
rect 8000 5290 8040 5300
rect 8060 5290 8120 5300
rect 8140 5290 8170 5300
rect 8230 5290 8310 5300
rect 8380 5290 8410 5300
rect 8440 5290 8490 5300
rect 8550 5290 8590 5300
rect 9130 5290 9160 5300
rect 9270 5290 9370 5300
rect 9430 5290 9460 5300
rect 9530 5290 9560 5300
rect 9580 5290 9620 5300
rect 9950 5290 9970 5300
rect 0 5280 190 5290
rect 3540 5280 4660 5290
rect 4670 5280 4710 5290
rect 4750 5280 5070 5290
rect 5230 5280 5580 5290
rect 5920 5280 6170 5290
rect 6500 5280 6590 5290
rect 6790 5280 6910 5290
rect 6920 5280 7240 5290
rect 8000 5280 8040 5290
rect 8060 5280 8130 5290
rect 8140 5280 8180 5290
rect 8230 5280 8260 5290
rect 8280 5280 8320 5290
rect 8380 5280 8410 5290
rect 8450 5280 8500 5290
rect 8550 5280 8590 5290
rect 9050 5280 9070 5290
rect 9130 5280 9160 5290
rect 9280 5280 9380 5290
rect 9440 5280 9470 5290
rect 9520 5280 9550 5290
rect 9590 5280 9610 5290
rect 9950 5280 9970 5290
rect 0 5270 180 5280
rect 3530 5270 4710 5280
rect 4780 5270 5090 5280
rect 5220 5270 5490 5280
rect 5500 5270 5570 5280
rect 5910 5270 6170 5280
rect 6470 5270 6580 5280
rect 6680 5270 6750 5280
rect 6800 5270 6910 5280
rect 6930 5270 7230 5280
rect 8010 5270 8050 5280
rect 8060 5270 8130 5280
rect 8140 5270 8180 5280
rect 8230 5270 8270 5280
rect 8290 5270 8330 5280
rect 8380 5270 8420 5280
rect 8460 5270 8510 5280
rect 8560 5270 8580 5280
rect 9040 5270 9080 5280
rect 9130 5270 9170 5280
rect 9290 5270 9330 5280
rect 9360 5270 9390 5280
rect 9440 5270 9470 5280
rect 9520 5270 9550 5280
rect 9950 5270 9980 5280
rect 0 5260 180 5270
rect 3530 5260 4710 5270
rect 4720 5260 4740 5270
rect 4760 5260 5070 5270
rect 5220 5260 5480 5270
rect 5880 5260 6170 5270
rect 6470 5260 6500 5270
rect 6640 5260 6780 5270
rect 6800 5260 6910 5270
rect 6930 5260 7230 5270
rect 7250 5260 7260 5270
rect 8010 5260 8050 5270
rect 8060 5260 8180 5270
rect 8230 5260 8260 5270
rect 8290 5260 8330 5270
rect 8380 5260 8420 5270
rect 8470 5260 8510 5270
rect 9040 5260 9090 5270
rect 9140 5260 9170 5270
rect 9370 5260 9390 5270
rect 9440 5260 9470 5270
rect 9850 5260 9880 5270
rect 9950 5260 9980 5270
rect 0 5250 170 5260
rect 3520 5250 4710 5260
rect 4720 5250 4740 5260
rect 4760 5250 5070 5260
rect 5220 5250 5520 5260
rect 5850 5250 6180 5260
rect 6620 5250 7230 5260
rect 7240 5250 7260 5260
rect 8010 5250 8050 5260
rect 8060 5250 8180 5260
rect 8230 5250 8260 5260
rect 8290 5250 8340 5260
rect 8380 5250 8420 5260
rect 8480 5250 8510 5260
rect 8940 5250 8970 5260
rect 9050 5250 9100 5260
rect 9140 5250 9170 5260
rect 9370 5250 9390 5260
rect 9440 5250 9470 5260
rect 9850 5250 9890 5260
rect 9960 5250 9980 5260
rect 0 5240 150 5250
rect 3520 5240 4710 5250
rect 4740 5240 5060 5250
rect 5230 5240 5560 5250
rect 5820 5240 6180 5250
rect 6630 5240 7260 5250
rect 8020 5240 8180 5250
rect 8230 5240 8340 5250
rect 8390 5240 8420 5250
rect 8940 5240 8980 5250
rect 9050 5240 9120 5250
rect 9140 5240 9170 5250
rect 9360 5240 9390 5250
rect 9450 5240 9470 5250
rect 9760 5240 9800 5250
rect 9850 5240 9910 5250
rect 9960 5240 9980 5250
rect 0 5230 140 5240
rect 3510 5230 4670 5240
rect 4680 5230 4720 5240
rect 4740 5230 5060 5240
rect 5230 5230 5600 5240
rect 5790 5230 6180 5240
rect 6610 5230 7270 5240
rect 8020 5230 8100 5240
rect 8110 5230 8180 5240
rect 8230 5230 8350 5240
rect 8390 5230 8420 5240
rect 8940 5230 8980 5240
rect 9050 5230 9130 5240
rect 9150 5230 9180 5240
rect 9290 5230 9320 5240
rect 9350 5230 9390 5240
rect 9730 5230 9820 5240
rect 9860 5230 9920 5240
rect 9970 5230 9990 5240
rect 0 5220 120 5230
rect 3510 5220 4740 5230
rect 4780 5220 5060 5230
rect 5230 5220 5670 5230
rect 5720 5220 6180 5230
rect 6600 5220 7270 5230
rect 7290 5220 7300 5230
rect 8020 5220 8100 5230
rect 8110 5220 8180 5230
rect 8230 5220 8300 5230
rect 8310 5220 8350 5230
rect 8400 5220 8410 5230
rect 8840 5220 8870 5230
rect 8940 5220 8990 5230
rect 9060 5220 9090 5230
rect 9100 5220 9140 5230
rect 9150 5220 9180 5230
rect 9290 5220 9380 5230
rect 9720 5220 9820 5230
rect 9860 5220 9930 5230
rect 9970 5220 9990 5230
rect 0 5210 100 5220
rect 2570 5210 2610 5220
rect 3500 5210 4770 5220
rect 4780 5210 5060 5220
rect 5230 5210 6180 5220
rect 6270 5210 6330 5220
rect 6580 5210 7190 5220
rect 8030 5210 8100 5220
rect 8120 5210 8180 5220
rect 8230 5210 8270 5220
rect 8320 5210 8350 5220
rect 8840 5210 8870 5220
rect 8940 5210 8990 5220
rect 9060 5210 9090 5220
rect 9110 5210 9180 5220
rect 9300 5210 9370 5220
rect 9720 5210 9750 5220
rect 9800 5210 9830 5220
rect 9870 5210 9900 5220
rect 9910 5210 9940 5220
rect 0 5200 90 5210
rect 2570 5200 2620 5210
rect 2650 5200 2660 5210
rect 3500 5200 5060 5210
rect 5230 5200 6190 5210
rect 6270 5200 6350 5210
rect 6560 5200 7140 5210
rect 7160 5200 7180 5210
rect 8030 5200 8100 5210
rect 8120 5200 8180 5210
rect 8230 5200 8260 5210
rect 8320 5200 8340 5210
rect 8760 5200 8780 5210
rect 8840 5200 8870 5210
rect 8940 5200 9000 5210
rect 9060 5200 9090 5210
rect 9120 5200 9180 5210
rect 9710 5200 9750 5210
rect 9800 5200 9830 5210
rect 9870 5200 9900 5210
rect 9930 5200 9950 5210
rect 9980 5200 9990 5210
rect 0 5190 70 5200
rect 2560 5190 2660 5200
rect 3490 5190 5060 5200
rect 5230 5190 6190 5200
rect 6270 5190 6360 5200
rect 6400 5190 7220 5200
rect 8030 5190 8100 5200
rect 8130 5190 8180 5200
rect 8230 5190 8260 5200
rect 8750 5190 8780 5200
rect 8850 5190 8870 5200
rect 8940 5190 9010 5200
rect 9070 5190 9090 5200
rect 9130 5190 9190 5200
rect 9710 5190 9740 5200
rect 9800 5190 9830 5200
rect 9880 5190 9890 5200
rect 9940 5190 9990 5200
rect 0 5180 60 5190
rect 2510 5180 2520 5190
rect 2560 5180 2670 5190
rect 3490 5180 5070 5190
rect 5220 5180 6220 5190
rect 6270 5180 7260 5190
rect 8040 5180 8090 5190
rect 8130 5180 8190 5190
rect 8230 5180 8260 5190
rect 8680 5180 8720 5190
rect 8760 5180 8780 5190
rect 8850 5180 8870 5190
rect 8940 5180 8970 5190
rect 8980 5180 9010 5190
rect 9070 5180 9100 5190
rect 9150 5180 9190 5190
rect 9540 5180 9600 5190
rect 9710 5180 9750 5190
rect 9810 5180 9840 5190
rect 9880 5180 9900 5190
rect 9960 5180 9990 5190
rect 0 5170 40 5180
rect 2550 5170 2680 5180
rect 3480 5170 5070 5180
rect 5220 5170 6230 5180
rect 6280 5170 7280 5180
rect 8040 5170 8090 5180
rect 8140 5170 8190 5180
rect 8640 5170 8720 5180
rect 8760 5170 8790 5180
rect 8850 5170 8880 5180
rect 8940 5170 8960 5180
rect 8990 5170 9020 5180
rect 9070 5170 9100 5180
rect 9160 5170 9190 5180
rect 9520 5170 9610 5180
rect 9720 5170 9750 5180
rect 9820 5170 9840 5180
rect 9880 5170 9910 5180
rect 9970 5170 9990 5180
rect 0 5160 30 5170
rect 2550 5160 2670 5170
rect 3480 5160 5080 5170
rect 5220 5160 7290 5170
rect 8040 5160 8090 5170
rect 8140 5160 8180 5170
rect 8620 5160 8700 5170
rect 8760 5160 8790 5170
rect 8820 5160 8880 5170
rect 8940 5160 8960 5170
rect 8990 5160 9030 5170
rect 9070 5160 9100 5170
rect 9510 5160 9560 5170
rect 9580 5160 9620 5170
rect 9720 5160 9750 5170
rect 9820 5160 9840 5170
rect 9890 5160 9910 5170
rect 9980 5160 9990 5170
rect 0 5150 20 5160
rect 2530 5150 2660 5160
rect 2810 5150 2820 5160
rect 3470 5150 5090 5160
rect 5230 5150 7290 5160
rect 8050 5150 8090 5160
rect 8160 5150 8170 5160
rect 8610 5150 8690 5160
rect 8770 5150 8880 5160
rect 8940 5150 9030 5160
rect 9080 5150 9100 5160
rect 9420 5150 9470 5160
rect 9510 5150 9540 5160
rect 9590 5150 9620 5160
rect 9720 5150 9750 5160
rect 9820 5150 9840 5160
rect 9890 5150 9910 5160
rect 9990 5150 9990 5160
rect 2530 5140 2650 5150
rect 2680 5140 2690 5150
rect 3460 5140 3470 5150
rect 3490 5140 5090 5150
rect 5220 5140 7300 5150
rect 8050 5140 8090 5150
rect 8660 5140 8690 5150
rect 8770 5140 8840 5150
rect 8860 5140 8880 5150
rect 8940 5140 9040 5150
rect 9400 5140 9470 5150
rect 9510 5140 9540 5150
rect 9600 5140 9620 5150
rect 9730 5140 9760 5150
rect 9820 5140 9850 5150
rect 9890 5140 9920 5150
rect 2540 5130 2660 5140
rect 3460 5130 3470 5140
rect 3490 5130 5110 5140
rect 5220 5130 7300 5140
rect 8060 5130 8080 5140
rect 8490 5130 8510 5140
rect 8670 5130 8690 5140
rect 8770 5130 8810 5140
rect 8860 5130 8890 5140
rect 8940 5130 8980 5140
rect 9010 5130 9040 5140
rect 9370 5130 9450 5140
rect 9520 5130 9550 5140
rect 9600 5130 9630 5140
rect 9730 5130 9760 5140
rect 9820 5130 9850 5140
rect 9890 5130 9920 5140
rect 2550 5120 2660 5130
rect 3450 5120 3460 5130
rect 3490 5120 5110 5130
rect 5220 5120 7300 5130
rect 8450 5120 8520 5130
rect 8670 5120 8690 5130
rect 8770 5120 8800 5130
rect 8860 5120 8890 5130
rect 8930 5120 8960 5130
rect 9310 5120 9330 5130
rect 9370 5120 9410 5130
rect 9520 5120 9550 5130
rect 9600 5120 9630 5130
rect 9730 5120 9760 5130
rect 9820 5120 9850 5130
rect 9900 5120 9910 5130
rect 2560 5110 2610 5120
rect 3440 5110 3450 5120
rect 3490 5110 5130 5120
rect 5220 5110 7300 5120
rect 8430 5110 8510 5120
rect 8670 5110 8700 5120
rect 8780 5110 8800 5120
rect 8860 5110 8890 5120
rect 8930 5110 8960 5120
rect 9270 5110 9340 5120
rect 9370 5110 9400 5120
rect 9520 5110 9550 5120
rect 9610 5110 9630 5120
rect 9740 5110 9770 5120
rect 9810 5110 9840 5120
rect 2580 5100 2590 5110
rect 2650 5100 2660 5110
rect 3440 5100 3450 5110
rect 3500 5100 5140 5110
rect 5220 5100 7290 5110
rect 8420 5100 8480 5110
rect 8670 5100 8700 5110
rect 8780 5100 8800 5110
rect 8870 5100 8890 5110
rect 8940 5100 8950 5110
rect 9240 5100 9330 5110
rect 9380 5100 9410 5110
rect 9520 5100 9550 5110
rect 9610 5100 9640 5110
rect 9740 5100 9840 5110
rect 3430 5090 3450 5100
rect 3470 5090 5150 5100
rect 5220 5090 7290 5100
rect 8430 5090 8460 5100
rect 8680 5090 8700 5100
rect 8780 5090 8810 5100
rect 8870 5090 8890 5100
rect 9230 5090 9310 5100
rect 9380 5090 9410 5100
rect 9440 5090 9470 5100
rect 9530 5090 9550 5100
rect 9610 5090 9640 5100
rect 9750 5090 9820 5100
rect 3420 5080 3450 5090
rect 3460 5080 3500 5090
rect 3510 5080 5150 5090
rect 5220 5080 7290 5090
rect 8300 5080 8380 5090
rect 8430 5080 8460 5090
rect 8680 5080 8700 5090
rect 8780 5080 8810 5090
rect 9160 5080 9200 5090
rect 9240 5080 9260 5090
rect 9270 5080 9310 5090
rect 9380 5080 9480 5090
rect 9530 5080 9550 5090
rect 9610 5080 9640 5090
rect 3420 5070 3510 5080
rect 3520 5070 5150 5080
rect 5230 5070 7240 5080
rect 7250 5070 7290 5080
rect 8290 5070 8400 5080
rect 8430 5070 8460 5080
rect 8500 5070 8510 5080
rect 8680 5070 8710 5080
rect 8780 5070 8810 5080
rect 9120 5070 9200 5080
rect 9280 5070 9310 5080
rect 9390 5070 9460 5080
rect 9530 5070 9560 5080
rect 9610 5070 9640 5080
rect 3420 5060 3520 5070
rect 3530 5060 5150 5070
rect 5230 5060 6300 5070
rect 6320 5060 7290 5070
rect 8290 5060 8350 5070
rect 8360 5060 8400 5070
rect 8440 5060 8520 5070
rect 8680 5060 8710 5070
rect 9100 5060 9190 5070
rect 9280 5060 9310 5070
rect 9390 5060 9430 5070
rect 9540 5060 9560 5070
rect 9600 5060 9630 5070
rect 3410 5050 5150 5060
rect 5230 5050 6300 5060
rect 6320 5050 7300 5060
rect 8190 5050 8240 5060
rect 8290 5050 8320 5060
rect 8370 5050 8400 5060
rect 8440 5050 8510 5060
rect 8680 5050 8710 5060
rect 9100 5050 9170 5060
rect 9280 5050 9310 5060
rect 9390 5050 9420 5060
rect 9540 5050 9570 5060
rect 9580 5050 9630 5060
rect 3410 5040 5150 5050
rect 5230 5040 5710 5050
rect 5800 5040 6310 5050
rect 6330 5040 7210 5050
rect 7230 5040 7290 5050
rect 8170 5040 8250 5050
rect 8290 5040 8320 5050
rect 8370 5040 8400 5050
rect 8440 5040 8490 5050
rect 8690 5040 8710 5050
rect 9040 5040 9060 5050
rect 9140 5040 9170 5050
rect 9290 5040 9320 5050
rect 9400 5040 9420 5050
rect 9540 5040 9620 5050
rect 3420 5030 5150 5040
rect 5230 5030 5680 5040
rect 5800 5030 6300 5040
rect 6350 5030 7210 5040
rect 7230 5030 7300 5040
rect 8160 5030 8260 5040
rect 8290 5030 8320 5040
rect 8370 5030 8400 5040
rect 8440 5030 8470 5040
rect 8980 5030 8990 5040
rect 9040 5030 9070 5040
rect 9140 5030 9180 5040
rect 9290 5030 9320 5040
rect 9400 5030 9420 5040
rect 9550 5030 9580 5040
rect 3420 5020 3510 5030
rect 3520 5020 5160 5030
rect 5230 5020 5660 5030
rect 5800 5020 6310 5030
rect 6370 5020 7300 5030
rect 8150 5020 8200 5030
rect 8230 5020 8260 5030
rect 8290 5020 8320 5030
rect 8350 5020 8390 5030
rect 8450 5020 8470 5030
rect 8970 5020 9000 5030
rect 9040 5020 9070 5030
rect 9150 5020 9180 5030
rect 9290 5020 9320 5030
rect 9400 5020 9430 5030
rect 9460 5020 9500 5030
rect 3410 5010 3510 5020
rect 3520 5010 4160 5020
rect 4170 5010 5160 5020
rect 5230 5010 5630 5020
rect 5800 5010 6310 5020
rect 6390 5010 6400 5020
rect 6410 5010 7210 5020
rect 7230 5010 7300 5020
rect 8090 5010 8110 5020
rect 8150 5010 8190 5020
rect 8230 5010 8260 5020
rect 8300 5010 8380 5020
rect 8450 5010 8480 5020
rect 8510 5010 8540 5020
rect 8970 5010 9000 5020
rect 9040 5010 9070 5020
rect 9150 5010 9180 5020
rect 9290 5010 9320 5020
rect 9400 5010 9500 5020
rect 3410 5000 3510 5010
rect 3520 5000 4120 5010
rect 4130 5000 4160 5010
rect 4190 5000 5160 5010
rect 5230 5000 5620 5010
rect 5790 5000 6320 5010
rect 6420 5000 7210 5010
rect 7230 5000 7300 5010
rect 8010 5000 8030 5010
rect 8080 5000 8120 5010
rect 8150 5000 8180 5010
rect 8230 5000 8270 5010
rect 8300 5000 8370 5010
rect 8450 5000 8550 5010
rect 8890 5000 8920 5010
rect 8970 5000 9010 5010
rect 9040 5000 9080 5010
rect 9150 5000 9180 5010
rect 9300 5000 9330 5010
rect 9400 5000 9480 5010
rect 3410 4990 3510 5000
rect 3530 4990 4020 5000
rect 4030 4990 4200 5000
rect 4220 4990 4270 5000
rect 4300 4990 5170 5000
rect 5230 4990 5600 5000
rect 5790 4990 6330 5000
rect 6470 4990 7300 5000
rect 8000 4990 8040 5000
rect 8080 4990 8120 5000
rect 8150 4990 8190 5000
rect 8240 4990 8270 5000
rect 8300 4990 8380 5000
rect 8450 4990 8540 5000
rect 8890 4990 8930 5000
rect 8960 4990 9010 5000
rect 9050 4990 9080 5000
rect 9160 4990 9190 5000
rect 9310 4990 9330 5000
rect 3400 4980 3510 4990
rect 3520 4980 4010 4990
rect 4030 4980 4210 4990
rect 4230 4980 4280 4990
rect 4340 4980 4510 4990
rect 4570 4980 5200 4990
rect 5230 4980 5570 4990
rect 5780 4980 6330 4990
rect 6480 4980 7310 4990
rect 8000 4980 8050 4990
rect 8080 4980 8120 4990
rect 8150 4980 8190 4990
rect 8240 4980 8270 4990
rect 8300 4980 8330 4990
rect 8350 4980 8400 4990
rect 8450 4980 8510 4990
rect 8770 4980 8820 4990
rect 8890 4980 8940 4990
rect 8960 4980 9010 4990
rect 9050 4980 9080 4990
rect 9160 4980 9190 4990
rect 9310 4980 9330 4990
rect 3400 4970 3510 4980
rect 3520 4970 4000 4980
rect 4070 4970 4080 4980
rect 4090 4970 4200 4980
rect 4290 4970 4310 4980
rect 4370 4970 4390 4980
rect 4410 4970 4510 4980
rect 4590 4970 5200 4980
rect 5230 4970 5510 4980
rect 5780 4970 6120 4980
rect 6150 4970 6330 4980
rect 6500 4970 7310 4980
rect 8010 4970 8050 4980
rect 8080 4970 8120 4980
rect 8160 4970 8190 4980
rect 8240 4970 8270 4980
rect 8310 4970 8340 4980
rect 8360 4970 8410 4980
rect 8750 4970 8840 4980
rect 8890 4970 8940 4980
rect 8960 4970 9010 4980
rect 9050 4970 9080 4980
rect 9160 4970 9190 4980
rect 9310 4970 9330 4980
rect 9680 4970 9710 4980
rect 3390 4960 3500 4970
rect 3520 4960 4000 4970
rect 4070 4960 4080 4970
rect 4100 4960 4190 4970
rect 4390 4960 4400 4970
rect 4420 4960 4620 4970
rect 4690 4960 5200 4970
rect 5240 4960 5510 4970
rect 5790 4960 5810 4970
rect 5820 4960 5830 4970
rect 5880 4960 5920 4970
rect 5980 4960 6040 4970
rect 6200 4960 6320 4970
rect 6540 4960 7310 4970
rect 7870 4960 7910 4970
rect 8010 4960 8060 4970
rect 8070 4960 8130 4970
rect 8160 4960 8190 4970
rect 8240 4960 8270 4970
rect 8310 4960 8340 4970
rect 8380 4960 8410 4970
rect 8750 4960 8850 4970
rect 8890 4960 8950 4970
rect 8960 4960 9020 4970
rect 9060 4960 9080 4970
rect 9170 4960 9190 4970
rect 9640 4960 9710 4970
rect 3390 4950 3500 4960
rect 3520 4950 4000 4960
rect 4080 4950 4190 4960
rect 4420 4950 4450 4960
rect 4490 4950 4590 4960
rect 4710 4950 5190 4960
rect 5240 4950 5500 4960
rect 5980 4950 6010 4960
rect 6230 4950 6240 4960
rect 6610 4950 7320 4960
rect 7850 4950 7930 4960
rect 8010 4950 8130 4960
rect 8160 4950 8190 4960
rect 8240 4950 8270 4960
rect 8310 4950 8340 4960
rect 8670 4950 8710 4960
rect 8740 4950 8770 4960
rect 8820 4950 8850 4960
rect 8900 4950 9020 4960
rect 9060 4950 9090 4960
rect 9170 4950 9200 4960
rect 9620 4950 9690 4960
rect 3380 4940 3510 4950
rect 3520 4940 4000 4950
rect 4100 4940 4180 4950
rect 4440 4940 4480 4950
rect 4530 4940 4640 4950
rect 4720 4940 4740 4950
rect 4750 4940 4760 4950
rect 4780 4940 5190 4950
rect 5240 4940 5490 4950
rect 6580 4940 6590 4950
rect 6640 4940 6670 4950
rect 6680 4940 7320 4950
rect 7840 4940 7930 4950
rect 8010 4940 8130 4950
rect 8160 4940 8200 4950
rect 8240 4940 8270 4950
rect 8320 4940 8340 4950
rect 8640 4940 8710 4950
rect 8750 4940 8770 4950
rect 8830 4940 8860 4950
rect 8900 4940 8980 4950
rect 8990 4940 9020 4950
rect 9060 4940 9090 4950
rect 9170 4940 9240 4950
rect 9560 4940 9570 4950
rect 9610 4940 9660 4950
rect 3380 4930 3510 4940
rect 3520 4930 3990 4940
rect 4070 4930 4180 4940
rect 4450 4930 4510 4940
rect 4560 4930 4710 4940
rect 4790 4930 5060 4940
rect 5070 4930 5190 4940
rect 5240 4930 5470 4940
rect 6680 4930 7230 4940
rect 7240 4930 7320 4940
rect 7770 4930 7790 4940
rect 7830 4930 7870 4940
rect 7900 4930 7940 4940
rect 8010 4930 8130 4940
rect 8170 4930 8210 4940
rect 8220 4930 8270 4940
rect 8610 4930 8700 4940
rect 8750 4930 8780 4940
rect 8830 4930 8860 4940
rect 8900 4930 8930 4940
rect 8940 4930 8980 4940
rect 9000 4930 9020 4940
rect 9060 4930 9090 4940
rect 9150 4930 9260 4940
rect 9550 4930 9580 4940
rect 9620 4930 9650 4940
rect 3380 4920 3480 4930
rect 3500 4920 3510 4930
rect 3520 4920 3990 4930
rect 4070 4920 4120 4930
rect 4150 4920 4170 4930
rect 4380 4920 4390 4930
rect 4490 4920 4540 4930
rect 4610 4920 4740 4930
rect 4770 4920 4790 4930
rect 4820 4920 5040 4930
rect 5090 4920 5190 4930
rect 5240 4920 5450 4930
rect 6690 4920 7320 4930
rect 7770 4920 7790 4930
rect 7830 4920 7860 4930
rect 7910 4920 7940 4930
rect 8010 4920 8130 4930
rect 8170 4920 8260 4930
rect 8610 4920 8660 4930
rect 8750 4920 8780 4930
rect 8820 4920 8850 4930
rect 8910 4920 8930 4930
rect 8950 4920 8980 4930
rect 9000 4920 9020 4930
rect 9070 4920 9090 4930
rect 9140 4920 9280 4930
rect 9540 4920 9580 4930
rect 9620 4920 9650 4930
rect 3380 4910 3480 4920
rect 3500 4910 3910 4920
rect 3930 4910 3970 4920
rect 4050 4910 4110 4920
rect 4160 4910 4170 4920
rect 4530 4910 4570 4920
rect 4680 4910 4790 4920
rect 4830 4910 5030 4920
rect 5080 4910 5190 4920
rect 5250 4910 5420 4920
rect 6690 4910 7320 4920
rect 7700 4910 7710 4920
rect 7770 4910 7800 4920
rect 7830 4910 7860 4920
rect 7910 4910 7940 4920
rect 8020 4910 8140 4920
rect 8180 4910 8250 4920
rect 8530 4910 8540 4920
rect 8610 4910 8640 4920
rect 8750 4910 8780 4920
rect 8800 4910 8850 4920
rect 8910 4910 8940 4920
rect 8950 4910 8980 4920
rect 9000 4910 9030 4920
rect 9070 4910 9090 4920
rect 9130 4910 9290 4920
rect 9460 4910 9480 4920
rect 9540 4910 9580 4920
rect 9620 4910 9660 4920
rect 3330 4900 3340 4910
rect 3410 4900 3470 4910
rect 3490 4900 3900 4910
rect 3940 4900 3950 4910
rect 4030 4900 4070 4910
rect 4580 4900 4600 4910
rect 4730 4900 4830 4910
rect 4840 4900 4850 4910
rect 4870 4900 5020 4910
rect 5070 4900 5180 4910
rect 5250 4900 5380 4910
rect 6700 4900 7230 4910
rect 7240 4900 7320 4910
rect 7690 4900 7720 4910
rect 7770 4900 7800 4910
rect 7830 4900 7860 4910
rect 7910 4900 7940 4910
rect 8020 4900 8060 4910
rect 8070 4900 8090 4910
rect 8110 4900 8140 4910
rect 8490 4900 8560 4910
rect 8610 4900 8640 4910
rect 8750 4900 8840 4910
rect 8910 4900 8940 4910
rect 9000 4900 9030 4910
rect 9120 4900 9300 4910
rect 9460 4900 9490 4910
rect 9540 4900 9580 4910
rect 9630 4900 9720 4910
rect 3410 4890 3460 4900
rect 3480 4890 3750 4900
rect 3760 4890 3860 4900
rect 3870 4890 3890 4900
rect 3920 4890 3930 4900
rect 4020 4890 4050 4900
rect 4790 4890 4820 4900
rect 4880 4890 5030 4900
rect 5060 4890 5100 4900
rect 5110 4890 5180 4900
rect 5250 4890 5380 4900
rect 6700 4890 7230 4900
rect 7240 4890 7320 4900
rect 7690 4890 7730 4900
rect 7770 4890 7800 4900
rect 7830 4890 7870 4900
rect 7910 4890 7950 4900
rect 8020 4890 8060 4900
rect 8110 4890 8140 4900
rect 8480 4890 8570 4900
rect 8610 4890 8640 4900
rect 8680 4890 8700 4900
rect 8760 4890 8830 4900
rect 8910 4890 8940 4900
rect 9010 4890 9030 4900
rect 9110 4890 9300 4900
rect 9390 4890 9410 4900
rect 9460 4890 9500 4900
rect 9540 4890 9590 4900
rect 9630 4890 9710 4900
rect 3340 4880 3360 4890
rect 3430 4880 3470 4890
rect 3480 4880 3710 4890
rect 3760 4880 3840 4890
rect 3850 4880 3870 4890
rect 3920 4880 3930 4890
rect 4010 4880 4030 4890
rect 4910 4880 5180 4890
rect 5250 4880 5380 4890
rect 6710 4880 7190 4890
rect 7210 4880 7230 4890
rect 7240 4880 7320 4890
rect 7690 4880 7740 4890
rect 7780 4880 7800 4890
rect 7830 4880 7870 4890
rect 7910 4880 7950 4890
rect 8020 4880 8060 4890
rect 8120 4880 8130 4890
rect 8470 4880 8510 4890
rect 8550 4880 8580 4890
rect 8620 4880 8700 4890
rect 8760 4880 8790 4890
rect 8810 4880 8840 4890
rect 8920 4880 8940 4890
rect 9100 4880 9310 4890
rect 9340 4880 9350 4890
rect 9390 4880 9420 4890
rect 9460 4880 9510 4890
rect 9540 4880 9590 4890
rect 9630 4880 9680 4890
rect 3330 4870 3350 4880
rect 3430 4870 3700 4880
rect 3750 4870 3790 4880
rect 3800 4870 3870 4880
rect 4000 4870 4020 4880
rect 4850 4870 4880 4880
rect 4930 4870 5180 4880
rect 5250 4870 5380 4880
rect 6710 4870 7210 4880
rect 7250 4870 7330 4880
rect 7690 4870 7750 4880
rect 7780 4870 7810 4880
rect 7840 4870 7870 4880
rect 7920 4870 7950 4880
rect 8030 4870 8060 4880
rect 8470 4870 8500 4880
rect 8550 4870 8580 4880
rect 8620 4870 8700 4880
rect 8760 4870 8790 4880
rect 8820 4870 8850 4880
rect 8920 4870 8940 4880
rect 9100 4870 9360 4880
rect 9390 4870 9420 4880
rect 9470 4870 9520 4880
rect 9540 4870 9560 4880
rect 9570 4870 9590 4880
rect 9630 4870 9670 4880
rect 3330 4860 3340 4870
rect 3420 4860 3690 4870
rect 3790 4860 3830 4870
rect 3850 4860 3860 4870
rect 3990 4860 4000 4870
rect 4880 4860 4920 4870
rect 4950 4860 5180 4870
rect 5240 4860 5370 4870
rect 6700 4860 7330 4870
rect 7700 4860 7760 4870
rect 7780 4860 7810 4870
rect 7840 4860 7870 4870
rect 7920 4860 7950 4870
rect 8030 4860 8060 4870
rect 8480 4860 8510 4870
rect 8550 4860 8580 4870
rect 8620 4860 8670 4870
rect 8770 4860 8790 4870
rect 8830 4860 8870 4870
rect 9090 4860 9350 4870
rect 9400 4860 9420 4870
rect 9470 4860 9560 4870
rect 9570 4860 9590 4870
rect 9640 4860 9670 4870
rect 3410 4850 3670 4860
rect 3970 4850 3980 4860
rect 4910 4850 4930 4860
rect 4960 4850 5190 4860
rect 5240 4850 5370 4860
rect 6710 4850 7330 4860
rect 7700 4850 7810 4860
rect 7840 4850 7870 4860
rect 7910 4850 7950 4860
rect 8310 4850 8370 4860
rect 8480 4850 8510 4860
rect 8550 4850 8580 4860
rect 8630 4850 8650 4860
rect 8770 4850 8800 4860
rect 8840 4850 8870 4860
rect 9080 4850 9330 4860
rect 9400 4850 9420 4860
rect 9470 4850 9490 4860
rect 9510 4850 9550 4860
rect 9570 4850 9600 4860
rect 9640 4850 9670 4860
rect 3410 4840 3670 4850
rect 4970 4840 5180 4850
rect 5240 4840 5370 4850
rect 6710 4840 7330 4850
rect 7710 4840 7730 4850
rect 7750 4840 7810 4850
rect 7840 4840 7940 4850
rect 8290 4840 8370 4850
rect 8480 4840 8510 4850
rect 8530 4840 8570 4850
rect 8630 4840 8650 4850
rect 8770 4840 8800 4850
rect 9080 4840 9320 4850
rect 9400 4840 9430 4850
rect 9470 4840 9500 4850
rect 9510 4840 9550 4850
rect 9570 4840 9600 4850
rect 9640 4840 9670 4850
rect 9710 4840 9750 4850
rect 3400 4830 3570 4840
rect 3590 4830 3660 4840
rect 3950 4830 3960 4840
rect 4990 4830 5180 4840
rect 5240 4830 5370 4840
rect 6720 4830 7270 4840
rect 7290 4830 7340 4840
rect 7710 4830 7740 4840
rect 7760 4830 7820 4840
rect 7850 4830 7940 4840
rect 8280 4830 8370 4840
rect 8480 4830 8570 4840
rect 8630 4830 8650 4840
rect 8710 4830 8730 4840
rect 8780 4830 8790 4840
rect 9070 4830 9330 4840
rect 9400 4830 9430 4840
rect 9480 4830 9500 4840
rect 9520 4830 9550 4840
rect 9570 4830 9600 4840
rect 9640 4830 9750 4840
rect 3390 4820 3560 4830
rect 3590 4820 3640 4830
rect 5000 4820 5170 4830
rect 5240 4820 5370 4830
rect 6720 4820 7240 4830
rect 7250 4820 7340 4830
rect 7710 4820 7740 4830
rect 7770 4820 7820 4830
rect 7850 4820 7920 4830
rect 8200 4820 8230 4830
rect 8270 4820 8310 4830
rect 8490 4820 8550 4830
rect 8630 4820 8660 4830
rect 8670 4820 8740 4830
rect 9070 4820 9330 4830
rect 9410 4820 9430 4830
rect 9480 4820 9510 4830
rect 9530 4820 9550 4830
rect 9580 4820 9600 4830
rect 9650 4820 9730 4830
rect 2420 4810 2430 4820
rect 3390 4810 3550 4820
rect 3580 4810 3630 4820
rect 5030 4810 5170 4820
rect 5240 4810 5360 4820
rect 6720 4810 7340 4820
rect 7710 4810 7740 4820
rect 7780 4810 7820 4820
rect 8200 4810 8230 4820
rect 8270 4810 8300 4820
rect 8490 4810 8520 4820
rect 8630 4810 8730 4820
rect 9060 4810 9330 4820
rect 9410 4810 9440 4820
rect 9480 4810 9510 4820
rect 9580 4810 9610 4820
rect 9650 4810 9690 4820
rect 3260 4800 3270 4810
rect 3380 4800 3550 4810
rect 3570 4800 3620 4810
rect 5040 4800 5170 4810
rect 5240 4800 5360 4810
rect 6730 4800 7350 4810
rect 7720 4800 7740 4810
rect 7790 4800 7820 4810
rect 8120 4800 8150 4810
rect 8200 4800 8240 4810
rect 8270 4800 8310 4810
rect 8490 4800 8520 4810
rect 8630 4800 8700 4810
rect 9060 4800 9330 4810
rect 9410 4800 9440 4810
rect 9480 4800 9510 4810
rect 9580 4800 9610 4810
rect 3380 4790 3540 4800
rect 3560 4790 3610 4800
rect 5050 4790 5180 4800
rect 5240 4790 5350 4800
rect 6720 4790 7350 4800
rect 7720 4790 7750 4800
rect 8120 4790 8160 4800
rect 8210 4790 8240 4800
rect 8280 4790 8370 4800
rect 8500 4790 8520 4800
rect 9000 4790 9030 4800
rect 9050 4790 9340 4800
rect 9410 4790 9440 4800
rect 9490 4790 9520 4800
rect 9590 4790 9600 4800
rect 3370 4780 3540 4790
rect 3560 4780 3600 4790
rect 5040 4780 5200 4790
rect 5240 4780 5340 4790
rect 5780 4780 5840 4790
rect 6720 4780 7340 4790
rect 7720 4780 7740 4790
rect 8030 4780 8080 4790
rect 8120 4780 8170 4790
rect 8210 4780 8240 4790
rect 8280 4780 8390 4790
rect 8500 4780 8530 4790
rect 9000 4780 9030 4790
rect 9050 4780 9340 4790
rect 9420 4780 9450 4790
rect 9490 4780 9520 4790
rect 3360 4770 3530 4780
rect 3550 4770 3590 4780
rect 5060 4770 5230 4780
rect 5240 4770 5340 4780
rect 5780 4770 5880 4780
rect 6720 4770 7340 4780
rect 8010 4770 8090 4780
rect 8130 4770 8180 4780
rect 8210 4770 8240 4780
rect 8300 4770 8390 4780
rect 8500 4770 8530 4780
rect 8920 4770 8940 4780
rect 9010 4770 9300 4780
rect 9310 4770 9340 4780
rect 9420 4770 9450 4780
rect 9490 4770 9520 4780
rect 3260 4760 3280 4770
rect 3360 4760 3520 4770
rect 3560 4760 3580 4770
rect 5090 4760 5340 4770
rect 5760 4760 5900 4770
rect 6720 4760 7350 4770
rect 8000 4760 8100 4770
rect 8130 4760 8200 4770
rect 8210 4760 8250 4770
rect 8360 4760 8390 4770
rect 8500 4760 8530 4770
rect 8920 4760 8950 4770
rect 9010 4760 9300 4770
rect 9320 4760 9340 4770
rect 9420 4760 9450 4770
rect 3260 4750 3280 4760
rect 3370 4750 3520 4760
rect 3560 4750 3570 4760
rect 3840 4750 3850 4760
rect 5100 4750 5340 4760
rect 5760 4750 5910 4760
rect 6730 4750 7310 4760
rect 7320 4750 7360 4760
rect 7990 4750 8040 4760
rect 8070 4750 8100 4760
rect 8130 4750 8200 4760
rect 8220 4750 8250 4760
rect 8370 4750 8390 4760
rect 8810 4750 8870 4760
rect 8920 4750 8960 4760
rect 9010 4750 9300 4760
rect 9320 4750 9350 4760
rect 9430 4750 9440 4760
rect 3260 4740 3280 4750
rect 3370 4740 3510 4750
rect 5110 4740 5340 4750
rect 5750 4740 5920 4750
rect 6720 4740 6730 4750
rect 6740 4740 7300 4750
rect 7310 4740 7360 4750
rect 7880 4740 7950 4750
rect 7990 4740 8030 4750
rect 8070 4740 8100 4750
rect 8130 4740 8250 4750
rect 8300 4740 8310 4750
rect 8360 4740 8390 4750
rect 8800 4740 8880 4750
rect 8930 4740 8980 4750
rect 9010 4740 9300 4750
rect 9320 4740 9350 4750
rect 9890 4740 9990 4750
rect 3270 4730 3290 4740
rect 3360 4730 3510 4740
rect 5120 4730 5330 4740
rect 5740 4730 5920 4740
rect 6750 4730 7360 4740
rect 7870 4730 7950 4740
rect 7990 4730 8020 4740
rect 8070 4730 8110 4740
rect 8140 4730 8170 4740
rect 8190 4730 8250 4740
rect 8290 4730 8380 4740
rect 8790 4730 8830 4740
rect 8850 4730 8890 4740
rect 8930 4730 8990 4740
rect 9020 4730 9290 4740
rect 9320 4730 9350 4740
rect 9870 4730 9990 4740
rect 3270 4720 3290 4730
rect 3360 4720 3500 4730
rect 5140 4720 5330 4730
rect 5740 4720 5940 4730
rect 6760 4720 7290 4730
rect 7310 4720 7360 4730
rect 7860 4720 7950 4730
rect 7990 4720 8030 4730
rect 8070 4720 8110 4730
rect 8140 4720 8170 4730
rect 8200 4720 8260 4730
rect 8290 4720 8380 4730
rect 8790 4720 8820 4730
rect 8860 4720 8890 4730
rect 8930 4720 9000 4730
rect 9020 4720 9290 4730
rect 9850 4720 9990 4730
rect 3070 4710 3080 4720
rect 3270 4710 3290 4720
rect 3370 4710 3500 4720
rect 5150 4710 5200 4720
rect 5220 4710 5330 4720
rect 5770 4710 5930 4720
rect 6760 4710 7360 4720
rect 7760 4710 7800 4720
rect 7860 4710 7890 4720
rect 7990 4710 8030 4720
rect 8080 4710 8110 4720
rect 8140 4710 8170 4720
rect 8210 4710 8260 4720
rect 8300 4710 8360 4720
rect 8790 4710 8820 4720
rect 8860 4710 8890 4720
rect 8930 4710 8960 4720
rect 8970 4710 9280 4720
rect 9840 4710 9990 4720
rect 3270 4700 3290 4710
rect 3370 4700 3500 4710
rect 5110 4700 5120 4710
rect 5160 4700 5190 4710
rect 5230 4700 5320 4710
rect 5780 4700 5930 4710
rect 6750 4700 7360 4710
rect 7740 4700 7820 4710
rect 7860 4700 7890 4710
rect 8000 4700 8030 4710
rect 8080 4700 8110 4710
rect 8150 4700 8180 4710
rect 8220 4700 8260 4710
rect 8630 4700 8670 4710
rect 8790 4700 8810 4710
rect 8870 4700 8900 4710
rect 8930 4700 8960 4710
rect 8980 4700 9280 4710
rect 9840 4700 9990 4710
rect 3270 4690 3290 4700
rect 3370 4690 3490 4700
rect 5120 4690 5130 4700
rect 5170 4690 5310 4700
rect 5800 4690 5820 4700
rect 5830 4690 5920 4700
rect 6700 4690 6710 4700
rect 6760 4690 7370 4700
rect 7730 4690 7830 4700
rect 7860 4690 7890 4700
rect 8000 4690 8030 4700
rect 8080 4690 8110 4700
rect 8150 4690 8180 4700
rect 8230 4690 8260 4700
rect 8580 4690 8670 4700
rect 8790 4690 8820 4700
rect 8870 4690 8900 4700
rect 8940 4690 8960 4700
rect 8990 4690 9280 4700
rect 9830 4690 9990 4700
rect 3270 4680 3290 4690
rect 3390 4680 3480 4690
rect 5120 4680 5140 4690
rect 5180 4680 5240 4690
rect 5250 4680 5310 4690
rect 6700 4680 6710 4690
rect 6750 4680 7370 4690
rect 7660 4680 7690 4690
rect 7730 4680 7760 4690
rect 7790 4680 7830 4690
rect 7860 4680 7960 4690
rect 8000 4680 8030 4690
rect 8080 4680 8110 4690
rect 8150 4680 8180 4690
rect 8570 4680 8640 4690
rect 8790 4680 8820 4690
rect 8870 4680 8900 4690
rect 8940 4680 8970 4690
rect 9000 4680 9270 4690
rect 9820 4680 9990 4690
rect 3150 4670 3170 4680
rect 3270 4670 3280 4680
rect 3390 4670 3480 4680
rect 5130 4670 5140 4680
rect 5180 4670 5240 4680
rect 5250 4670 5300 4680
rect 6750 4670 7300 4680
rect 7330 4670 7380 4680
rect 7620 4670 7690 4680
rect 7730 4670 7760 4680
rect 7800 4670 7830 4680
rect 7870 4670 7970 4680
rect 8000 4670 8030 4680
rect 8080 4670 8110 4680
rect 8150 4670 8180 4680
rect 8510 4670 8520 4680
rect 8570 4670 8640 4680
rect 8790 4670 8820 4680
rect 8880 4670 8900 4680
rect 8940 4670 8970 4680
rect 9000 4670 9270 4680
rect 9810 4670 9990 4680
rect 3150 4660 3160 4670
rect 3380 4660 3400 4670
rect 3420 4660 3480 4670
rect 5140 4660 5150 4670
rect 5190 4660 5220 4670
rect 5250 4660 5300 4670
rect 6690 4660 6700 4670
rect 6750 4660 7310 4670
rect 7320 4660 7380 4670
rect 7610 4660 7680 4670
rect 7730 4660 7760 4670
rect 7800 4660 7830 4670
rect 7890 4660 7970 4670
rect 8010 4660 8040 4670
rect 8060 4660 8110 4670
rect 8510 4660 8540 4670
rect 8610 4660 8640 4670
rect 8800 4660 8830 4670
rect 8880 4660 8900 4670
rect 8940 4660 8970 4670
rect 9000 4660 9260 4670
rect 9800 4660 9990 4670
rect 3370 4650 3400 4660
rect 3420 4650 3470 4660
rect 5200 4650 5240 4660
rect 5250 4650 5300 4660
rect 6690 4650 6700 4660
rect 6750 4650 7240 4660
rect 7260 4650 7380 4660
rect 7600 4650 7650 4660
rect 7730 4650 7770 4660
rect 7790 4650 7830 4660
rect 7940 4650 7980 4660
rect 8010 4650 8110 4660
rect 8500 4650 8540 4660
rect 8610 4650 8640 4660
rect 8800 4650 8830 4660
rect 8880 4650 8910 4660
rect 8940 4650 8970 4660
rect 8990 4650 9260 4660
rect 9790 4650 9990 4660
rect 3330 4640 3340 4650
rect 3370 4640 3390 4650
rect 3410 4640 3460 4650
rect 5210 4640 5300 4650
rect 6750 4640 7380 4650
rect 7500 4640 7570 4650
rect 7610 4640 7640 4650
rect 7740 4640 7820 4650
rect 7950 4640 7980 4650
rect 8020 4640 8090 4650
rect 8500 4640 8550 4650
rect 8620 4640 8650 4650
rect 8800 4640 8830 4650
rect 8880 4640 8910 4650
rect 8950 4640 8980 4650
rect 8990 4640 9250 4650
rect 9780 4640 9990 4650
rect 3320 4630 3340 4640
rect 3410 4630 3460 4640
rect 5210 4630 5290 4640
rect 6750 4630 7380 4640
rect 7480 4630 7580 4640
rect 7610 4630 7640 4640
rect 7740 4630 7810 4640
rect 7940 4630 7970 4640
rect 8330 4630 8340 4640
rect 8500 4630 8550 4640
rect 8620 4630 8650 4640
rect 8800 4630 8840 4640
rect 8870 4630 8910 4640
rect 8960 4630 8970 4640
rect 8990 4630 9250 4640
rect 9770 4630 9990 4640
rect 3310 4620 3340 4630
rect 3410 4620 3420 4630
rect 5220 4620 5280 4630
rect 6750 4620 7380 4630
rect 7480 4620 7530 4630
rect 7540 4620 7580 4630
rect 7610 4620 7640 4630
rect 7650 4620 7690 4630
rect 7740 4620 7810 4630
rect 7880 4620 7970 4630
rect 8290 4620 8370 4630
rect 8500 4620 8560 4630
rect 8620 4620 8650 4630
rect 8810 4620 8900 4630
rect 8980 4620 9250 4630
rect 9760 4620 9990 4630
rect 3310 4610 3340 4620
rect 3430 4610 3450 4620
rect 5220 4610 5280 4620
rect 6740 4610 7380 4620
rect 7480 4610 7510 4620
rect 7550 4610 7580 4620
rect 7610 4610 7690 4620
rect 7740 4610 7770 4620
rect 7780 4610 7820 4620
rect 7880 4610 7960 4620
rect 8280 4610 8380 4620
rect 8500 4610 8560 4620
rect 8620 4610 8650 4620
rect 8820 4610 8890 4620
rect 8980 4610 9240 4620
rect 9750 4610 9990 4620
rect 3300 4600 3350 4610
rect 3420 4600 3450 4610
rect 5230 4600 5280 4610
rect 6740 4600 7310 4610
rect 7330 4600 7390 4610
rect 7480 4600 7520 4610
rect 7550 4600 7580 4610
rect 7610 4600 7680 4610
rect 7750 4600 7770 4610
rect 7790 4600 7830 4610
rect 7890 4600 7940 4610
rect 8220 4600 8250 4610
rect 8280 4600 8320 4610
rect 8350 4600 8380 4610
rect 8500 4600 8530 4610
rect 8540 4600 8570 4610
rect 8630 4600 8650 4610
rect 8980 4600 9240 4610
rect 9740 4600 9990 4610
rect 3300 4590 3340 4600
rect 3380 4590 3440 4600
rect 5240 4590 5280 4600
rect 6740 4590 7320 4600
rect 7340 4590 7380 4600
rect 7490 4590 7520 4600
rect 7550 4590 7580 4600
rect 7620 4590 7650 4600
rect 7750 4590 7780 4600
rect 7800 4590 7840 4600
rect 8180 4590 8250 4600
rect 8280 4590 8310 4600
rect 8360 4590 8390 4600
rect 8500 4590 8530 4600
rect 8540 4590 8580 4600
rect 8630 4590 8660 4600
rect 8970 4590 9240 4600
rect 9730 4590 9990 4600
rect 3270 4580 3330 4590
rect 3380 4580 3440 4590
rect 3460 4580 3470 4590
rect 5240 4580 5280 4590
rect 5810 4580 5820 4590
rect 5960 4580 5980 4590
rect 6740 4580 7320 4590
rect 7350 4580 7380 4590
rect 7490 4580 7520 4590
rect 7530 4580 7580 4590
rect 7620 4580 7650 4590
rect 7750 4580 7780 4590
rect 7810 4580 7840 4590
rect 8160 4580 8240 4590
rect 8280 4580 8320 4590
rect 8360 4580 8390 4590
rect 8500 4580 8520 4590
rect 8550 4580 8580 4590
rect 8630 4580 8660 4590
rect 8970 4580 9240 4590
rect 9720 4580 9990 4590
rect 3270 4570 3330 4580
rect 3360 4570 3440 4580
rect 5240 4570 5280 4580
rect 5800 4570 5810 4580
rect 6740 4570 7320 4580
rect 7330 4570 7380 4580
rect 7490 4570 7570 4580
rect 7620 4570 7650 4580
rect 7750 4570 7780 4580
rect 8110 4570 8120 4580
rect 8160 4570 8210 4580
rect 8290 4570 8320 4580
rect 8350 4570 8390 4580
rect 8500 4570 8520 4580
rect 8550 4570 8590 4580
rect 8630 4570 8660 4580
rect 8970 4570 9240 4580
rect 9710 4570 9980 4580
rect 3270 4560 3330 4570
rect 3360 4560 3380 4570
rect 3390 4560 3440 4570
rect 5250 4560 5290 4570
rect 5800 4560 5830 4570
rect 5870 4560 5900 4570
rect 5950 4560 6000 4570
rect 6730 4560 7320 4570
rect 7360 4560 7370 4570
rect 7490 4560 7560 4570
rect 7620 4560 7650 4570
rect 7680 4560 7720 4570
rect 7760 4560 7770 4570
rect 8100 4560 8130 4570
rect 8160 4560 8190 4570
rect 8290 4560 8320 4570
rect 8340 4560 8390 4570
rect 8490 4560 8600 4570
rect 8640 4560 8660 4570
rect 8960 4560 9230 4570
rect 9700 4560 9980 4570
rect 3260 4550 3270 4560
rect 3280 4550 3320 4560
rect 3340 4550 3440 4560
rect 5250 4550 5290 4560
rect 5810 4550 5830 4560
rect 5870 4550 5910 4560
rect 5930 4550 6010 4560
rect 6090 4550 6110 4560
rect 6730 4550 7320 4560
rect 7360 4550 7370 4560
rect 7500 4550 7530 4560
rect 7620 4550 7720 4560
rect 8100 4550 8130 4560
rect 8160 4550 8190 4560
rect 8290 4550 8380 4560
rect 8490 4550 8600 4560
rect 8960 4550 9230 4560
rect 9700 4550 9980 4560
rect 3280 4540 3320 4550
rect 3340 4540 3420 4550
rect 3430 4540 3440 4550
rect 5260 4540 5290 4550
rect 5810 4540 5840 4550
rect 5870 4540 6020 4550
rect 6060 4540 6120 4550
rect 6720 4540 7330 4550
rect 7360 4540 7370 4550
rect 7500 4540 7530 4550
rect 7630 4540 7700 4550
rect 8010 4540 8040 4550
rect 8070 4540 8090 4550
rect 8100 4540 8130 4550
rect 8160 4540 8200 4550
rect 8230 4540 8240 4550
rect 8300 4540 8370 4550
rect 8490 4540 8530 4550
rect 8580 4540 8600 4550
rect 8950 4540 9230 4550
rect 9690 4540 9960 4550
rect 3270 4530 3310 4540
rect 3320 4530 3340 4540
rect 3350 4530 3420 4540
rect 5260 4530 5290 4540
rect 5820 4530 5840 4540
rect 5870 4530 6020 4540
rect 6040 4530 6130 4540
rect 6160 4530 6170 4540
rect 6720 4530 7330 4540
rect 7360 4530 7380 4540
rect 7500 4530 7530 4540
rect 7630 4530 7670 4540
rect 7930 4530 7960 4540
rect 8010 4530 8040 4540
rect 8060 4530 8090 4540
rect 8100 4530 8130 4540
rect 8170 4530 8250 4540
rect 8300 4530 8370 4540
rect 8490 4530 8520 4540
rect 8950 4530 9230 4540
rect 9680 4530 9950 4540
rect 3270 4520 3300 4530
rect 3330 4520 3420 4530
rect 5270 4520 5290 4530
rect 5830 4520 5850 4530
rect 5870 4520 6130 4530
rect 6150 4520 6180 4530
rect 6720 4520 7330 4530
rect 7360 4520 7390 4530
rect 7500 4520 7530 4530
rect 7910 4520 7980 4530
rect 8020 4520 8050 4530
rect 8060 4520 8130 4530
rect 8170 4520 8250 4530
rect 8300 4520 8330 4530
rect 8340 4520 8390 4530
rect 8490 4520 8520 4530
rect 8950 4520 9230 4530
rect 9670 4520 9940 4530
rect 3010 4510 3020 4520
rect 3260 4510 3300 4520
rect 3330 4510 3410 4520
rect 5280 4510 5300 4520
rect 5830 4510 5840 4520
rect 5870 4510 6190 4520
rect 6710 4510 7330 4520
rect 7360 4510 7400 4520
rect 7500 4510 7540 4520
rect 7900 4510 7990 4520
rect 8020 4510 8050 4520
rect 8060 4510 8140 4520
rect 8170 4510 8230 4520
rect 8300 4510 8330 4520
rect 8350 4510 8400 4520
rect 8940 4510 9220 4520
rect 9660 4510 9940 4520
rect 3010 4500 3030 4510
rect 3260 4500 3300 4510
rect 3310 4500 3410 4510
rect 5280 4500 5300 4510
rect 5870 4500 6170 4510
rect 6710 4500 7330 4510
rect 7380 4500 7400 4510
rect 7510 4500 7530 4510
rect 7820 4500 7850 4510
rect 7890 4500 7940 4510
rect 7950 4500 7990 4510
rect 8020 4500 8140 4510
rect 8170 4500 8200 4510
rect 8300 4500 8330 4510
rect 8360 4500 8400 4510
rect 8940 4500 9220 4510
rect 9650 4500 9930 4510
rect 3010 4490 3030 4500
rect 3270 4490 3400 4500
rect 5280 4490 5310 4500
rect 5880 4490 6170 4500
rect 6710 4490 7330 4500
rect 7370 4490 7410 4500
rect 7780 4490 7860 4500
rect 7890 4490 7920 4500
rect 7960 4490 7990 4500
rect 8030 4490 8140 4500
rect 8180 4490 8210 4500
rect 8300 4490 8340 4500
rect 8370 4490 8400 4500
rect 8930 4490 9220 4500
rect 9640 4490 9930 4500
rect 3280 4480 3400 4490
rect 5290 4480 5310 4490
rect 5900 4480 6160 4490
rect 6710 4480 7340 4490
rect 7370 4480 7420 4490
rect 7760 4480 7850 4490
rect 7890 4480 7920 4490
rect 7960 4480 8000 4490
rect 8030 4480 8140 4490
rect 8180 4480 8210 4490
rect 8310 4480 8340 4490
rect 8930 4480 9220 4490
rect 9630 4480 9910 4490
rect 3000 4470 3030 4480
rect 3090 4470 3110 4480
rect 3280 4470 3400 4480
rect 5300 4470 5310 4480
rect 5920 4470 6140 4480
rect 6710 4470 7340 4480
rect 7370 4470 7420 4480
rect 7760 4470 7830 4480
rect 7890 4470 7920 4480
rect 7960 4470 8000 4480
rect 8030 4470 8080 4480
rect 8090 4470 8140 4480
rect 8180 4470 8280 4480
rect 8310 4470 8330 4480
rect 8920 4470 9210 4480
rect 9620 4470 9890 4480
rect 3010 4460 3030 4470
rect 3090 4460 3110 4470
rect 3290 4460 3390 4470
rect 5310 4460 5320 4470
rect 5930 4460 6130 4470
rect 6710 4460 7340 4470
rect 7360 4460 7410 4470
rect 7800 4460 7830 4470
rect 7890 4460 7920 4470
rect 7970 4460 8000 4470
rect 8040 4460 8080 4470
rect 8090 4460 8140 4470
rect 8180 4460 8280 4470
rect 8920 4460 9210 4470
rect 9610 4460 9880 4470
rect 2850 4450 2860 4460
rect 3000 4450 3020 4460
rect 3090 4450 3110 4460
rect 3300 4450 3390 4460
rect 5310 4450 5320 4460
rect 5960 4450 6120 4460
rect 6710 4450 7340 4460
rect 7350 4450 7410 4460
rect 7800 4450 7830 4460
rect 7890 4450 7920 4460
rect 7970 4450 8000 4460
rect 8040 4450 8080 4460
rect 8100 4450 8140 4460
rect 8190 4450 8260 4460
rect 8910 4450 9210 4460
rect 9600 4450 9870 4460
rect 3030 4440 3040 4450
rect 3300 4440 3390 4450
rect 5320 4440 5330 4450
rect 6070 4440 6100 4450
rect 6700 4440 7410 4450
rect 7800 4440 7840 4450
rect 7890 4440 7920 4450
rect 7970 4440 8010 4450
rect 8040 4440 8080 4450
rect 8110 4440 8140 4450
rect 8190 4440 8210 4450
rect 8910 4440 9210 4450
rect 9590 4440 9870 4450
rect 2830 4430 2840 4440
rect 3020 4430 3040 4440
rect 3260 4430 3270 4440
rect 3310 4430 3380 4440
rect 5320 4430 5340 4440
rect 6690 4430 7340 4440
rect 7370 4430 7410 4440
rect 7810 4430 7840 4440
rect 7900 4430 7930 4440
rect 7970 4430 8010 4440
rect 8050 4430 8080 4440
rect 8110 4430 8140 4440
rect 8870 4430 9210 4440
rect 9580 4430 9840 4440
rect 2980 4420 2990 4430
rect 3020 4420 3050 4430
rect 3260 4420 3270 4430
rect 3310 4420 3370 4430
rect 5330 4420 5340 4430
rect 6680 4420 7240 4430
rect 7250 4420 7270 4430
rect 7280 4420 7340 4430
rect 7380 4420 7410 4430
rect 7810 4420 7840 4430
rect 7900 4420 7930 4430
rect 7970 4420 8010 4430
rect 8050 4420 8080 4430
rect 8120 4420 8130 4430
rect 8850 4420 9200 4430
rect 9570 4420 9830 4430
rect 3000 4410 3010 4420
rect 3020 4410 3050 4420
rect 3270 4410 3290 4420
rect 3320 4410 3370 4420
rect 5330 4410 5350 4420
rect 6680 4410 7240 4420
rect 7250 4410 7260 4420
rect 7300 4410 7340 4420
rect 7370 4410 7420 4420
rect 7810 4410 7840 4420
rect 7900 4410 7940 4420
rect 7970 4410 8000 4420
rect 8060 4410 8080 4420
rect 8850 4410 8880 4420
rect 8900 4410 9200 4420
rect 9560 4410 9840 4420
rect 3000 4400 3010 4410
rect 3020 4400 3050 4410
rect 3240 4400 3260 4410
rect 3320 4400 3360 4410
rect 5330 4400 5360 4410
rect 5810 4400 5820 4410
rect 6680 4400 7240 4410
rect 7250 4400 7290 4410
rect 7300 4400 7340 4410
rect 7370 4400 7420 4410
rect 7810 4400 7850 4410
rect 7910 4400 8000 4410
rect 8860 4400 8880 4410
rect 8890 4400 9200 4410
rect 9550 4400 9840 4410
rect 3010 4390 3050 4400
rect 3240 4390 3260 4400
rect 3320 4390 3360 4400
rect 5320 4390 5360 4400
rect 5800 4390 5840 4400
rect 6680 4390 7240 4400
rect 7250 4390 7270 4400
rect 7280 4390 7340 4400
rect 7370 4390 7420 4400
rect 7810 4390 7850 4400
rect 7910 4390 7990 4400
rect 8860 4390 8880 4400
rect 8890 4390 9190 4400
rect 9540 4390 9850 4400
rect 2960 4380 2970 4390
rect 3010 4380 3040 4390
rect 3250 4380 3260 4390
rect 3330 4380 3360 4390
rect 5340 4380 5370 4390
rect 5800 4380 5880 4390
rect 6680 4380 7240 4390
rect 7250 4380 7270 4390
rect 7280 4380 7300 4390
rect 7310 4380 7330 4390
rect 7370 4380 7420 4390
rect 7820 4380 7850 4390
rect 7930 4380 7970 4390
rect 8670 4380 8720 4390
rect 8860 4380 9190 4390
rect 9530 4380 9850 4390
rect 2960 4370 2970 4380
rect 3010 4370 3040 4380
rect 3060 4370 3070 4380
rect 3330 4370 3360 4380
rect 5350 4370 5370 4380
rect 5800 4370 5900 4380
rect 6680 4370 7250 4380
rect 7290 4370 7330 4380
rect 7370 4370 7420 4380
rect 7820 4370 7850 4380
rect 8660 4370 8690 4380
rect 8710 4370 8720 4380
rect 8860 4370 9190 4380
rect 9510 4370 9840 4380
rect 3000 4360 3040 4370
rect 3330 4360 3350 4370
rect 5350 4360 5380 4370
rect 5810 4360 5940 4370
rect 6670 4360 7250 4370
rect 7260 4360 7270 4370
rect 7280 4360 7330 4370
rect 7380 4360 7410 4370
rect 7820 4360 7850 4370
rect 8600 4360 8620 4370
rect 8660 4360 8670 4370
rect 8860 4360 9180 4370
rect 9500 4360 9830 4370
rect 3000 4350 3030 4360
rect 3330 4350 3340 4360
rect 5350 4350 5390 4360
rect 5820 4350 5950 4360
rect 6670 4350 7350 4360
rect 7830 4350 7840 4360
rect 8540 4350 8570 4360
rect 8600 4350 8620 4360
rect 8650 4350 8670 4360
rect 8870 4350 9180 4360
rect 9490 4350 9820 4360
rect 9980 4350 9990 4360
rect 2940 4340 2950 4350
rect 3000 4340 3020 4350
rect 3280 4340 3300 4350
rect 5350 4340 5390 4350
rect 5860 4340 5950 4350
rect 6670 4340 7240 4350
rect 7260 4340 7280 4350
rect 7290 4340 7350 4350
rect 8550 4340 8580 4350
rect 8590 4340 8610 4350
rect 8660 4340 8720 4350
rect 8870 4340 9180 4350
rect 9480 4340 9800 4350
rect 9910 4340 9950 4350
rect 9990 4340 9990 4350
rect 2940 4330 2950 4340
rect 2960 4330 2980 4340
rect 3000 4330 3020 4340
rect 3280 4330 3300 4340
rect 5350 4330 5400 4340
rect 5880 4330 5940 4340
rect 6670 4330 7350 4340
rect 8490 4330 8510 4340
rect 8560 4330 8610 4340
rect 8670 4330 8730 4340
rect 8870 4330 9180 4340
rect 9470 4330 9800 4340
rect 9860 4330 9880 4340
rect 9900 4330 9960 4340
rect 9980 4330 9990 4340
rect 2960 4320 2970 4330
rect 5350 4320 5410 4330
rect 5900 4320 5910 4330
rect 6660 4320 7340 4330
rect 8440 4320 8460 4330
rect 8490 4320 8510 4330
rect 8570 4320 8610 4330
rect 8720 4320 8740 4330
rect 8870 4320 9180 4330
rect 9460 4320 9790 4330
rect 9820 4320 9840 4330
rect 9860 4320 9880 4330
rect 9900 4320 9920 4330
rect 9970 4320 9990 4330
rect 3160 4310 3170 4320
rect 4680 4310 4780 4320
rect 5360 4310 5410 4320
rect 6660 4310 7190 4320
rect 7200 4310 7290 4320
rect 8440 4310 8470 4320
rect 8500 4310 8520 4320
rect 8580 4310 8600 4320
rect 8720 4310 8740 4320
rect 8870 4310 9180 4320
rect 9450 4310 9780 4320
rect 9810 4310 9880 4320
rect 9900 4310 9910 4320
rect 9980 4310 9990 4320
rect 2930 4300 2940 4310
rect 3230 4300 3240 4310
rect 4650 4300 4810 4310
rect 5350 4300 5420 4310
rect 6660 4300 7250 4310
rect 8440 4300 8480 4310
rect 8500 4300 8520 4310
rect 8580 4300 8600 4310
rect 8670 4300 8690 4310
rect 8720 4300 8740 4310
rect 8870 4300 9180 4310
rect 9440 4300 9770 4310
rect 9800 4300 9880 4310
rect 9900 4300 9910 4310
rect 9970 4300 9990 4310
rect 3220 4290 3240 4300
rect 4650 4290 4820 4300
rect 5350 4290 5430 4300
rect 6650 4290 7200 4300
rect 8450 4290 8490 4300
rect 8500 4290 8520 4300
rect 8590 4290 8610 4300
rect 8670 4290 8730 4300
rect 8860 4290 9180 4300
rect 9430 4290 9760 4300
rect 9800 4290 9880 4300
rect 9900 4290 9910 4300
rect 9960 4290 9990 4300
rect 3210 4280 3240 4290
rect 4610 4280 4620 4290
rect 4630 4280 4820 4290
rect 5360 4280 5430 4290
rect 6650 4280 7180 4290
rect 8450 4280 8520 4290
rect 8590 4280 8610 4290
rect 8860 4280 9180 4290
rect 9430 4280 9750 4290
rect 9800 4280 9830 4290
rect 9840 4280 9860 4290
rect 9900 4280 9910 4290
rect 9950 4280 9990 4290
rect 3210 4270 3230 4280
rect 4610 4270 4820 4280
rect 5360 4270 5390 4280
rect 5410 4270 5440 4280
rect 6650 4270 7150 4280
rect 8450 4270 8470 4280
rect 8480 4270 8530 4280
rect 8590 4270 8610 4280
rect 8860 4270 9180 4280
rect 9420 4270 9740 4280
rect 9850 4270 9860 4280
rect 9890 4270 9910 4280
rect 9940 4270 9990 4280
rect 3140 4260 3160 4270
rect 3210 4260 3230 4270
rect 4610 4260 4840 4270
rect 5370 4260 5390 4270
rect 5410 4260 5430 4270
rect 5650 4260 5660 4270
rect 6650 4260 7050 4270
rect 7070 4260 7080 4270
rect 8450 4260 8470 4270
rect 8490 4260 8530 4270
rect 8850 4260 9180 4270
rect 9410 4260 9740 4270
rect 9890 4260 9900 4270
rect 9930 4260 9990 4270
rect 3210 4250 3230 4260
rect 4610 4250 4840 4260
rect 5380 4250 5460 4260
rect 5660 4250 5670 4260
rect 6660 4250 7040 4260
rect 8450 4250 8470 4260
rect 8500 4250 8530 4260
rect 8850 4250 9180 4260
rect 9400 4250 9730 4260
rect 9820 4250 9830 4260
rect 9880 4250 9900 4260
rect 9920 4250 9990 4260
rect 3210 4240 3220 4250
rect 4600 4240 4850 4250
rect 5380 4240 5470 4250
rect 5650 4240 5690 4250
rect 6660 4240 7050 4250
rect 8460 4240 8470 4250
rect 8850 4240 9180 4250
rect 9400 4240 9730 4250
rect 9810 4240 9820 4250
rect 9880 4240 9990 4250
rect 3140 4230 3150 4240
rect 3200 4230 3220 4240
rect 4600 4230 4830 4240
rect 5380 4230 5480 4240
rect 5650 4230 5720 4240
rect 6660 4230 7090 4240
rect 8840 4230 9180 4240
rect 9390 4230 9720 4240
rect 9880 4230 9940 4240
rect 9950 4230 9970 4240
rect 3190 4220 3210 4230
rect 4600 4220 4770 4230
rect 5390 4220 5480 4230
rect 5650 4220 5720 4230
rect 6670 4220 7120 4230
rect 8840 4220 9180 4230
rect 9380 4220 9710 4230
rect 9840 4220 9860 4230
rect 9880 4220 9930 4230
rect 3050 4210 3070 4220
rect 3190 4210 3210 4220
rect 4270 4210 4280 4220
rect 4590 4210 4710 4220
rect 5400 4210 5490 4220
rect 5650 4210 5750 4220
rect 5840 4210 5910 4220
rect 6670 4210 7150 4220
rect 7210 4210 7230 4220
rect 7380 4210 7460 4220
rect 8840 4210 9180 4220
rect 9340 4210 9680 4220
rect 9830 4210 9870 4220
rect 9890 4210 9920 4220
rect 4230 4200 4300 4210
rect 5410 4200 5490 4210
rect 5660 4200 5810 4210
rect 5830 4200 5920 4210
rect 6660 4200 7230 4210
rect 7340 4200 7460 4210
rect 8830 4200 9180 4210
rect 9320 4200 9670 4210
rect 9820 4200 9880 4210
rect 9900 4200 9930 4210
rect 9950 4200 9960 4210
rect 4220 4190 4300 4200
rect 5430 4190 5490 4200
rect 5660 4190 5920 4200
rect 6670 4190 7220 4200
rect 7290 4190 7470 4200
rect 8830 4190 9180 4200
rect 9240 4190 9270 4200
rect 9320 4190 9670 4200
rect 9820 4190 9860 4200
rect 9910 4190 9980 4200
rect 9990 4190 9990 4200
rect 3150 4180 3160 4190
rect 4200 4180 4330 4190
rect 4800 4180 4820 4190
rect 4960 4180 4970 4190
rect 5420 4180 5490 4190
rect 5670 4180 5930 4190
rect 6670 4180 7230 4190
rect 7320 4180 7470 4190
rect 8830 4180 9180 4190
rect 9200 4180 9280 4190
rect 9340 4180 9670 4190
rect 9760 4180 9790 4190
rect 9900 4180 9990 4190
rect 4190 4170 4340 4180
rect 5420 4170 5490 4180
rect 5670 4170 5920 4180
rect 6670 4170 7250 4180
rect 7340 4170 7470 4180
rect 8830 4170 9280 4180
rect 9340 4170 9660 4180
rect 9700 4170 9800 4180
rect 9890 4170 9990 4180
rect 4210 4160 4340 4170
rect 5440 4160 5490 4170
rect 5680 4160 5920 4170
rect 6670 4160 7250 4170
rect 7350 4160 7470 4170
rect 8820 4160 9210 4170
rect 9230 4160 9280 4170
rect 9320 4160 9660 4170
rect 9690 4160 9790 4170
rect 9890 4160 9990 4170
rect 4180 4150 4340 4160
rect 5450 4150 5490 4160
rect 5690 4150 5940 4160
rect 6670 4150 7250 4160
rect 7370 4150 7410 4160
rect 8820 4150 9260 4160
rect 9320 4150 9650 4160
rect 9680 4150 9780 4160
rect 9900 4150 9990 4160
rect 3270 4140 3280 4150
rect 4190 4140 4350 4150
rect 5460 4140 5490 4150
rect 5690 4140 5950 4150
rect 6670 4140 7250 4150
rect 8820 4140 9280 4150
rect 9300 4140 9630 4150
rect 9670 4140 9800 4150
rect 9920 4140 9940 4150
rect 3260 4130 3270 4140
rect 4180 4130 4350 4140
rect 5460 4130 5490 4140
rect 5700 4130 5950 4140
rect 6670 4130 7240 4140
rect 8820 4130 9630 4140
rect 9660 4130 9820 4140
rect 3260 4120 3270 4130
rect 4170 4120 4390 4130
rect 4400 4120 4410 4130
rect 5460 4120 5490 4130
rect 5710 4120 5950 4130
rect 6670 4120 7240 4130
rect 8810 4120 9630 4130
rect 9660 4120 9820 4130
rect 3240 4110 3260 4120
rect 4170 4110 4420 4120
rect 5470 4110 5490 4120
rect 5710 4110 5950 4120
rect 6480 4110 6490 4120
rect 6660 4110 7240 4120
rect 8810 4110 9630 4120
rect 9650 4110 9770 4120
rect 9780 4110 9800 4120
rect 3220 4100 3240 4110
rect 3250 4100 3270 4110
rect 4160 4100 4440 4110
rect 5460 4100 5490 4110
rect 5720 4100 5730 4110
rect 5780 4100 5950 4110
rect 6470 4100 6490 4110
rect 6660 4100 7230 4110
rect 8810 4100 9620 4110
rect 9640 4100 9760 4110
rect 9990 4100 9990 4110
rect 3210 4090 3260 4100
rect 4160 4090 4440 4100
rect 5020 4090 5030 4100
rect 5470 4090 5500 4100
rect 5800 4090 5960 4100
rect 6460 4090 6490 4100
rect 6650 4090 7230 4100
rect 8810 4090 9210 4100
rect 9220 4090 9610 4100
rect 9650 4090 9710 4100
rect 3220 4080 3240 4090
rect 4120 4080 4140 4090
rect 4160 4080 4440 4090
rect 4930 4080 5030 4090
rect 5450 4080 5460 4090
rect 5470 4080 5490 4090
rect 5810 4080 5960 4090
rect 6460 4080 6490 4090
rect 6650 4080 7220 4090
rect 8800 4080 9200 4090
rect 9220 4080 9600 4090
rect 9840 4080 9890 4090
rect 3130 4070 3180 4080
rect 3220 4070 3240 4080
rect 4120 4070 4440 4080
rect 4840 4070 4870 4080
rect 4910 4070 5030 4080
rect 5440 4070 5490 4080
rect 5840 4070 5910 4080
rect 5920 4070 5930 4080
rect 5940 4070 5950 4080
rect 6460 4070 6490 4080
rect 6650 4070 7220 4080
rect 8800 4070 9200 4080
rect 9220 4070 9600 4080
rect 9620 4070 9630 4080
rect 9760 4070 9770 4080
rect 9790 4070 9910 4080
rect 3150 4060 3180 4070
rect 3220 4060 3240 4070
rect 4130 4060 4210 4070
rect 4220 4060 4450 4070
rect 4830 4060 4880 4070
rect 4900 4060 5020 4070
rect 5430 4060 5490 4070
rect 6470 4060 6490 4070
rect 6540 4060 6560 4070
rect 6660 4060 6680 4070
rect 6700 4060 7210 4070
rect 8800 4060 9210 4070
rect 9220 4060 9590 4070
rect 9610 4060 9660 4070
rect 9730 4060 9930 4070
rect 3070 4050 3090 4060
rect 3220 4050 3240 4060
rect 4130 4050 4170 4060
rect 4180 4050 4200 4060
rect 4250 4050 4470 4060
rect 4810 4050 4870 4060
rect 4900 4050 5030 4060
rect 5040 4050 5050 4060
rect 5430 4050 5490 4060
rect 6470 4050 6490 4060
rect 6550 4050 6570 4060
rect 6690 4050 7200 4060
rect 7640 4050 7650 4060
rect 8630 4050 8650 4060
rect 8790 4050 9210 4060
rect 9220 4050 9580 4060
rect 9600 4050 9950 4060
rect 3100 4040 3110 4050
rect 3180 4040 3200 4050
rect 3230 4040 3240 4050
rect 3250 4040 3270 4050
rect 4100 4040 4170 4050
rect 4270 4040 4290 4050
rect 4300 4040 4470 4050
rect 4800 4040 4870 4050
rect 4900 4040 5040 4050
rect 5430 4040 5490 4050
rect 6480 4040 6490 4050
rect 6540 4040 6570 4050
rect 6670 4040 7190 4050
rect 7670 4040 7680 4050
rect 8640 4040 8660 4050
rect 8790 4040 9210 4050
rect 9220 4040 9570 4050
rect 9590 4040 9970 4050
rect 3230 4030 3240 4040
rect 3260 4030 3270 4040
rect 4090 4030 4170 4040
rect 4310 4030 4480 4040
rect 4780 4030 4860 4040
rect 4910 4030 5030 4040
rect 5430 4030 5490 4040
rect 6480 4030 6490 4040
rect 6540 4030 6590 4040
rect 6650 4030 7180 4040
rect 8650 4030 8660 4040
rect 8780 4030 9560 4040
rect 9580 4030 9990 4040
rect 3230 4020 3240 4030
rect 4080 4020 4150 4030
rect 4170 4020 4180 4030
rect 4320 4020 4480 4030
rect 4770 4020 4830 4030
rect 4910 4020 5010 4030
rect 5430 4020 5490 4030
rect 6630 4020 7160 4030
rect 8540 4020 8560 4030
rect 8780 4020 9560 4030
rect 9570 4020 9990 4030
rect 3230 4010 3240 4020
rect 3260 4010 3270 4020
rect 4070 4010 4170 4020
rect 4330 4010 4500 4020
rect 4750 4010 4820 4020
rect 4900 4010 5020 4020
rect 5430 4010 5490 4020
rect 6610 4010 7010 4020
rect 7020 4010 7130 4020
rect 7150 4010 7160 4020
rect 7740 4010 7750 4020
rect 8550 4010 8570 4020
rect 8610 4010 8640 4020
rect 8780 4010 9550 4020
rect 9560 4010 9990 4020
rect 3200 4000 3210 4010
rect 3230 4000 3240 4010
rect 3260 4000 3270 4010
rect 4070 4000 4160 4010
rect 4330 4000 4500 4010
rect 4720 4000 4790 4010
rect 4890 4000 5020 4010
rect 5420 4000 5490 4010
rect 6580 4000 7010 4010
rect 7030 4000 7140 4010
rect 8440 4000 8470 4010
rect 8570 4000 8580 4010
rect 8620 4000 8640 4010
rect 8770 4000 9990 4010
rect 3230 3990 3240 4000
rect 4070 3990 4150 4000
rect 4340 3990 4500 4000
rect 4700 3990 4770 4000
rect 4880 3990 5060 4000
rect 5420 3990 5490 4000
rect 6580 3990 7020 4000
rect 7030 3990 7130 4000
rect 8360 3990 8400 4000
rect 8440 3990 8480 4000
rect 8570 3990 8620 4000
rect 8770 3990 9990 4000
rect 3150 3980 3170 3990
rect 3230 3980 3240 3990
rect 4050 3980 4140 3990
rect 4350 3980 4510 3990
rect 4680 3980 4710 3990
rect 4730 3980 4740 3990
rect 4860 3980 5070 3990
rect 5410 3980 5450 3990
rect 5470 3980 5480 3990
rect 6580 3980 7020 3990
rect 7030 3980 7130 3990
rect 7820 3980 7830 3990
rect 8340 3980 8400 3990
rect 8460 3980 8490 3990
rect 8570 3980 8620 3990
rect 8760 3980 9990 3990
rect 3150 3970 3160 3980
rect 3230 3970 3240 3980
rect 4050 3970 4130 3980
rect 4350 3970 4520 3980
rect 4850 3970 5080 3980
rect 6580 3970 7020 3980
rect 7040 3970 7120 3980
rect 8330 3970 8400 3980
rect 8480 3970 8500 3980
rect 8580 3970 8630 3980
rect 8680 3970 8700 3980
rect 8750 3970 9990 3980
rect 3150 3960 3160 3970
rect 3210 3960 3250 3970
rect 4040 3960 4120 3970
rect 4350 3960 4520 3970
rect 4650 3960 4660 3970
rect 4830 3960 5100 3970
rect 6580 3960 7020 3970
rect 7040 3960 7110 3970
rect 7870 3960 7880 3970
rect 8240 3960 8270 3970
rect 8340 3960 8410 3970
rect 8490 3960 8510 3970
rect 8580 3960 8650 3970
rect 8750 3960 9990 3970
rect 3230 3950 3250 3960
rect 4030 3950 4100 3960
rect 4350 3950 4530 3960
rect 4650 3950 4660 3960
rect 4810 3950 5100 3960
rect 6580 3950 7110 3960
rect 8250 3950 8290 3960
rect 8340 3950 8410 3960
rect 8450 3950 8480 3960
rect 8490 3950 8500 3960
rect 8580 3950 8660 3960
rect 8670 3950 8680 3960
rect 8720 3950 8730 3960
rect 8750 3950 9670 3960
rect 9710 3950 9990 3960
rect 3230 3940 3240 3950
rect 4010 3940 4100 3950
rect 4350 3940 4530 3950
rect 4810 3940 5120 3950
rect 6590 3940 7110 3950
rect 8270 3940 8320 3950
rect 8340 3940 8410 3950
rect 8460 3940 8500 3950
rect 8580 3940 8640 3950
rect 8670 3940 8680 3950
rect 8720 3940 9650 3950
rect 9730 3940 9990 3950
rect 3230 3930 3240 3940
rect 4000 3930 4080 3940
rect 4360 3930 4530 3940
rect 4780 3930 5130 3940
rect 6590 3930 7120 3940
rect 8210 3930 8240 3940
rect 8290 3930 8320 3940
rect 8350 3930 8410 3940
rect 8470 3930 8500 3940
rect 8590 3930 8630 3940
rect 8730 3930 9640 3940
rect 9750 3930 9990 3940
rect 3230 3920 3240 3930
rect 3250 3920 3260 3930
rect 3980 3920 4070 3930
rect 4360 3920 4530 3930
rect 4740 3920 5140 3930
rect 6590 3920 7140 3930
rect 8210 3920 8250 3930
rect 8300 3920 8330 3930
rect 8340 3920 8430 3930
rect 8470 3920 8510 3930
rect 8710 3920 9610 3930
rect 9760 3920 9940 3930
rect 9950 3920 9990 3930
rect 3970 3910 4060 3920
rect 4370 3910 4530 3920
rect 4660 3910 4670 3920
rect 4680 3910 4690 3920
rect 4700 3910 5130 3920
rect 6600 3910 7140 3920
rect 8010 3910 8050 3920
rect 8210 3910 8260 3920
rect 8320 3910 8480 3920
rect 8500 3910 8510 3920
rect 8710 3910 9600 3920
rect 9780 3910 9990 3920
rect 3240 3900 3270 3910
rect 3970 3900 4050 3910
rect 4380 3900 4540 3910
rect 4630 3900 5140 3910
rect 6600 3900 7140 3910
rect 7990 3900 8060 3910
rect 8200 3900 8260 3910
rect 8340 3900 8480 3910
rect 8500 3900 8510 3910
rect 8720 3900 9600 3910
rect 9790 3900 9990 3910
rect 3220 3890 3270 3900
rect 3950 3890 4020 3900
rect 4380 3890 4540 3900
rect 4640 3890 5150 3900
rect 6600 3890 7130 3900
rect 8010 3890 8060 3900
rect 8200 3890 8270 3900
rect 8350 3890 8420 3900
rect 8470 3890 8510 3900
rect 8720 3890 9490 3900
rect 9500 3890 9550 3900
rect 9770 3890 9990 3900
rect 3220 3880 3270 3890
rect 3950 3880 4000 3890
rect 4390 3880 4550 3890
rect 4640 3880 5150 3890
rect 6600 3880 7130 3890
rect 8020 3880 8050 3890
rect 8210 3880 8270 3890
rect 8350 3880 8420 3890
rect 8480 3880 8510 3890
rect 8620 3880 8630 3890
rect 8700 3880 9460 3890
rect 9730 3880 9800 3890
rect 9820 3880 9990 3890
rect 3180 3870 3200 3880
rect 3210 3870 3270 3880
rect 3940 3870 3990 3880
rect 4390 3870 4550 3880
rect 4650 3870 5160 3880
rect 6600 3870 7120 3880
rect 8230 3870 8280 3880
rect 8350 3870 8420 3880
rect 8490 3870 8520 3880
rect 8700 3870 9440 3880
rect 9730 3870 9790 3880
rect 9840 3870 9990 3880
rect 3130 3860 3140 3870
rect 3190 3860 3200 3870
rect 3220 3860 3260 3870
rect 3930 3860 3980 3870
rect 4400 3860 4550 3870
rect 4640 3860 5160 3870
rect 6610 3860 7120 3870
rect 8240 3860 8290 3870
rect 8360 3860 8420 3870
rect 8480 3860 8530 3870
rect 8580 3860 8610 3870
rect 8650 3860 8660 3870
rect 8700 3860 9430 3870
rect 9730 3860 9770 3870
rect 9860 3860 9990 3870
rect 3200 3850 3260 3860
rect 3920 3850 3970 3860
rect 4400 3850 4580 3860
rect 4640 3850 5160 3860
rect 6610 3850 7110 3860
rect 8250 3850 8310 3860
rect 8370 3850 8430 3860
rect 8470 3850 8550 3860
rect 8590 3850 8610 3860
rect 8650 3850 8670 3860
rect 8700 3850 9430 3860
rect 9480 3850 9550 3860
rect 9740 3850 9800 3860
rect 9870 3850 9990 3860
rect 3190 3840 3260 3850
rect 3920 3840 3960 3850
rect 4410 3840 4590 3850
rect 4640 3840 5160 3850
rect 6610 3840 7110 3850
rect 8260 3840 8320 3850
rect 8410 3840 8460 3850
rect 8480 3840 8520 3850
rect 8530 3840 8570 3850
rect 8620 3840 8630 3850
rect 8680 3840 9430 3850
rect 9440 3840 9580 3850
rect 9740 3840 9800 3850
rect 9890 3840 9990 3850
rect 3170 3830 3240 3840
rect 3250 3830 3260 3840
rect 3920 3830 3950 3840
rect 4410 3830 4600 3840
rect 4650 3830 5160 3840
rect 6610 3830 7100 3840
rect 8270 3830 8340 3840
rect 8410 3830 8460 3840
rect 8500 3830 8530 3840
rect 8550 3830 8590 3840
rect 8690 3830 9590 3840
rect 9740 3830 9800 3840
rect 9870 3830 9890 3840
rect 9900 3830 9990 3840
rect 3210 3820 3250 3830
rect 3920 3820 3950 3830
rect 4410 3820 4610 3830
rect 4650 3820 5160 3830
rect 6610 3820 7090 3830
rect 8270 3820 8350 3830
rect 8420 3820 8430 3830
rect 8450 3820 8480 3830
rect 8510 3820 8550 3830
rect 8560 3820 8590 3830
rect 8660 3820 8670 3830
rect 8690 3820 9600 3830
rect 9750 3820 9790 3830
rect 9830 3820 9990 3830
rect 3210 3810 3250 3820
rect 3920 3810 3940 3820
rect 4420 3810 5160 3820
rect 6610 3810 7090 3820
rect 8260 3810 8290 3820
rect 8320 3810 8360 3820
rect 8470 3810 8490 3820
rect 8530 3810 8610 3820
rect 8650 3810 8670 3820
rect 8680 3810 9600 3820
rect 9820 3810 9990 3820
rect 3210 3800 3250 3810
rect 4430 3800 5160 3810
rect 6610 3800 7080 3810
rect 8330 3800 8380 3810
rect 8480 3800 8510 3810
rect 8540 3800 8620 3810
rect 8670 3800 9610 3810
rect 9830 3800 9990 3810
rect 3200 3790 3240 3800
rect 4440 3790 5160 3800
rect 6610 3790 7070 3800
rect 8120 3790 8140 3800
rect 8360 3790 8380 3800
rect 8490 3790 8520 3800
rect 8540 3790 8640 3800
rect 8670 3790 9610 3800
rect 9840 3790 9990 3800
rect 3200 3780 3210 3790
rect 3230 3780 3260 3790
rect 4270 3780 4300 3790
rect 4450 3780 5150 3790
rect 6610 3780 7060 3790
rect 8130 3780 8140 3790
rect 8370 3780 8420 3790
rect 8430 3780 8450 3790
rect 8510 3780 8640 3790
rect 8670 3780 9620 3790
rect 9750 3780 9770 3790
rect 9850 3780 9990 3790
rect 2950 3770 2970 3780
rect 3200 3770 3230 3780
rect 3250 3770 3260 3780
rect 4450 3770 4870 3780
rect 4900 3770 5150 3780
rect 6610 3770 7060 3780
rect 8380 3770 8480 3780
rect 8530 3770 8630 3780
rect 8660 3770 9640 3780
rect 9750 3770 9760 3780
rect 9890 3770 9990 3780
rect 3200 3760 3260 3770
rect 4210 3760 4220 3770
rect 4450 3760 4840 3770
rect 4930 3760 5150 3770
rect 6610 3760 7050 3770
rect 8390 3760 8490 3770
rect 8540 3760 8630 3770
rect 8660 3760 9650 3770
rect 9870 3760 9900 3770
rect 9910 3760 9990 3770
rect 3240 3750 3270 3760
rect 4160 3750 4200 3760
rect 4450 3750 4810 3760
rect 4950 3750 5140 3760
rect 6610 3750 7040 3760
rect 8160 3750 8170 3760
rect 8400 3750 8510 3760
rect 8550 3750 8640 3760
rect 8650 3750 9660 3760
rect 9800 3750 9820 3760
rect 9870 3750 9990 3760
rect 3190 3740 3200 3750
rect 3250 3740 3260 3750
rect 4110 3740 4180 3750
rect 4440 3740 4780 3750
rect 4970 3740 5130 3750
rect 6610 3740 7040 3750
rect 8410 3740 8520 3750
rect 8570 3740 9670 3750
rect 9800 3740 9820 3750
rect 9880 3740 9990 3750
rect 2960 3730 2990 3740
rect 3190 3730 3230 3740
rect 4090 3730 4160 3740
rect 4440 3730 4780 3740
rect 4990 3730 5110 3740
rect 6610 3730 7030 3740
rect 8430 3730 8530 3740
rect 8580 3730 9680 3740
rect 9850 3730 9870 3740
rect 9900 3730 9920 3740
rect 9990 3730 9990 3740
rect 3180 3720 3220 3730
rect 3260 3720 3270 3730
rect 4070 3720 4140 3730
rect 4440 3720 4780 3730
rect 5060 3720 5080 3730
rect 6610 3720 7020 3730
rect 8440 3720 8530 3730
rect 8600 3720 9690 3730
rect 9830 3720 9870 3730
rect 9990 3720 9990 3730
rect 3030 3710 3040 3720
rect 3250 3710 3270 3720
rect 4060 3710 4130 3720
rect 4450 3710 4780 3720
rect 6610 3710 7020 3720
rect 8190 3710 8210 3720
rect 8350 3710 8370 3720
rect 8460 3710 8540 3720
rect 8610 3710 9600 3720
rect 9610 3710 9690 3720
rect 9710 3710 9720 3720
rect 9730 3710 9870 3720
rect 9990 3710 9990 3720
rect 3090 3700 3110 3710
rect 3180 3700 3190 3710
rect 3260 3700 3280 3710
rect 4050 3700 4080 3710
rect 4440 3700 4810 3710
rect 6610 3700 7010 3710
rect 8200 3700 8220 3710
rect 8270 3700 8290 3710
rect 8350 3700 8370 3710
rect 8470 3700 8550 3710
rect 8620 3700 9560 3710
rect 9570 3700 9590 3710
rect 9620 3700 9870 3710
rect 9970 3700 9990 3710
rect 3090 3690 3170 3700
rect 3270 3690 3280 3700
rect 4050 3690 4070 3700
rect 4260 3690 4280 3700
rect 4450 3690 4810 3700
rect 6600 3690 7000 3700
rect 8210 3690 8320 3700
rect 8330 3690 8370 3700
rect 8490 3690 8550 3700
rect 8620 3690 9540 3700
rect 9570 3690 9590 3700
rect 9630 3690 9830 3700
rect 9840 3690 9860 3700
rect 9970 3690 9990 3700
rect 3110 3680 3180 3690
rect 3260 3680 3290 3690
rect 4040 3680 4060 3690
rect 4230 3680 4310 3690
rect 4440 3680 4810 3690
rect 6600 3680 6990 3690
rect 8210 3680 8320 3690
rect 8330 3680 8360 3690
rect 8380 3680 8390 3690
rect 8500 3680 8550 3690
rect 8620 3680 9520 3690
rect 9550 3680 9580 3690
rect 9640 3680 9830 3690
rect 9930 3680 9990 3690
rect 3110 3670 3120 3680
rect 3140 3670 3170 3680
rect 3260 3670 3280 3680
rect 4220 3670 4320 3680
rect 4450 3670 4810 3680
rect 6600 3670 6980 3680
rect 8210 3670 8390 3680
rect 8520 3670 8560 3680
rect 8610 3670 9510 3680
rect 9520 3670 9570 3680
rect 9650 3670 9840 3680
rect 9930 3670 9990 3680
rect 3170 3660 3180 3670
rect 4180 3660 4320 3670
rect 4440 3660 4810 3670
rect 6600 3660 6960 3670
rect 8210 3660 8400 3670
rect 8530 3660 8560 3670
rect 8610 3660 9570 3670
rect 9660 3660 9850 3670
rect 9890 3660 9990 3670
rect 4100 3650 4340 3660
rect 4440 3650 4810 3660
rect 6600 3650 6960 3660
rect 8220 3650 8310 3660
rect 8320 3650 8350 3660
rect 8370 3650 8380 3660
rect 8390 3650 8400 3660
rect 8560 3650 9550 3660
rect 9680 3650 9870 3660
rect 9890 3650 9930 3660
rect 9940 3650 9990 3660
rect 3150 3640 3170 3650
rect 4050 3640 4340 3650
rect 4420 3640 4810 3650
rect 4840 3640 4870 3650
rect 6590 3640 6950 3650
rect 8230 3640 8320 3650
rect 8570 3640 9530 3650
rect 9680 3640 9870 3650
rect 9900 3640 9990 3650
rect 4040 3630 4330 3640
rect 4400 3630 4800 3640
rect 4850 3630 4870 3640
rect 6600 3630 6950 3640
rect 8250 3630 8340 3640
rect 8520 3630 8530 3640
rect 8560 3630 9520 3640
rect 9690 3630 9860 3640
rect 9920 3630 9990 3640
rect 3190 3620 3200 3630
rect 4040 3620 4270 3630
rect 4280 3620 4330 3630
rect 4420 3620 4800 3630
rect 6590 3620 6940 3630
rect 8260 3620 8340 3630
rect 8560 3620 9510 3630
rect 9690 3620 9820 3630
rect 9860 3620 9900 3630
rect 9950 3620 9990 3630
rect 4050 3610 4340 3620
rect 4430 3610 4800 3620
rect 6590 3610 6930 3620
rect 8270 3610 8340 3620
rect 8530 3610 9500 3620
rect 9700 3610 9910 3620
rect 9950 3610 9990 3620
rect 4050 3600 4340 3610
rect 4440 3600 4780 3610
rect 4850 3600 4880 3610
rect 6590 3600 6930 3610
rect 8270 3600 8340 3610
rect 8530 3600 9460 3610
rect 9700 3600 9910 3610
rect 9950 3600 9990 3610
rect 3350 3590 3370 3600
rect 4060 3590 4340 3600
rect 4450 3590 4730 3600
rect 4740 3590 4760 3600
rect 4850 3590 4910 3600
rect 6590 3590 6920 3600
rect 8290 3590 8340 3600
rect 8510 3590 9440 3600
rect 9580 3590 9610 3600
rect 9690 3590 9750 3600
rect 9760 3590 9920 3600
rect 9940 3590 9990 3600
rect 4060 3580 4310 3590
rect 4330 3580 4350 3590
rect 4470 3580 4700 3590
rect 4850 3580 4920 3590
rect 4930 3580 4970 3590
rect 6580 3580 6910 3590
rect 8310 3580 8330 3590
rect 8350 3580 8360 3590
rect 8370 3580 8380 3590
rect 8510 3580 9300 3590
rect 9370 3580 9380 3590
rect 9390 3580 9400 3590
rect 9410 3580 9420 3590
rect 9560 3580 9630 3590
rect 9680 3580 9730 3590
rect 9760 3580 9990 3590
rect 3290 3570 3320 3580
rect 3360 3570 3370 3580
rect 4060 3570 4310 3580
rect 4470 3570 4690 3580
rect 4850 3570 4990 3580
rect 6580 3570 6900 3580
rect 8320 3570 8360 3580
rect 8510 3570 9260 3580
rect 9550 3570 9630 3580
rect 9680 3570 9720 3580
rect 9750 3570 9990 3580
rect 3290 3560 3310 3570
rect 3360 3560 3370 3570
rect 4050 3560 4290 3570
rect 4480 3560 4680 3570
rect 4840 3560 4990 3570
rect 6580 3560 6900 3570
rect 8320 3560 8370 3570
rect 8510 3560 8820 3570
rect 8830 3560 9250 3570
rect 9540 3560 9630 3570
rect 9670 3560 9720 3570
rect 9740 3560 9990 3570
rect 3280 3550 3330 3560
rect 3360 3550 3380 3560
rect 4040 3550 4280 3560
rect 4490 3550 4670 3560
rect 4840 3550 5000 3560
rect 6580 3550 6890 3560
rect 8340 3550 8380 3560
rect 8400 3550 8410 3560
rect 8510 3550 9230 3560
rect 9530 3550 9630 3560
rect 9670 3550 9710 3560
rect 9720 3550 9990 3560
rect 3290 3540 3330 3550
rect 3370 3540 3380 3550
rect 4050 3540 4270 3550
rect 4490 3540 4650 3550
rect 4830 3540 5010 3550
rect 6590 3540 6870 3550
rect 8340 3540 8410 3550
rect 8500 3540 9210 3550
rect 9520 3540 9630 3550
rect 9690 3540 9990 3550
rect 3310 3530 3340 3540
rect 3370 3530 3390 3540
rect 4050 3530 4260 3540
rect 4490 3530 4630 3540
rect 4830 3530 5000 3540
rect 6580 3530 6870 3540
rect 8350 3530 8390 3540
rect 8500 3530 9180 3540
rect 9500 3530 9620 3540
rect 9670 3530 9990 3540
rect 3330 3520 3350 3530
rect 3360 3520 3370 3530
rect 3380 3520 3390 3530
rect 4050 3520 4260 3530
rect 4500 3520 4600 3530
rect 4830 3520 5000 3530
rect 6580 3520 6860 3530
rect 8360 3520 8380 3530
rect 8500 3520 9180 3530
rect 9480 3520 9590 3530
rect 9660 3520 9990 3530
rect 3340 3510 3390 3520
rect 4060 3510 4240 3520
rect 4530 3510 4570 3520
rect 4820 3510 4990 3520
rect 6580 3510 6850 3520
rect 8370 3510 8410 3520
rect 8500 3510 9170 3520
rect 9460 3510 9570 3520
rect 9660 3510 9990 3520
rect 3350 3500 3380 3510
rect 3390 3500 3400 3510
rect 4070 3500 4220 3510
rect 4820 3500 4980 3510
rect 6580 3500 6850 3510
rect 8390 3500 8410 3510
rect 8510 3500 9150 3510
rect 9430 3500 9570 3510
rect 9640 3500 9990 3510
rect 3370 3490 3390 3500
rect 4070 3490 4210 3500
rect 4810 3490 4960 3500
rect 6580 3490 6830 3500
rect 8400 3490 8410 3500
rect 8520 3490 9150 3500
rect 9410 3490 9550 3500
rect 9640 3490 9990 3500
rect 2480 3480 2510 3490
rect 2530 3480 2600 3490
rect 2610 3480 2620 3490
rect 2640 3480 2650 3490
rect 2660 3480 2670 3490
rect 3380 3480 3410 3490
rect 4070 3480 4210 3490
rect 4810 3480 4950 3490
rect 6570 3480 6830 3490
rect 8420 3480 8440 3490
rect 8530 3480 9130 3490
rect 9400 3480 9540 3490
rect 9640 3480 9990 3490
rect 2420 3470 2680 3480
rect 3390 3470 3410 3480
rect 4070 3470 4200 3480
rect 4800 3470 4930 3480
rect 6570 3470 6820 3480
rect 8430 3470 8450 3480
rect 8550 3470 9120 3480
rect 9410 3470 9530 3480
rect 9640 3470 9990 3480
rect 2410 3460 2710 3470
rect 3420 3460 3430 3470
rect 4070 3460 4190 3470
rect 4800 3460 4910 3470
rect 5050 3460 5090 3470
rect 6570 3460 6820 3470
rect 8460 3460 8470 3470
rect 8560 3460 9100 3470
rect 9330 3460 9380 3470
rect 9430 3460 9480 3470
rect 9490 3460 9500 3470
rect 9630 3460 9990 3470
rect 2370 3450 2720 3460
rect 2740 3450 2750 3460
rect 2760 3450 2800 3460
rect 4080 3450 4170 3460
rect 4790 3450 4880 3460
rect 5040 3450 5110 3460
rect 6570 3450 6800 3460
rect 8470 3450 8480 3460
rect 8550 3450 9090 3460
rect 9300 3450 9420 3460
rect 9640 3450 9990 3460
rect 2350 3440 2740 3450
rect 2750 3440 2830 3450
rect 4080 3440 4150 3450
rect 4790 3440 4850 3450
rect 5040 3440 5120 3450
rect 5150 3440 5170 3450
rect 6560 3440 6800 3450
rect 8550 3440 9080 3450
rect 9280 3440 9430 3450
rect 9610 3440 9990 3450
rect 2310 3430 2740 3440
rect 2750 3430 2870 3440
rect 4080 3430 4140 3440
rect 4780 3430 4830 3440
rect 5030 3430 5120 3440
rect 5150 3430 5180 3440
rect 6560 3430 6780 3440
rect 8550 3430 9070 3440
rect 9260 3430 9430 3440
rect 9600 3430 9990 3440
rect 2290 3420 2880 3430
rect 4090 3420 4120 3430
rect 5030 3420 5120 3430
rect 5150 3420 5180 3430
rect 6550 3420 6780 3430
rect 8550 3420 9040 3430
rect 9240 3420 9420 3430
rect 9590 3420 9990 3430
rect 2280 3410 2900 3420
rect 5030 3410 5130 3420
rect 5150 3410 5180 3420
rect 6550 3410 6760 3420
rect 8550 3410 9030 3420
rect 9230 3410 9400 3420
rect 9580 3410 9650 3420
rect 9670 3410 9990 3420
rect 2260 3400 2880 3410
rect 5020 3400 5130 3410
rect 5150 3400 5180 3410
rect 6540 3400 6750 3410
rect 8530 3400 9020 3410
rect 9220 3400 9400 3410
rect 9570 3400 9650 3410
rect 9700 3400 9770 3410
rect 9780 3400 9990 3410
rect 2250 3390 2810 3400
rect 2830 3390 2920 3400
rect 5020 3390 5130 3400
rect 5150 3390 5190 3400
rect 6530 3390 6740 3400
rect 8540 3390 9010 3400
rect 9200 3390 9400 3400
rect 9560 3390 9650 3400
rect 9700 3390 9990 3400
rect 2240 3380 2980 3390
rect 4940 3380 4950 3390
rect 5020 3380 5140 3390
rect 5150 3380 5190 3390
rect 6530 3380 6730 3390
rect 8540 3380 9020 3390
rect 9190 3380 9400 3390
rect 9550 3380 9650 3390
rect 9710 3380 9760 3390
rect 9770 3380 9990 3390
rect 2230 3370 3010 3380
rect 4930 3370 4960 3380
rect 5020 3370 5140 3380
rect 5150 3370 5190 3380
rect 6520 3370 6720 3380
rect 8530 3370 9030 3380
rect 9180 3370 9410 3380
rect 9540 3370 9660 3380
rect 9700 3370 9740 3380
rect 9830 3370 9990 3380
rect 2210 3360 3030 3370
rect 3530 3360 3550 3370
rect 4930 3360 4950 3370
rect 5020 3360 5190 3370
rect 6520 3360 6710 3370
rect 8530 3360 9060 3370
rect 9170 3360 9410 3370
rect 9530 3360 9660 3370
rect 9720 3360 9730 3370
rect 9820 3360 9990 3370
rect 2200 3350 3050 3360
rect 3530 3350 3560 3360
rect 4430 3350 4450 3360
rect 4930 3350 4940 3360
rect 5020 3350 5190 3360
rect 6520 3350 6690 3360
rect 8530 3350 9060 3360
rect 9160 3350 9410 3360
rect 9520 3350 9650 3360
rect 9810 3350 9990 3360
rect 2190 3340 3060 3350
rect 3530 3340 3570 3350
rect 4420 3340 4480 3350
rect 4930 3340 4940 3350
rect 5020 3340 5190 3350
rect 6520 3340 6680 3350
rect 8520 3340 9040 3350
rect 9150 3340 9400 3350
rect 9510 3340 9640 3350
rect 9800 3340 9990 3350
rect 2180 3330 3070 3340
rect 3540 3330 3580 3340
rect 4410 3330 4500 3340
rect 4530 3330 4540 3340
rect 4930 3330 4940 3340
rect 5020 3330 5190 3340
rect 6510 3330 6660 3340
rect 8520 3330 8980 3340
rect 9140 3330 9330 3340
rect 9500 3330 9640 3340
rect 9790 3330 9990 3340
rect 2180 3320 3080 3330
rect 3540 3320 3590 3330
rect 4410 3320 4530 3330
rect 4920 3320 4940 3330
rect 5020 3320 5190 3330
rect 6510 3320 6650 3330
rect 8520 3320 8940 3330
rect 9130 3320 9330 3330
rect 9500 3320 9630 3330
rect 9780 3320 9990 3330
rect 2180 3310 3090 3320
rect 3550 3310 3590 3320
rect 4390 3310 4510 3320
rect 5020 3310 5190 3320
rect 6520 3310 6640 3320
rect 8520 3310 8920 3320
rect 9010 3310 9020 3320
rect 9130 3310 9330 3320
rect 9490 3310 9630 3320
rect 9770 3310 9990 3320
rect 2170 3300 3100 3310
rect 4400 3300 4490 3310
rect 4920 3300 4930 3310
rect 5020 3300 5200 3310
rect 6530 3300 6630 3310
rect 8480 3300 8490 3310
rect 8510 3300 8920 3310
rect 8970 3300 9020 3310
rect 9120 3300 9330 3310
rect 9490 3300 9610 3310
rect 9760 3300 9990 3310
rect 2170 3290 3110 3300
rect 4400 3290 4410 3300
rect 4420 3290 4440 3300
rect 4910 3290 4930 3300
rect 5010 3290 5200 3300
rect 6520 3290 6600 3300
rect 8480 3290 8920 3300
rect 9120 3290 9330 3300
rect 9470 3290 9600 3300
rect 9760 3290 9990 3300
rect 2150 3280 3110 3290
rect 4900 3280 4920 3290
rect 5010 3280 5200 3290
rect 6530 3280 6580 3290
rect 8480 3280 8860 3290
rect 9120 3280 9330 3290
rect 9460 3280 9590 3290
rect 9750 3280 9990 3290
rect 2150 3270 3120 3280
rect 4900 3270 4920 3280
rect 5010 3270 5200 3280
rect 6520 3270 6560 3280
rect 8500 3270 8830 3280
rect 9080 3270 9090 3280
rect 9120 3270 9320 3280
rect 9460 3270 9560 3280
rect 9740 3270 9980 3280
rect 2140 3260 3120 3270
rect 4900 3260 4920 3270
rect 5010 3260 5200 3270
rect 6520 3260 6540 3270
rect 8470 3260 8480 3270
rect 8510 3260 8820 3270
rect 8900 3260 8910 3270
rect 8930 3260 8990 3270
rect 9060 3260 9090 3270
rect 9130 3260 9310 3270
rect 9460 3260 9520 3270
rect 9730 3260 9970 3270
rect 2130 3250 3130 3260
rect 4900 3250 4910 3260
rect 5010 3250 5200 3260
rect 8460 3250 8830 3260
rect 8890 3250 8990 3260
rect 9040 3250 9090 3260
rect 9130 3250 9300 3260
rect 9720 3250 9960 3260
rect 2130 3240 3130 3250
rect 3590 3240 3610 3250
rect 4890 3240 4900 3250
rect 5000 3240 5200 3250
rect 8460 3240 8830 3250
rect 8850 3240 8990 3250
rect 9020 3240 9080 3250
rect 9150 3240 9290 3250
rect 9710 3240 9950 3250
rect 2140 3230 3140 3240
rect 3580 3230 3610 3240
rect 5000 3230 5200 3240
rect 8450 3230 8980 3240
rect 9010 3230 9080 3240
rect 9170 3230 9280 3240
rect 9620 3230 9630 3240
rect 9670 3230 9940 3240
rect 2140 3220 3140 3230
rect 3580 3220 3600 3230
rect 5000 3220 5210 3230
rect 8450 3220 8950 3230
rect 8990 3220 9070 3230
rect 9250 3220 9270 3230
rect 9610 3220 9640 3230
rect 9660 3220 9940 3230
rect 9980 3220 9990 3230
rect 2140 3210 3150 3220
rect 5000 3210 5210 3220
rect 8440 3210 8920 3220
rect 8970 3210 9060 3220
rect 9600 3210 9930 3220
rect 9980 3210 9990 3220
rect 2130 3200 3150 3210
rect 5000 3200 5210 3210
rect 8440 3200 8860 3210
rect 8940 3200 9040 3210
rect 9600 3200 9660 3210
rect 9670 3200 9910 3210
rect 9960 3200 9990 3210
rect 2130 3190 3160 3200
rect 5000 3190 5210 3200
rect 8430 3190 8760 3200
rect 8900 3190 9010 3200
rect 9600 3190 9640 3200
rect 9670 3190 9900 3200
rect 9940 3190 9990 3200
rect 2130 3180 3160 3190
rect 4860 3180 4870 3190
rect 5010 3180 5210 3190
rect 8430 3180 8990 3190
rect 9660 3180 9900 3190
rect 9950 3180 9990 3190
rect 2120 3170 3170 3180
rect 4850 3170 4860 3180
rect 5010 3170 5210 3180
rect 8420 3170 8960 3180
rect 9650 3170 9890 3180
rect 9960 3170 9990 3180
rect 2120 3160 3170 3170
rect 5010 3160 5210 3170
rect 8420 3160 8910 3170
rect 9640 3160 9880 3170
rect 9970 3160 9990 3170
rect 2120 3150 3170 3160
rect 5000 3150 5210 3160
rect 8410 3150 8870 3160
rect 9630 3150 9870 3160
rect 9980 3150 9990 3160
rect 2120 3140 3160 3150
rect 5000 3140 5200 3150
rect 8410 3140 8800 3150
rect 8810 3140 8820 3150
rect 9620 3140 9860 3150
rect 9990 3140 9990 3150
rect 2110 3130 3160 3140
rect 4420 3130 4430 3140
rect 5000 3130 5200 3140
rect 8400 3130 8790 3140
rect 9570 3130 9590 3140
rect 9610 3130 9850 3140
rect 2110 3120 3160 3130
rect 4420 3120 4450 3130
rect 4990 3120 5190 3130
rect 8390 3120 8770 3130
rect 8880 3120 8910 3130
rect 9570 3120 9840 3130
rect 2110 3110 3150 3120
rect 4420 3110 4460 3120
rect 4770 3110 4780 3120
rect 4980 3110 5190 3120
rect 8390 3110 8720 3120
rect 8780 3110 8800 3120
rect 8810 3110 8900 3120
rect 9000 3110 9020 3120
rect 9570 3110 9830 3120
rect 2110 3100 3160 3110
rect 4430 3100 4470 3110
rect 4630 3100 4640 3110
rect 4990 3100 5180 3110
rect 8390 3100 8430 3110
rect 8450 3100 8870 3110
rect 8980 3100 9010 3110
rect 9540 3100 9820 3110
rect 9890 3100 9930 3110
rect 2110 3090 3160 3100
rect 3910 3090 3930 3100
rect 4430 3090 4480 3100
rect 4990 3090 5180 3100
rect 8390 3090 8410 3100
rect 8450 3090 8860 3100
rect 8960 3090 9010 3100
rect 9530 3090 9810 3100
rect 9900 3090 9930 3100
rect 2110 3080 3150 3090
rect 3910 3080 3950 3090
rect 4400 3080 4410 3090
rect 4460 3080 4470 3090
rect 4980 3080 5170 3090
rect 8380 3080 8400 3090
rect 8450 3080 8840 3090
rect 8950 3080 9000 3090
rect 9530 3080 9800 3090
rect 9900 3080 9930 3090
rect 2110 3070 3150 3080
rect 3910 3070 3990 3080
rect 4980 3070 5160 3080
rect 8380 3070 8390 3080
rect 8450 3070 8830 3080
rect 8920 3070 8970 3080
rect 9520 3070 9790 3080
rect 9900 3070 9960 3080
rect 2110 3060 3140 3070
rect 3910 3060 4010 3070
rect 4990 3060 5160 3070
rect 8370 3060 8390 3070
rect 8450 3060 8790 3070
rect 8910 3060 8950 3070
rect 9520 3060 9790 3070
rect 9900 3060 9980 3070
rect 2110 3050 3140 3060
rect 3910 3050 4020 3060
rect 5000 3050 5150 3060
rect 8370 3050 8390 3060
rect 8410 3050 8430 3060
rect 8450 3050 8760 3060
rect 8870 3050 8920 3060
rect 9530 3050 9780 3060
rect 9910 3050 9990 3060
rect 2100 3040 3130 3050
rect 3910 3040 4030 3050
rect 4360 3040 4400 3050
rect 5000 3040 5130 3050
rect 8360 3040 8430 3050
rect 8440 3040 8720 3050
rect 8730 3040 8750 3050
rect 8840 3040 8900 3050
rect 9510 3040 9770 3050
rect 9910 3040 9990 3050
rect 2100 3030 3130 3040
rect 3920 3030 4030 3040
rect 4360 3030 4400 3040
rect 5010 3030 5120 3040
rect 8360 3030 8430 3040
rect 8450 3030 8640 3040
rect 8650 3030 8660 3040
rect 9510 3030 9760 3040
rect 9910 3030 9990 3040
rect 2100 3020 3130 3030
rect 3930 3020 4040 3030
rect 4370 3020 4410 3030
rect 5030 3020 5080 3030
rect 5090 3020 5110 3030
rect 8350 3020 8400 3030
rect 8450 3020 8630 3030
rect 9500 3020 9750 3030
rect 9920 3020 9990 3030
rect 2090 3010 3130 3020
rect 3920 3010 4040 3020
rect 4380 3010 4420 3020
rect 5100 3010 5120 3020
rect 8350 3010 8400 3020
rect 8450 3010 8590 3020
rect 8600 3010 8620 3020
rect 9490 3010 9750 3020
rect 9940 3010 9990 3020
rect 2090 3000 3130 3010
rect 3910 3000 4030 3010
rect 4390 3000 4430 3010
rect 8340 3000 8400 3010
rect 8450 3000 8600 3010
rect 9480 3000 9750 3010
rect 9960 3000 9990 3010
rect 2090 2990 3130 3000
rect 3900 2990 4020 3000
rect 4410 2990 4430 3000
rect 8340 2990 8400 3000
rect 8460 2990 8570 3000
rect 9470 2990 9770 3000
rect 9960 2990 9990 3000
rect 2080 2980 3130 2990
rect 3900 2980 4010 2990
rect 8330 2980 8400 2990
rect 8450 2980 8560 2990
rect 9470 2980 9790 2990
rect 9970 2980 9990 2990
rect 2080 2970 3120 2980
rect 3900 2970 4000 2980
rect 4080 2970 4110 2980
rect 8320 2970 8400 2980
rect 8450 2970 8550 2980
rect 9460 2970 9800 2980
rect 9870 2970 9890 2980
rect 9960 2970 9990 2980
rect 2080 2960 3120 2970
rect 3900 2960 3990 2970
rect 4000 2960 4010 2970
rect 4050 2960 4120 2970
rect 8320 2960 8410 2970
rect 8450 2960 8550 2970
rect 9460 2960 9810 2970
rect 9820 2960 9890 2970
rect 9950 2960 9990 2970
rect 2080 2950 3120 2960
rect 3900 2950 3980 2960
rect 4060 2950 4140 2960
rect 4150 2950 4160 2960
rect 8310 2950 8420 2960
rect 8450 2950 8550 2960
rect 9450 2950 9690 2960
rect 9720 2950 9910 2960
rect 9950 2950 9990 2960
rect 2090 2940 3120 2950
rect 3900 2940 3980 2950
rect 4060 2940 4150 2950
rect 4160 2940 4170 2950
rect 8310 2940 8550 2950
rect 9440 2940 9680 2950
rect 9740 2940 9920 2950
rect 9960 2940 9990 2950
rect 2080 2930 3110 2940
rect 3900 2930 3970 2940
rect 4050 2930 4080 2940
rect 4090 2930 4190 2940
rect 8300 2930 8550 2940
rect 9440 2930 9680 2940
rect 9740 2930 9930 2940
rect 9960 2930 9990 2940
rect 2080 2920 3110 2930
rect 4040 2920 4100 2930
rect 4110 2920 4200 2930
rect 8290 2920 8540 2930
rect 9430 2920 9670 2930
rect 9740 2920 9990 2930
rect 2080 2910 3110 2920
rect 4020 2910 4210 2920
rect 8290 2910 8500 2920
rect 9420 2910 9660 2920
rect 9730 2910 9990 2920
rect 2080 2900 3100 2910
rect 4020 2900 4220 2910
rect 8280 2900 8500 2910
rect 9420 2900 9650 2910
rect 9730 2900 9900 2910
rect 9970 2900 9990 2910
rect 2070 2890 3100 2900
rect 4010 2890 4230 2900
rect 8280 2890 8500 2900
rect 9410 2890 9640 2900
rect 9730 2890 9900 2900
rect 9980 2890 9990 2900
rect 2070 2880 3100 2890
rect 4010 2880 4240 2890
rect 8270 2880 8500 2890
rect 9400 2880 9650 2890
rect 9750 2880 9920 2890
rect 2070 2870 3100 2880
rect 4000 2870 4240 2880
rect 8260 2870 8500 2880
rect 9380 2870 9660 2880
rect 9740 2870 9920 2880
rect 2060 2860 3110 2870
rect 3990 2860 4240 2870
rect 7430 2860 7480 2870
rect 8250 2860 8500 2870
rect 9370 2860 9680 2870
rect 9740 2860 9930 2870
rect 2060 2850 3110 2860
rect 3990 2850 4250 2860
rect 7280 2850 7340 2860
rect 7390 2850 7510 2860
rect 8250 2850 8500 2860
rect 9370 2850 9690 2860
rect 9740 2850 9930 2860
rect 2050 2840 3110 2850
rect 3990 2840 4250 2850
rect 7250 2840 7520 2850
rect 8240 2840 8510 2850
rect 9370 2840 9710 2850
rect 9740 2840 9940 2850
rect 2050 2830 3090 2840
rect 3100 2830 3110 2840
rect 3990 2830 4080 2840
rect 4100 2830 4150 2840
rect 4160 2830 4250 2840
rect 7230 2830 7530 2840
rect 8230 2830 8520 2840
rect 9400 2830 9650 2840
rect 9670 2830 9720 2840
rect 9750 2830 9940 2840
rect 9950 2830 9990 2840
rect 2040 2820 3050 2830
rect 3990 2820 4070 2830
rect 4090 2820 4250 2830
rect 7220 2820 7540 2830
rect 8220 2820 8530 2830
rect 9420 2820 9600 2830
rect 9610 2820 9630 2830
rect 9680 2820 9730 2830
rect 9770 2820 9970 2830
rect 2050 2810 2900 2820
rect 2920 2810 3030 2820
rect 4010 2810 4070 2820
rect 4090 2810 4260 2820
rect 7200 2810 7550 2820
rect 8220 2810 8510 2820
rect 8520 2810 8530 2820
rect 9430 2810 9560 2820
rect 9660 2810 9670 2820
rect 9690 2810 9730 2820
rect 9780 2810 9920 2820
rect 9930 2810 9980 2820
rect 2060 2800 2250 2810
rect 2270 2800 2290 2810
rect 2390 2800 2840 2810
rect 2850 2800 2860 2810
rect 2970 2800 2990 2810
rect 3000 2800 3010 2810
rect 3990 2800 4260 2810
rect 7180 2800 7550 2810
rect 8210 2800 8500 2810
rect 9360 2800 9380 2810
rect 9450 2800 9550 2810
rect 9600 2800 9620 2810
rect 9670 2800 9760 2810
rect 9780 2800 9920 2810
rect 9940 2800 9990 2810
rect 2080 2790 2220 2800
rect 2410 2790 2810 2800
rect 3980 2790 4170 2800
rect 4180 2790 4260 2800
rect 7170 2790 7560 2800
rect 8200 2790 8500 2800
rect 9350 2790 9400 2800
rect 9470 2790 9580 2800
rect 9670 2790 9920 2800
rect 9990 2790 9990 2800
rect 2080 2780 2220 2790
rect 2430 2780 2800 2790
rect 3960 2780 4260 2790
rect 7150 2780 7590 2790
rect 8190 2780 8500 2790
rect 9340 2780 9380 2790
rect 9490 2780 9590 2790
rect 9620 2780 9630 2790
rect 9680 2780 9920 2790
rect 9990 2780 9990 2790
rect 2080 2770 2210 2780
rect 2430 2770 2790 2780
rect 3950 2770 4260 2780
rect 7140 2770 7600 2780
rect 8180 2770 8510 2780
rect 9340 2770 9390 2780
rect 9510 2770 9630 2780
rect 9690 2770 9920 2780
rect 9990 2770 9990 2780
rect 2090 2760 2200 2770
rect 2440 2760 2780 2770
rect 3950 2760 4150 2770
rect 4180 2760 4260 2770
rect 7120 2760 7610 2770
rect 8180 2760 8530 2770
rect 9330 2760 9400 2770
rect 9530 2760 9630 2770
rect 9690 2760 9710 2770
rect 9730 2760 9910 2770
rect 2080 2750 2180 2760
rect 2450 2750 2780 2760
rect 2990 2750 3030 2760
rect 3040 2750 3100 2760
rect 3950 2750 4170 2760
rect 4200 2750 4270 2760
rect 7100 2750 7620 2760
rect 8160 2750 8570 2760
rect 9320 2750 9400 2760
rect 9460 2750 9490 2760
rect 9550 2750 9630 2760
rect 9730 2750 9740 2760
rect 9750 2750 9900 2760
rect 2070 2740 2220 2750
rect 2460 2740 2770 2750
rect 2980 2740 3100 2750
rect 3950 2740 4170 2750
rect 4220 2740 4270 2750
rect 7080 2740 7630 2750
rect 8160 2740 8580 2750
rect 9320 2740 9400 2750
rect 9440 2740 9500 2750
rect 9570 2740 9620 2750
rect 9750 2740 9890 2750
rect 2080 2730 2260 2740
rect 2460 2730 2770 2740
rect 2950 2730 3100 2740
rect 3940 2730 4220 2740
rect 4250 2730 4270 2740
rect 7060 2730 7640 2740
rect 8150 2730 8570 2740
rect 9310 2730 9380 2740
rect 9430 2730 9530 2740
rect 9600 2730 9630 2740
rect 9710 2730 9730 2740
rect 9740 2730 9890 2740
rect 2080 2720 2270 2730
rect 2470 2720 2760 2730
rect 2940 2720 3110 2730
rect 3940 2720 4210 2730
rect 4250 2720 4270 2730
rect 7040 2720 7650 2730
rect 8140 2720 8580 2730
rect 9310 2720 9380 2730
rect 9420 2720 9550 2730
rect 9620 2720 9640 2730
rect 9700 2720 9730 2730
rect 9740 2720 9890 2730
rect 2080 2710 2280 2720
rect 2470 2710 2760 2720
rect 2950 2710 3110 2720
rect 3930 2710 4220 2720
rect 4250 2710 4270 2720
rect 7020 2710 7650 2720
rect 8130 2710 8550 2720
rect 9300 2710 9350 2720
rect 9410 2710 9570 2720
rect 9640 2710 9660 2720
rect 9690 2710 9710 2720
rect 9740 2710 9810 2720
rect 9820 2710 9890 2720
rect 2050 2700 2270 2710
rect 2470 2700 2750 2710
rect 2950 2700 3110 2710
rect 3930 2700 4230 2710
rect 4240 2700 4270 2710
rect 7000 2700 7660 2710
rect 8120 2700 8560 2710
rect 9290 2700 9370 2710
rect 9390 2700 9590 2710
rect 9660 2700 9710 2710
rect 9730 2700 9900 2710
rect 2050 2690 2220 2700
rect 2470 2690 2750 2700
rect 2950 2690 3110 2700
rect 3930 2690 4270 2700
rect 6990 2690 7160 2700
rect 7170 2690 7670 2700
rect 8120 2690 8540 2700
rect 8550 2690 8560 2700
rect 9300 2690 9610 2700
rect 9680 2690 9910 2700
rect 2040 2680 2200 2690
rect 2480 2680 2740 2690
rect 3060 2680 3090 2690
rect 3930 2680 4240 2690
rect 4250 2680 4270 2690
rect 6970 2680 7160 2690
rect 7170 2680 7670 2690
rect 8110 2680 8510 2690
rect 8530 2680 8550 2690
rect 8570 2680 8580 2690
rect 9280 2680 9630 2690
rect 9700 2680 9940 2690
rect 2030 2670 2160 2680
rect 2480 2670 2740 2680
rect 3920 2670 4220 2680
rect 4250 2670 4270 2680
rect 6960 2670 7160 2680
rect 7170 2670 7680 2680
rect 8100 2670 8540 2680
rect 8550 2670 8560 2680
rect 8570 2670 8580 2680
rect 9260 2670 9650 2680
rect 9720 2670 9950 2680
rect 2030 2660 2140 2670
rect 2480 2660 2740 2670
rect 3910 2660 4200 2670
rect 4250 2660 4270 2670
rect 6940 2660 7160 2670
rect 7180 2660 7690 2670
rect 8090 2660 8520 2670
rect 8560 2660 8590 2670
rect 9250 2660 9670 2670
rect 9740 2660 9960 2670
rect 2020 2650 2090 2660
rect 2480 2650 2740 2660
rect 3920 2650 4190 2660
rect 4240 2650 4260 2660
rect 6930 2650 7140 2660
rect 7150 2650 7170 2660
rect 7190 2650 7690 2660
rect 8080 2650 8500 2660
rect 8550 2650 8590 2660
rect 9230 2650 9690 2660
rect 9760 2650 9970 2660
rect 2030 2640 2070 2650
rect 2480 2640 2730 2650
rect 2980 2640 3020 2650
rect 3930 2640 4180 2650
rect 4240 2640 4260 2650
rect 6920 2640 7130 2650
rect 7190 2640 7700 2650
rect 8070 2640 8500 2650
rect 8520 2640 8530 2650
rect 8550 2640 8600 2650
rect 9220 2640 9710 2650
rect 9780 2640 9880 2650
rect 9890 2640 9930 2650
rect 9940 2640 9950 2650
rect 2480 2630 2730 2640
rect 2970 2630 3050 2640
rect 3930 2630 4190 2640
rect 4240 2630 4260 2640
rect 6910 2630 7130 2640
rect 7220 2630 7240 2640
rect 7250 2630 7700 2640
rect 8060 2630 8430 2640
rect 8470 2630 8510 2640
rect 8520 2630 8540 2640
rect 8550 2630 8600 2640
rect 9210 2630 9730 2640
rect 9800 2630 9840 2640
rect 2200 2620 2250 2630
rect 2490 2620 2730 2630
rect 2940 2620 2950 2630
rect 3020 2620 3030 2630
rect 3940 2620 4190 2630
rect 4230 2620 4260 2630
rect 6900 2620 7140 2630
rect 7220 2620 7240 2630
rect 7260 2620 7710 2630
rect 8050 2620 8410 2630
rect 8480 2620 8520 2630
rect 8560 2620 8590 2630
rect 8610 2620 8620 2630
rect 9200 2620 9750 2630
rect 9820 2620 9850 2630
rect 2480 2610 2730 2620
rect 3950 2610 4200 2620
rect 4230 2610 4260 2620
rect 6890 2610 7130 2620
rect 7230 2610 7240 2620
rect 7260 2610 7270 2620
rect 7280 2610 7720 2620
rect 8040 2610 8400 2620
rect 8490 2610 8530 2620
rect 8570 2610 8580 2620
rect 9200 2610 9770 2620
rect 9830 2610 9860 2620
rect 2480 2600 2730 2610
rect 3950 2600 4200 2610
rect 4230 2600 4260 2610
rect 6880 2600 7130 2610
rect 7140 2600 7150 2610
rect 7280 2600 7720 2610
rect 8030 2600 8400 2610
rect 8490 2600 8550 2610
rect 9200 2600 9790 2610
rect 2470 2590 2730 2600
rect 3950 2590 4080 2600
rect 4100 2590 4200 2600
rect 4230 2590 4250 2600
rect 6870 2590 7130 2600
rect 7290 2590 7730 2600
rect 8020 2590 8400 2600
rect 8500 2590 8560 2600
rect 9200 2590 9800 2600
rect 9880 2590 9900 2600
rect 2460 2580 2730 2590
rect 3960 2580 4060 2590
rect 4080 2580 4190 2590
rect 4240 2580 4250 2590
rect 6860 2580 7100 2590
rect 7150 2580 7160 2590
rect 7290 2580 7740 2590
rect 8010 2580 8400 2590
rect 8490 2580 8500 2590
rect 8510 2580 8520 2590
rect 8540 2580 8580 2590
rect 9190 2580 9830 2590
rect 9900 2580 9920 2590
rect 2450 2570 2730 2580
rect 3920 2570 4040 2580
rect 4070 2570 4090 2580
rect 4110 2570 4180 2580
rect 6850 2570 7100 2580
rect 7160 2570 7170 2580
rect 7300 2570 7750 2580
rect 8000 2570 8400 2580
rect 9190 2570 9320 2580
rect 9330 2570 9490 2580
rect 9530 2570 9850 2580
rect 9920 2570 9940 2580
rect 2430 2560 2730 2570
rect 3950 2560 4040 2570
rect 4080 2560 4090 2570
rect 4110 2560 4170 2570
rect 6850 2560 7110 2570
rect 7170 2560 7180 2570
rect 7310 2560 7760 2570
rect 7990 2560 8400 2570
rect 8490 2560 8500 2570
rect 8580 2560 8630 2570
rect 9190 2560 9310 2570
rect 9330 2560 9390 2570
rect 9420 2560 9470 2570
rect 9550 2560 9870 2570
rect 2430 2550 2740 2560
rect 2800 2550 2820 2560
rect 4020 2550 4030 2560
rect 4100 2550 4150 2560
rect 6840 2550 7120 2560
rect 7180 2550 7190 2560
rect 7320 2550 7770 2560
rect 7980 2550 8400 2560
rect 8490 2550 8500 2560
rect 8580 2550 8640 2560
rect 9190 2550 9340 2560
rect 9360 2550 9380 2560
rect 9480 2550 9490 2560
rect 9570 2550 9890 2560
rect 9970 2550 9980 2560
rect 2430 2540 2740 2550
rect 2790 2540 2820 2550
rect 3960 2540 3990 2550
rect 4010 2540 4030 2550
rect 4060 2540 4070 2550
rect 4110 2540 4120 2550
rect 6830 2540 7130 2550
rect 7190 2540 7210 2550
rect 7330 2540 7770 2550
rect 7960 2540 8390 2550
rect 8580 2540 8590 2550
rect 8660 2540 8670 2550
rect 9180 2540 9340 2550
rect 9360 2540 9380 2550
rect 9480 2540 9500 2550
rect 9590 2540 9910 2550
rect 9980 2540 9990 2550
rect 2420 2530 2750 2540
rect 2760 2530 2820 2540
rect 2970 2530 3010 2540
rect 3970 2530 4050 2540
rect 4060 2530 4080 2540
rect 6820 2530 6830 2540
rect 6840 2530 7160 2540
rect 7210 2530 7230 2540
rect 7340 2530 7780 2540
rect 7950 2530 8390 2540
rect 8670 2530 8680 2540
rect 9180 2530 9340 2540
rect 9610 2530 9930 2540
rect 2410 2520 2840 2530
rect 2920 2520 3100 2530
rect 4070 2520 4080 2530
rect 6810 2520 6830 2530
rect 6850 2520 7180 2530
rect 7340 2520 7780 2530
rect 7940 2520 8390 2530
rect 9170 2520 9330 2530
rect 9630 2520 9950 2530
rect 2390 2510 2870 2520
rect 2900 2510 3120 2520
rect 6800 2510 6830 2520
rect 6850 2510 7190 2520
rect 7340 2510 7790 2520
rect 7920 2510 8390 2520
rect 8690 2510 8700 2520
rect 9170 2510 9300 2520
rect 9420 2510 9440 2520
rect 9650 2510 9970 2520
rect 2020 2500 2040 2510
rect 2120 2500 2200 2510
rect 2370 2500 3120 2510
rect 6790 2500 6820 2510
rect 6830 2500 6840 2510
rect 6860 2500 7210 2510
rect 7350 2500 7800 2510
rect 7910 2500 8390 2510
rect 9170 2500 9270 2510
rect 9420 2500 9430 2510
rect 9590 2500 9600 2510
rect 9670 2500 9990 2510
rect 2000 2490 2060 2500
rect 2120 2490 2230 2500
rect 2360 2490 3100 2500
rect 3190 2490 3200 2500
rect 6790 2490 6810 2500
rect 6860 2490 7220 2500
rect 7360 2490 7800 2500
rect 7890 2490 8390 2500
rect 8750 2490 8760 2500
rect 9160 2490 9260 2500
rect 9590 2490 9600 2500
rect 9690 2490 9990 2500
rect 1980 2480 2180 2490
rect 2190 2480 2200 2490
rect 2310 2480 3070 2490
rect 3150 2480 3200 2490
rect 6780 2480 6790 2490
rect 6870 2480 7230 2490
rect 7370 2480 7810 2490
rect 7870 2480 8390 2490
rect 8780 2480 8790 2490
rect 9160 2480 9250 2490
rect 9710 2480 9990 2490
rect 1970 2470 2190 2480
rect 2250 2470 2300 2480
rect 2310 2470 2920 2480
rect 3130 2470 3200 2480
rect 6870 2470 7240 2480
rect 7380 2470 7810 2480
rect 7850 2470 8390 2480
rect 8770 2470 8800 2480
rect 9160 2470 9240 2480
rect 9730 2470 9990 2480
rect 1960 2460 2280 2470
rect 2330 2460 2930 2470
rect 3110 2460 3190 2470
rect 6870 2460 7250 2470
rect 7430 2460 7820 2470
rect 7830 2460 8390 2470
rect 9160 2460 9240 2470
rect 9740 2460 9990 2470
rect 1950 2450 2060 2460
rect 2140 2450 2230 2460
rect 2320 2450 2960 2460
rect 3070 2450 3200 2460
rect 6880 2450 7260 2460
rect 7440 2450 8390 2460
rect 9150 2450 9230 2460
rect 9740 2450 9990 2460
rect 1940 2440 2060 2450
rect 2310 2440 3200 2450
rect 6890 2440 7280 2450
rect 7440 2440 8390 2450
rect 9150 2440 9230 2450
rect 9270 2440 9290 2450
rect 9790 2440 9990 2450
rect 1960 2430 2100 2440
rect 2290 2430 3210 2440
rect 6910 2430 7290 2440
rect 7450 2430 8390 2440
rect 9160 2430 9220 2440
rect 9270 2430 9290 2440
rect 9680 2430 9700 2440
rect 9790 2430 9990 2440
rect 1960 2420 2130 2430
rect 2270 2420 3210 2430
rect 6920 2420 7310 2430
rect 7450 2420 8400 2430
rect 9160 2420 9210 2430
rect 9280 2420 9300 2430
rect 9650 2420 9660 2430
rect 9680 2420 9710 2430
rect 9800 2420 9990 2430
rect 1960 2410 2150 2420
rect 2220 2410 3210 2420
rect 6930 2410 7330 2420
rect 7460 2410 8390 2420
rect 9170 2410 9200 2420
rect 9210 2410 9220 2420
rect 9270 2410 9300 2420
rect 9360 2410 9370 2420
rect 9380 2410 9390 2420
rect 9490 2410 9560 2420
rect 9650 2410 9670 2420
rect 9810 2410 9990 2420
rect 1970 2400 3220 2410
rect 6970 2400 7350 2410
rect 7470 2400 8390 2410
rect 9180 2400 9240 2410
rect 9260 2400 9290 2410
rect 9340 2400 9390 2410
rect 9420 2400 9440 2410
rect 9490 2400 9570 2410
rect 9650 2400 9680 2410
rect 9820 2400 9830 2410
rect 9850 2400 9990 2410
rect 1970 2390 3220 2400
rect 6990 2390 7370 2400
rect 7480 2390 8390 2400
rect 9190 2390 9280 2400
rect 9330 2390 9400 2400
rect 9480 2390 9520 2400
rect 9550 2390 9580 2400
rect 9650 2390 9670 2400
rect 9850 2390 9990 2400
rect 1970 2380 3220 2390
rect 7010 2380 7020 2390
rect 7040 2380 7380 2390
rect 7490 2380 8390 2390
rect 9200 2380 9260 2390
rect 9320 2380 9390 2390
rect 9470 2380 9520 2390
rect 9560 2380 9570 2390
rect 9850 2380 9990 2390
rect 1970 2370 3220 2380
rect 7090 2370 7390 2380
rect 7500 2370 8390 2380
rect 8700 2370 8710 2380
rect 8740 2370 8760 2380
rect 8860 2370 8900 2380
rect 9210 2370 9260 2380
rect 9320 2370 9380 2380
rect 9470 2370 9530 2380
rect 9830 2370 9990 2380
rect 1950 2360 3230 2370
rect 7090 2360 7410 2370
rect 7510 2360 8390 2370
rect 8670 2360 8760 2370
rect 8850 2360 8860 2370
rect 8870 2360 8890 2370
rect 9210 2360 9250 2370
rect 9280 2360 9300 2370
rect 9340 2360 9370 2370
rect 9480 2360 9630 2370
rect 9650 2360 9670 2370
rect 9840 2360 9990 2370
rect 1960 2350 3230 2360
rect 7150 2350 7420 2360
rect 7510 2350 8390 2360
rect 8650 2350 8760 2360
rect 8870 2350 8890 2360
rect 9220 2350 9240 2360
rect 9270 2350 9300 2360
rect 9500 2350 9550 2360
rect 9590 2350 9600 2360
rect 9610 2350 9630 2360
rect 9640 2350 9670 2360
rect 9860 2350 9990 2360
rect 1950 2340 3230 2350
rect 7170 2340 7440 2350
rect 7520 2340 8390 2350
rect 8660 2340 8750 2350
rect 9140 2340 9150 2350
rect 9220 2340 9230 2350
rect 9270 2340 9310 2350
rect 9500 2340 9540 2350
rect 9860 2340 9920 2350
rect 9930 2340 9990 2350
rect 1950 2330 3230 2340
rect 7180 2330 7460 2340
rect 7530 2330 8390 2340
rect 8660 2330 8750 2340
rect 8850 2330 8860 2340
rect 8930 2330 8980 2340
rect 9140 2330 9150 2340
rect 9220 2330 9230 2340
rect 9290 2330 9300 2340
rect 9420 2330 9430 2340
rect 9500 2330 9540 2340
rect 9850 2330 9910 2340
rect 9930 2330 9990 2340
rect 1940 2320 3230 2330
rect 7210 2320 7470 2330
rect 7550 2320 8370 2330
rect 8660 2320 8750 2330
rect 8840 2320 8880 2330
rect 8920 2320 8980 2330
rect 9140 2320 9150 2330
rect 9220 2320 9230 2330
rect 9410 2320 9430 2330
rect 9510 2320 9530 2330
rect 9840 2320 9990 2330
rect 1930 2310 3230 2320
rect 7230 2310 7480 2320
rect 7590 2310 8370 2320
rect 8660 2310 8740 2320
rect 8830 2310 8960 2320
rect 9130 2310 9150 2320
rect 9210 2310 9220 2320
rect 9420 2310 9430 2320
rect 9840 2310 9990 2320
rect 1930 2300 3240 2310
rect 7240 2300 7260 2310
rect 7270 2300 7490 2310
rect 7590 2300 8360 2310
rect 8660 2300 8720 2310
rect 8830 2300 8930 2310
rect 9140 2300 9150 2310
rect 9210 2300 9220 2310
rect 9840 2300 9990 2310
rect 1930 2290 3240 2300
rect 7270 2290 7330 2300
rect 7340 2290 7490 2300
rect 7620 2290 8360 2300
rect 8660 2290 8720 2300
rect 8860 2290 8900 2300
rect 9140 2290 9150 2300
rect 9490 2290 9520 2300
rect 9830 2290 9990 2300
rect 1930 2280 3250 2290
rect 7290 2280 7320 2290
rect 7340 2280 7360 2290
rect 7400 2280 7490 2290
rect 7620 2280 8360 2290
rect 8670 2280 8720 2290
rect 8860 2280 8870 2290
rect 9140 2280 9150 2290
rect 9500 2280 9570 2290
rect 9800 2280 9990 2290
rect 1930 2270 3250 2280
rect 7290 2270 7300 2280
rect 7420 2270 7480 2280
rect 7630 2270 8360 2280
rect 8680 2270 8690 2280
rect 9510 2270 9530 2280
rect 9540 2270 9560 2280
rect 9800 2270 9990 2280
rect 1930 2260 3250 2270
rect 7430 2260 7500 2270
rect 7630 2260 8360 2270
rect 9800 2260 9870 2270
rect 9880 2260 9990 2270
rect 1930 2250 3250 2260
rect 7440 2250 7500 2260
rect 7640 2250 8360 2260
rect 8890 2250 8910 2260
rect 9010 2250 9020 2260
rect 9800 2250 9990 2260
rect 1910 2240 2690 2250
rect 2720 2240 3250 2250
rect 7430 2240 7500 2250
rect 7650 2240 8360 2250
rect 8870 2240 9030 2250
rect 9800 2240 9990 2250
rect 1910 2230 2650 2240
rect 2730 2230 3250 2240
rect 6440 2230 6450 2240
rect 7400 2230 7420 2240
rect 7430 2230 7500 2240
rect 7660 2230 8360 2240
rect 8860 2230 9020 2240
rect 9250 2230 9270 2240
rect 9800 2230 9990 2240
rect 1910 2220 2490 2230
rect 2510 2220 2610 2230
rect 2740 2220 3250 2230
rect 7400 2220 7500 2230
rect 7680 2220 8360 2230
rect 8850 2220 8990 2230
rect 9250 2220 9300 2230
rect 9580 2220 9590 2230
rect 9820 2220 9990 2230
rect 1910 2210 2470 2220
rect 2750 2210 3250 2220
rect 6440 2210 6450 2220
rect 7400 2210 7490 2220
rect 7690 2210 8360 2220
rect 8870 2210 8970 2220
rect 9250 2210 9320 2220
rect 9580 2210 9590 2220
rect 9820 2210 9980 2220
rect 9990 2210 9990 2220
rect 1910 2200 2470 2210
rect 2770 2200 2820 2210
rect 2850 2200 3250 2210
rect 6440 2200 6460 2210
rect 7390 2200 7420 2210
rect 7430 2200 7480 2210
rect 7710 2200 8360 2210
rect 9250 2200 9350 2210
rect 9680 2200 9700 2210
rect 9810 2200 9960 2210
rect 1910 2190 2450 2200
rect 2860 2190 3240 2200
rect 6440 2190 6460 2200
rect 7400 2190 7410 2200
rect 7430 2190 7470 2200
rect 7730 2190 8360 2200
rect 9250 2190 9370 2200
rect 9820 2190 9950 2200
rect 1910 2180 2280 2190
rect 2310 2180 2420 2190
rect 2860 2180 3240 2190
rect 6440 2180 6460 2190
rect 7440 2180 7450 2190
rect 7740 2180 8360 2190
rect 9250 2180 9390 2190
rect 9820 2180 9950 2190
rect 9990 2180 9990 2190
rect 1910 2170 2260 2180
rect 2310 2170 2350 2180
rect 2860 2170 3240 2180
rect 6460 2170 6470 2180
rect 7750 2170 8360 2180
rect 9250 2170 9410 2180
rect 9810 2170 9960 2180
rect 9990 2170 9990 2180
rect 1910 2160 2250 2170
rect 2300 2160 2350 2170
rect 2860 2160 3230 2170
rect 6450 2160 6460 2170
rect 7780 2160 8370 2170
rect 9250 2160 9430 2170
rect 9800 2160 9980 2170
rect 9990 2160 9990 2170
rect 1920 2150 2240 2160
rect 2300 2150 2350 2160
rect 2840 2150 3230 2160
rect 6450 2150 6460 2160
rect 7840 2150 8370 2160
rect 9280 2150 9440 2160
rect 9560 2150 9570 2160
rect 9580 2150 9590 2160
rect 9790 2150 9950 2160
rect 9960 2150 9980 2160
rect 9990 2150 9990 2160
rect 1920 2140 2230 2150
rect 2290 2140 2360 2150
rect 2830 2140 3230 2150
rect 6440 2140 6460 2150
rect 7850 2140 8370 2150
rect 9300 2140 9460 2150
rect 9570 2140 9590 2150
rect 9790 2140 9940 2150
rect 9950 2140 9980 2150
rect 9990 2140 9990 2150
rect 1930 2130 2220 2140
rect 2290 2130 2360 2140
rect 2820 2130 3220 2140
rect 6440 2130 6450 2140
rect 7860 2130 8380 2140
rect 9320 2130 9480 2140
rect 9570 2130 9590 2140
rect 9780 2130 9910 2140
rect 9920 2130 9990 2140
rect 1930 2120 2220 2130
rect 2280 2120 2370 2130
rect 2800 2120 3220 2130
rect 6440 2120 6450 2130
rect 7870 2120 8380 2130
rect 9230 2120 9250 2130
rect 9330 2120 9500 2130
rect 9570 2120 9580 2130
rect 9670 2120 9690 2130
rect 9770 2120 9990 2130
rect 1940 2110 2210 2120
rect 2270 2110 2380 2120
rect 2490 2110 2520 2120
rect 2670 2110 2740 2120
rect 2770 2110 3220 2120
rect 6430 2110 6450 2120
rect 7880 2110 8390 2120
rect 9350 2110 9520 2120
rect 9570 2110 9650 2120
rect 9700 2110 9720 2120
rect 9760 2110 9990 2120
rect 1930 2100 2210 2110
rect 2260 2100 2400 2110
rect 2430 2100 2540 2110
rect 2640 2100 3220 2110
rect 6430 2100 6450 2110
rect 7880 2100 8390 2110
rect 9370 2100 9610 2110
rect 9700 2100 9990 2110
rect 1940 2090 2200 2100
rect 2260 2090 2550 2100
rect 2620 2090 3200 2100
rect 6430 2090 6450 2100
rect 7880 2090 8390 2100
rect 9380 2090 9530 2100
rect 9710 2090 9990 2100
rect 1940 2080 2180 2090
rect 2250 2080 3200 2090
rect 7900 2080 8390 2090
rect 9240 2080 9260 2090
rect 9360 2080 9450 2090
rect 9710 2080 9990 2090
rect 1940 2070 2180 2080
rect 2240 2070 3190 2080
rect 6430 2070 6440 2080
rect 7900 2070 8380 2080
rect 9230 2070 9260 2080
rect 9290 2070 9370 2080
rect 9700 2070 9990 2080
rect 1960 2060 2170 2070
rect 2230 2060 3180 2070
rect 8000 2060 8380 2070
rect 9220 2060 9270 2070
rect 9690 2060 9990 2070
rect 1960 2050 2160 2060
rect 2220 2050 3170 2060
rect 8010 2050 8380 2060
rect 9160 2050 9210 2060
rect 9540 2050 9550 2060
rect 9680 2050 9990 2060
rect 1980 2040 2150 2050
rect 2220 2040 3160 2050
rect 8010 2040 8380 2050
rect 9490 2040 9620 2050
rect 9650 2040 9990 2050
rect 1990 2030 2100 2040
rect 2210 2030 3150 2040
rect 8010 2030 8380 2040
rect 9480 2030 9990 2040
rect 2000 2020 2080 2030
rect 2200 2020 3130 2030
rect 8010 2020 8380 2030
rect 9350 2020 9360 2030
rect 9470 2020 9990 2030
rect 2010 2010 2040 2020
rect 2200 2010 3120 2020
rect 8000 2010 8380 2020
rect 9280 2010 9390 2020
rect 9430 2010 9990 2020
rect 2010 2000 2020 2010
rect 2200 2000 3120 2010
rect 7980 2000 8380 2010
rect 9090 2000 9110 2010
rect 9190 2000 9990 2010
rect 2190 1990 3110 2000
rect 7320 1990 7330 2000
rect 7980 1990 8380 2000
rect 9070 1990 9110 2000
rect 9140 1990 9680 2000
rect 9690 1990 9990 2000
rect 2180 1980 3110 1990
rect 7320 1980 7330 1990
rect 7990 1980 8380 1990
rect 9060 1980 9080 1990
rect 9100 1980 9110 1990
rect 9140 1980 9650 1990
rect 9680 1980 9990 1990
rect 2180 1970 3100 1980
rect 6410 1970 6420 1980
rect 7320 1970 7330 1980
rect 7980 1970 8380 1980
rect 9050 1970 9060 1980
rect 9130 1970 9990 1980
rect 2180 1960 3110 1970
rect 6410 1960 6430 1970
rect 7980 1960 8380 1970
rect 9130 1960 9670 1970
rect 9680 1960 9920 1970
rect 9960 1960 9990 1970
rect 2170 1950 3100 1960
rect 6410 1950 6430 1960
rect 7970 1950 8380 1960
rect 9130 1950 9670 1960
rect 9680 1950 9880 1960
rect 9960 1950 9990 1960
rect 2170 1940 3110 1950
rect 7960 1940 8380 1950
rect 9130 1940 9660 1950
rect 9690 1940 9850 1950
rect 9860 1940 9880 1950
rect 9910 1940 9940 1950
rect 9990 1940 9990 1950
rect 2170 1930 3030 1940
rect 3040 1930 3110 1940
rect 4800 1930 4830 1940
rect 7890 1930 8380 1940
rect 8830 1930 8900 1940
rect 9130 1930 9640 1940
rect 9690 1930 9850 1940
rect 9910 1930 9980 1940
rect 2160 1920 2650 1930
rect 2720 1920 3010 1930
rect 3030 1920 3110 1930
rect 4510 1920 4590 1930
rect 4610 1920 4630 1930
rect 4790 1920 4850 1930
rect 7900 1920 8380 1930
rect 8800 1920 8930 1930
rect 9130 1920 9600 1930
rect 9690 1920 9860 1930
rect 9920 1920 9960 1930
rect 9970 1920 9980 1930
rect 9990 1920 9990 1930
rect 2160 1910 2600 1920
rect 2760 1910 2850 1920
rect 2880 1910 2890 1920
rect 2900 1910 2990 1920
rect 3040 1910 3110 1920
rect 4490 1910 4530 1920
rect 4620 1910 4640 1920
rect 4780 1910 4800 1920
rect 4980 1910 5000 1920
rect 7910 1910 8370 1920
rect 8690 1910 8960 1920
rect 9120 1910 9600 1920
rect 9710 1910 9880 1920
rect 9910 1910 9960 1920
rect 9980 1910 9990 1920
rect 2160 1900 2450 1910
rect 2930 1900 2980 1910
rect 3030 1900 3110 1910
rect 4480 1900 4500 1910
rect 4630 1900 4640 1910
rect 4780 1900 4800 1910
rect 4980 1900 5000 1910
rect 5050 1900 5100 1910
rect 7910 1900 8370 1910
rect 8680 1900 8960 1910
rect 9120 1900 9590 1910
rect 9640 1900 9670 1910
rect 9740 1900 9950 1910
rect 9980 1900 9990 1910
rect 2160 1890 2430 1900
rect 2950 1890 2970 1900
rect 3020 1890 3110 1900
rect 4410 1890 4420 1900
rect 4480 1890 4500 1900
rect 4780 1890 4790 1900
rect 4850 1890 4870 1900
rect 4980 1890 5000 1900
rect 5070 1890 5130 1900
rect 7910 1890 8370 1900
rect 8660 1890 8980 1900
rect 9120 1890 9580 1900
rect 9620 1890 9670 1900
rect 9760 1890 9930 1900
rect 9980 1890 9990 1900
rect 2160 1880 2410 1890
rect 2950 1880 2970 1890
rect 3020 1880 3110 1890
rect 4350 1880 4360 1890
rect 4410 1880 4420 1890
rect 4480 1880 4500 1890
rect 4560 1880 4570 1890
rect 4640 1880 4650 1890
rect 4770 1880 4790 1890
rect 4850 1880 4870 1890
rect 4990 1880 5010 1890
rect 5110 1880 5140 1890
rect 7920 1880 8370 1890
rect 8640 1880 8990 1890
rect 9120 1880 9240 1890
rect 9250 1880 9580 1890
rect 9610 1880 9680 1890
rect 9770 1880 9990 1890
rect 2160 1870 2390 1880
rect 2950 1870 2970 1880
rect 3010 1870 3110 1880
rect 4410 1870 4420 1880
rect 4480 1870 4500 1880
rect 4550 1870 4560 1880
rect 4640 1870 4650 1880
rect 4770 1870 4790 1880
rect 4850 1870 4870 1880
rect 5000 1870 5030 1880
rect 5120 1870 5140 1880
rect 7920 1870 8370 1880
rect 8630 1870 8990 1880
rect 9120 1870 9140 1880
rect 9210 1870 9240 1880
rect 9260 1870 9530 1880
rect 9540 1870 9570 1880
rect 9600 1870 9690 1880
rect 9770 1870 9990 1880
rect 2170 1860 2370 1870
rect 2950 1860 3120 1870
rect 4390 1860 4400 1870
rect 4480 1860 4490 1870
rect 4540 1860 4550 1870
rect 4590 1860 4600 1870
rect 4640 1860 4650 1870
rect 4770 1860 4780 1870
rect 4860 1860 4870 1870
rect 5020 1860 5030 1870
rect 5120 1860 5140 1870
rect 5240 1860 5260 1870
rect 7930 1860 8370 1870
rect 8630 1860 8990 1870
rect 9210 1860 9250 1870
rect 9380 1860 9420 1870
rect 9430 1860 9520 1870
rect 9530 1860 9690 1870
rect 9770 1860 9980 1870
rect 2170 1850 2230 1860
rect 2280 1850 2290 1860
rect 2330 1850 2340 1860
rect 2950 1850 3120 1860
rect 4370 1850 4380 1860
rect 4480 1850 4490 1860
rect 4540 1850 4550 1860
rect 4590 1850 4600 1860
rect 4640 1850 4650 1860
rect 4760 1850 4780 1860
rect 4860 1850 4870 1860
rect 5020 1850 5040 1860
rect 5090 1850 5130 1860
rect 5190 1850 5220 1860
rect 5240 1850 5290 1860
rect 7920 1850 8370 1860
rect 8630 1850 8980 1860
rect 9230 1850 9250 1860
rect 9290 1850 9310 1860
rect 9340 1850 9360 1860
rect 9370 1850 9690 1860
rect 9780 1850 9970 1860
rect 2170 1840 2210 1850
rect 2960 1840 3120 1850
rect 4480 1840 4500 1850
rect 4540 1840 4550 1850
rect 4590 1840 4600 1850
rect 4640 1840 4650 1850
rect 4760 1840 4770 1850
rect 4860 1840 4870 1850
rect 5020 1840 5030 1850
rect 5180 1840 5210 1850
rect 5270 1840 5300 1850
rect 7920 1840 8360 1850
rect 8630 1840 8980 1850
rect 9240 1840 9310 1850
rect 9340 1840 9690 1850
rect 9780 1840 9970 1850
rect 2180 1830 2200 1840
rect 2950 1830 3130 1840
rect 4480 1830 4500 1840
rect 4540 1830 4550 1840
rect 4590 1830 4600 1840
rect 4640 1830 4650 1840
rect 4750 1830 4770 1840
rect 4860 1830 4870 1840
rect 5010 1830 5030 1840
rect 5070 1830 5080 1840
rect 5170 1830 5190 1840
rect 5290 1830 5310 1840
rect 7930 1830 8360 1840
rect 8630 1830 8960 1840
rect 9230 1830 9300 1840
rect 9330 1830 9370 1840
rect 9420 1830 9690 1840
rect 9780 1830 9960 1840
rect 2160 1820 2190 1830
rect 2960 1820 3130 1830
rect 4480 1820 4490 1830
rect 4540 1820 4550 1830
rect 4580 1820 4600 1830
rect 4640 1820 4650 1830
rect 4750 1820 4770 1830
rect 4860 1820 4870 1830
rect 5010 1820 5030 1830
rect 5060 1820 5080 1830
rect 5170 1820 5190 1830
rect 5300 1820 5320 1830
rect 7940 1820 8360 1830
rect 8630 1820 8950 1830
rect 9210 1820 9280 1830
rect 9330 1820 9380 1830
rect 9430 1820 9690 1830
rect 9770 1820 9960 1830
rect 2150 1810 2190 1820
rect 2950 1810 3130 1820
rect 4480 1810 4500 1820
rect 4570 1810 4590 1820
rect 4630 1810 4640 1820
rect 4750 1810 4760 1820
rect 4800 1810 4820 1820
rect 4860 1810 4870 1820
rect 5010 1810 5030 1820
rect 5060 1810 5080 1820
rect 5160 1810 5180 1820
rect 5320 1810 5330 1820
rect 7950 1810 8360 1820
rect 8630 1810 8930 1820
rect 9200 1810 9250 1820
rect 9330 1810 9380 1820
rect 9440 1810 9700 1820
rect 9770 1810 9950 1820
rect 9990 1810 9990 1820
rect 2140 1800 2190 1810
rect 2930 1800 3150 1810
rect 4280 1800 4290 1810
rect 4480 1800 4490 1810
rect 4560 1800 4580 1810
rect 4630 1800 4640 1810
rect 4750 1800 4760 1810
rect 4790 1800 4830 1810
rect 4860 1800 4880 1810
rect 5000 1800 5020 1810
rect 5060 1800 5070 1810
rect 5160 1800 5170 1810
rect 5260 1800 5270 1810
rect 5320 1800 5330 1810
rect 7940 1800 8360 1810
rect 8620 1800 8930 1810
rect 9210 1800 9250 1810
rect 9290 1800 9300 1810
rect 9310 1800 9320 1810
rect 9380 1800 9400 1810
rect 9460 1800 9700 1810
rect 9780 1800 9950 1810
rect 9980 1800 9990 1810
rect 2080 1790 2100 1800
rect 2110 1790 2200 1800
rect 2820 1790 3150 1800
rect 4120 1790 4180 1800
rect 4480 1790 4490 1800
rect 4620 1790 4630 1800
rect 4740 1790 4760 1800
rect 4790 1790 4800 1800
rect 4820 1790 4830 1800
rect 4860 1790 4880 1800
rect 5000 1790 5020 1800
rect 5050 1790 5070 1800
rect 5150 1790 5170 1800
rect 5260 1790 5280 1800
rect 5320 1790 5340 1800
rect 7940 1790 8360 1800
rect 8620 1790 8930 1800
rect 9230 1790 9240 1800
rect 9270 1790 9280 1800
rect 9290 1790 9320 1800
rect 9340 1790 9420 1800
rect 9470 1790 9600 1800
rect 9620 1790 9700 1800
rect 9780 1790 9920 1800
rect 9980 1790 9990 1800
rect 2080 1780 2190 1790
rect 2820 1780 3160 1790
rect 4100 1780 4190 1790
rect 4360 1780 4370 1790
rect 4480 1780 4490 1790
rect 4740 1780 4750 1790
rect 4780 1780 4800 1790
rect 4820 1780 4830 1790
rect 4860 1780 4880 1790
rect 5000 1780 5020 1790
rect 5050 1780 5070 1790
rect 5150 1780 5170 1790
rect 5260 1780 5280 1790
rect 5320 1780 5340 1790
rect 7940 1780 8350 1790
rect 8620 1780 8910 1790
rect 9250 1780 9270 1790
rect 9280 1780 9310 1790
rect 9340 1780 9690 1790
rect 9780 1780 9910 1790
rect 9970 1780 9990 1790
rect 2050 1770 2190 1780
rect 2320 1770 2330 1780
rect 2800 1770 3160 1780
rect 4090 1770 4200 1780
rect 4390 1770 4400 1780
rect 4480 1770 4490 1780
rect 4620 1770 4630 1780
rect 4730 1770 4750 1780
rect 4780 1770 4800 1780
rect 4820 1770 4830 1780
rect 4860 1770 4880 1780
rect 4990 1770 5010 1780
rect 5050 1770 5060 1780
rect 5140 1770 5160 1780
rect 5260 1770 5280 1780
rect 5320 1770 5340 1780
rect 5420 1770 5430 1780
rect 7070 1770 7080 1780
rect 7090 1770 7100 1780
rect 7930 1770 8350 1780
rect 8620 1770 8900 1780
rect 9240 1770 9320 1780
rect 9340 1770 9690 1780
rect 9780 1770 9910 1780
rect 9970 1770 9990 1780
rect 2040 1760 2200 1770
rect 2300 1760 2360 1770
rect 2780 1760 3170 1770
rect 4080 1760 4210 1770
rect 4390 1760 4400 1770
rect 4480 1760 4490 1770
rect 4620 1760 4630 1770
rect 4730 1760 4750 1770
rect 4860 1760 4880 1770
rect 4990 1760 5010 1770
rect 5050 1760 5060 1770
rect 5140 1760 5160 1770
rect 5260 1760 5280 1770
rect 5310 1760 5330 1770
rect 5410 1760 5430 1770
rect 5450 1760 5470 1770
rect 7040 1760 7110 1770
rect 7940 1760 8350 1770
rect 8610 1760 8920 1770
rect 9100 1760 9110 1770
rect 9240 1760 9360 1770
rect 9390 1760 9410 1770
rect 9430 1760 9700 1770
rect 9780 1760 9830 1770
rect 9850 1760 9920 1770
rect 9970 1760 9990 1770
rect 2030 1750 2210 1760
rect 2240 1750 2370 1760
rect 2760 1750 3170 1760
rect 4080 1750 4220 1760
rect 4390 1750 4400 1760
rect 4480 1750 4490 1760
rect 4550 1750 4560 1760
rect 4620 1750 4640 1760
rect 4730 1750 4740 1760
rect 4870 1750 4880 1760
rect 4990 1750 5010 1760
rect 5040 1750 5060 1760
rect 5140 1750 5150 1760
rect 5250 1750 5280 1760
rect 5310 1750 5330 1760
rect 5400 1750 5430 1760
rect 5460 1750 5480 1760
rect 7050 1750 7110 1760
rect 7940 1750 8350 1760
rect 8610 1750 8920 1760
rect 9090 1750 9110 1760
rect 9230 1750 9370 1760
rect 9390 1750 9410 1760
rect 9430 1750 9700 1760
rect 9780 1750 9830 1760
rect 9850 1750 9930 1760
rect 9960 1750 9990 1760
rect 2030 1740 2390 1750
rect 2730 1740 3150 1750
rect 4070 1740 4220 1750
rect 4290 1740 4300 1750
rect 4380 1740 4400 1750
rect 4480 1740 4500 1750
rect 4540 1740 4570 1750
rect 4630 1740 4640 1750
rect 4720 1740 4740 1750
rect 4870 1740 4880 1750
rect 4990 1740 5010 1750
rect 5040 1740 5060 1750
rect 5130 1740 5150 1750
rect 5250 1740 5270 1750
rect 5300 1740 5320 1750
rect 5390 1740 5420 1750
rect 5470 1740 5500 1750
rect 7040 1740 7120 1750
rect 7940 1740 8350 1750
rect 8610 1740 8910 1750
rect 9090 1740 9110 1750
rect 9210 1740 9390 1750
rect 9420 1740 9550 1750
rect 9560 1740 9710 1750
rect 9780 1740 9830 1750
rect 9850 1740 9920 1750
rect 9960 1740 9990 1750
rect 2040 1730 2410 1740
rect 2710 1730 3150 1740
rect 4070 1730 4220 1740
rect 4290 1730 4300 1740
rect 4370 1730 4380 1740
rect 4480 1730 4500 1740
rect 4540 1730 4550 1740
rect 4560 1730 4580 1740
rect 4630 1730 4650 1740
rect 4720 1730 4740 1740
rect 4870 1730 4880 1740
rect 4980 1730 5000 1740
rect 5040 1730 5050 1740
rect 5130 1730 5140 1740
rect 5240 1730 5270 1740
rect 5300 1730 5320 1740
rect 5390 1730 5410 1740
rect 5490 1730 5510 1740
rect 7020 1730 7030 1740
rect 7040 1730 7130 1740
rect 7950 1730 8340 1740
rect 8600 1730 8910 1740
rect 9090 1730 9110 1740
rect 9200 1730 9390 1740
rect 9410 1730 9540 1740
rect 9550 1730 9570 1740
rect 9580 1730 9710 1740
rect 9790 1730 9830 1740
rect 9860 1730 9910 1740
rect 9940 1730 9990 1740
rect 2020 1720 2030 1730
rect 2040 1720 2440 1730
rect 2690 1720 3140 1730
rect 4070 1720 4180 1730
rect 4290 1720 4300 1730
rect 4480 1720 4500 1730
rect 4540 1720 4550 1730
rect 4570 1720 4580 1730
rect 4630 1720 4650 1730
rect 4710 1720 4730 1730
rect 4770 1720 4820 1730
rect 4870 1720 4880 1730
rect 4980 1720 5000 1730
rect 5030 1720 5050 1730
rect 5120 1720 5140 1730
rect 5240 1720 5260 1730
rect 5290 1720 5310 1730
rect 5380 1720 5400 1730
rect 5500 1720 5520 1730
rect 7010 1720 7150 1730
rect 7950 1720 8340 1730
rect 8600 1720 8900 1730
rect 9090 1720 9110 1730
rect 9200 1720 9540 1730
rect 9580 1720 9710 1730
rect 9800 1720 9830 1730
rect 9870 1720 9910 1730
rect 9940 1720 9990 1730
rect 2020 1710 2030 1720
rect 2040 1710 2460 1720
rect 2670 1710 3140 1720
rect 4090 1710 4150 1720
rect 4480 1710 4500 1720
rect 4540 1710 4550 1720
rect 4570 1710 4590 1720
rect 4640 1710 4650 1720
rect 4710 1710 4730 1720
rect 4770 1710 4830 1720
rect 4870 1710 4890 1720
rect 4970 1710 4990 1720
rect 5030 1710 5040 1720
rect 5120 1710 5140 1720
rect 5230 1710 5250 1720
rect 5290 1710 5310 1720
rect 5370 1710 5390 1720
rect 5510 1710 5540 1720
rect 7010 1710 7150 1720
rect 7950 1710 8340 1720
rect 8610 1710 8870 1720
rect 9090 1710 9110 1720
rect 9220 1710 9320 1720
rect 9330 1710 9650 1720
rect 9660 1710 9700 1720
rect 9790 1710 9840 1720
rect 9860 1710 9900 1720
rect 9930 1710 9990 1720
rect 2020 1700 2030 1710
rect 2050 1700 2480 1710
rect 2660 1700 3130 1710
rect 4100 1700 4120 1710
rect 4480 1700 4490 1710
rect 4540 1700 4550 1710
rect 4580 1700 4590 1710
rect 4640 1700 4660 1710
rect 4710 1700 4720 1710
rect 4760 1700 4780 1710
rect 4820 1700 4830 1710
rect 4870 1700 4890 1710
rect 4970 1700 4990 1710
rect 5110 1700 5130 1710
rect 5230 1700 5250 1710
rect 5280 1700 5300 1710
rect 5370 1700 5390 1710
rect 5440 1700 5450 1710
rect 5460 1700 5470 1710
rect 5520 1700 5540 1710
rect 7010 1700 7120 1710
rect 7950 1700 8340 1710
rect 8610 1700 8850 1710
rect 9080 1700 9110 1710
rect 9220 1700 9320 1710
rect 9330 1700 9710 1710
rect 9790 1700 9900 1710
rect 9930 1700 9990 1710
rect 2030 1690 2480 1700
rect 2660 1690 3120 1700
rect 4490 1690 4500 1700
rect 4540 1690 4550 1700
rect 4580 1690 4600 1700
rect 4650 1690 4660 1700
rect 4700 1690 4720 1700
rect 4760 1690 4770 1700
rect 4820 1690 4830 1700
rect 4870 1690 4890 1700
rect 4970 1690 4990 1700
rect 5110 1690 5130 1700
rect 5220 1690 5240 1700
rect 5280 1690 5300 1700
rect 5360 1690 5380 1700
rect 5430 1690 5450 1700
rect 5460 1690 5480 1700
rect 5530 1690 5550 1700
rect 7020 1690 7130 1700
rect 7950 1690 8340 1700
rect 8610 1690 8850 1700
rect 9080 1690 9110 1700
rect 9230 1690 9350 1700
rect 9360 1690 9710 1700
rect 9800 1690 9890 1700
rect 9920 1690 9990 1700
rect 2030 1680 2480 1690
rect 2660 1680 3110 1690
rect 4490 1680 4500 1690
rect 4590 1680 4600 1690
rect 4650 1680 4660 1690
rect 4700 1680 4710 1690
rect 4750 1680 4770 1690
rect 4870 1680 4890 1690
rect 4960 1680 4980 1690
rect 5110 1680 5120 1690
rect 5220 1680 5240 1690
rect 5270 1680 5290 1690
rect 5350 1680 5370 1690
rect 5420 1680 5440 1690
rect 5470 1680 5480 1690
rect 5530 1680 5550 1690
rect 7020 1680 7130 1690
rect 7960 1680 8340 1690
rect 8620 1680 8860 1690
rect 9080 1680 9110 1690
rect 9220 1680 9350 1690
rect 9370 1680 9700 1690
rect 9800 1680 9880 1690
rect 9920 1680 9990 1690
rect 2040 1670 2470 1680
rect 2660 1670 2710 1680
rect 2720 1670 3110 1680
rect 4240 1670 4250 1680
rect 4390 1670 4400 1680
rect 4410 1670 4440 1680
rect 4590 1670 4610 1680
rect 4650 1670 4670 1680
rect 4700 1670 4710 1680
rect 4750 1670 4760 1680
rect 4870 1670 4890 1680
rect 4960 1670 4980 1680
rect 5020 1670 5030 1680
rect 5100 1670 5120 1680
rect 5210 1670 5230 1680
rect 5270 1670 5290 1680
rect 5340 1670 5370 1680
rect 5410 1670 5430 1680
rect 5470 1670 5490 1680
rect 5530 1670 5550 1680
rect 7020 1670 7140 1680
rect 7970 1670 8330 1680
rect 8620 1670 8840 1680
rect 9080 1670 9120 1680
rect 9210 1670 9530 1680
rect 9550 1670 9710 1680
rect 9800 1670 9880 1680
rect 9920 1670 9990 1680
rect 2050 1660 2450 1670
rect 2720 1660 3100 1670
rect 4390 1660 4400 1670
rect 4440 1660 4450 1670
rect 4480 1660 4490 1670
rect 4600 1660 4630 1670
rect 4650 1660 4670 1670
rect 4700 1660 4720 1670
rect 4740 1660 4760 1670
rect 4860 1660 4890 1670
rect 4960 1660 4980 1670
rect 5010 1660 5030 1670
rect 5100 1660 5120 1670
rect 5210 1660 5230 1670
rect 5260 1660 5280 1670
rect 5330 1660 5360 1670
rect 5400 1660 5430 1670
rect 5470 1660 5490 1670
rect 5530 1660 5550 1670
rect 7010 1660 7140 1670
rect 7970 1660 8330 1670
rect 8630 1660 8830 1670
rect 9080 1660 9120 1670
rect 9200 1660 9530 1670
rect 9540 1660 9610 1670
rect 9630 1660 9670 1670
rect 9690 1660 9710 1670
rect 9800 1660 9880 1670
rect 9910 1660 9960 1670
rect 9970 1660 9990 1670
rect 2050 1650 2420 1660
rect 2740 1650 3100 1660
rect 4250 1650 4260 1660
rect 4300 1650 4310 1660
rect 4440 1650 4450 1660
rect 4480 1650 4500 1660
rect 4610 1650 4640 1660
rect 4730 1650 4750 1660
rect 4840 1650 4890 1660
rect 4960 1650 4980 1660
rect 5010 1650 5020 1660
rect 5200 1650 5220 1660
rect 5260 1650 5280 1660
rect 5320 1650 5350 1660
rect 5400 1650 5420 1660
rect 5460 1650 5490 1660
rect 5530 1650 5550 1660
rect 7000 1650 7140 1660
rect 7970 1650 8330 1660
rect 8630 1650 8830 1660
rect 9080 1650 9120 1660
rect 9210 1650 9620 1660
rect 9630 1650 9660 1660
rect 9680 1650 9870 1660
rect 9900 1650 9950 1660
rect 9970 1650 9990 1660
rect 2060 1640 2420 1650
rect 2730 1640 3090 1650
rect 4300 1640 4310 1650
rect 4440 1640 4450 1650
rect 4490 1640 4530 1650
rect 4960 1640 4980 1650
rect 5010 1640 5020 1650
rect 5170 1640 5210 1650
rect 5250 1640 5270 1650
rect 5310 1640 5340 1650
rect 5410 1640 5430 1650
rect 5440 1640 5480 1650
rect 5530 1640 5550 1650
rect 7000 1640 7150 1650
rect 7980 1640 8330 1650
rect 8620 1640 8630 1650
rect 8650 1640 8820 1650
rect 9080 1640 9120 1650
rect 9230 1640 9860 1650
rect 9900 1640 9950 1650
rect 9970 1640 9990 1650
rect 2070 1630 2390 1640
rect 2750 1630 2760 1640
rect 2770 1630 3090 1640
rect 4430 1630 4450 1640
rect 4510 1630 4520 1640
rect 4960 1630 4980 1640
rect 4990 1630 5020 1640
rect 5100 1630 5120 1640
rect 5180 1630 5200 1640
rect 5240 1630 5270 1640
rect 5300 1630 5330 1640
rect 5410 1630 5470 1640
rect 5520 1630 5540 1640
rect 7000 1630 7150 1640
rect 7970 1630 8320 1640
rect 8620 1630 8630 1640
rect 8650 1630 8820 1640
rect 9080 1630 9120 1640
rect 9230 1630 9810 1640
rect 9890 1630 9950 1640
rect 9960 1630 9990 1640
rect 2070 1620 2370 1630
rect 2750 1620 2760 1630
rect 2770 1620 3070 1630
rect 4390 1620 4410 1630
rect 5110 1620 5130 1630
rect 5240 1620 5260 1630
rect 5290 1620 5320 1630
rect 5430 1620 5450 1630
rect 5510 1620 5540 1630
rect 7000 1620 7140 1630
rect 7970 1620 8320 1630
rect 8640 1620 8790 1630
rect 8800 1620 8810 1630
rect 9070 1620 9120 1630
rect 9270 1620 9710 1630
rect 9740 1620 9800 1630
rect 9840 1620 9850 1630
rect 9880 1620 9940 1630
rect 9950 1620 9990 1630
rect 2080 1610 2380 1620
rect 2750 1610 3060 1620
rect 4360 1610 4380 1620
rect 5110 1610 5130 1620
rect 5230 1610 5250 1620
rect 5290 1610 5310 1620
rect 5500 1610 5530 1620
rect 5620 1610 5650 1620
rect 7000 1610 7140 1620
rect 7960 1610 8320 1620
rect 8640 1610 8660 1620
rect 8700 1610 8790 1620
rect 9070 1610 9120 1620
rect 9250 1610 9370 1620
rect 9430 1610 9700 1620
rect 9740 1610 9840 1620
rect 9880 1610 9940 1620
rect 9950 1610 9990 1620
rect 2090 1600 2370 1610
rect 2730 1600 3060 1610
rect 5120 1600 5140 1610
rect 5220 1600 5240 1610
rect 5280 1600 5310 1610
rect 5360 1600 5400 1610
rect 5490 1600 5520 1610
rect 5590 1600 5670 1610
rect 7000 1600 7140 1610
rect 7950 1600 7960 1610
rect 7970 1600 8320 1610
rect 8610 1600 8630 1610
rect 8640 1600 8660 1610
rect 8710 1600 8780 1610
rect 9070 1600 9120 1610
rect 9170 1600 9380 1610
rect 9430 1600 9840 1610
rect 9870 1600 9930 1610
rect 9940 1600 9990 1610
rect 2100 1590 2370 1600
rect 2720 1590 3050 1600
rect 4280 1590 4290 1600
rect 5160 1590 5230 1600
rect 5270 1590 5300 1600
rect 5350 1590 5420 1600
rect 5470 1590 5510 1600
rect 5580 1590 5620 1600
rect 5660 1590 5690 1600
rect 7000 1590 7010 1600
rect 7030 1590 7130 1600
rect 7950 1590 7960 1600
rect 7970 1590 8320 1600
rect 8600 1590 8610 1600
rect 8620 1590 8660 1600
rect 8740 1590 8750 1600
rect 8760 1590 8770 1600
rect 9070 1590 9830 1600
rect 9870 1590 9920 1600
rect 9940 1590 9990 1600
rect 2110 1580 2370 1590
rect 2710 1580 3030 1590
rect 4280 1580 4300 1590
rect 5160 1580 5210 1590
rect 5260 1580 5290 1590
rect 5340 1580 5360 1590
rect 5410 1580 5420 1590
rect 5460 1580 5490 1590
rect 5580 1580 5590 1590
rect 5670 1580 5700 1590
rect 7030 1580 7130 1590
rect 7970 1580 8310 1590
rect 8620 1580 8670 1590
rect 9070 1580 9310 1590
rect 9330 1580 9830 1590
rect 9870 1580 9920 1590
rect 9940 1580 9960 1590
rect 9970 1580 9980 1590
rect 9990 1580 9990 1590
rect 2110 1570 2370 1580
rect 2700 1570 3000 1580
rect 4280 1570 4310 1580
rect 5260 1570 5280 1580
rect 5340 1570 5360 1580
rect 5570 1570 5590 1580
rect 5680 1570 5700 1580
rect 7000 1570 7150 1580
rect 7970 1570 8310 1580
rect 8610 1570 8660 1580
rect 9070 1570 9300 1580
rect 9340 1570 9820 1580
rect 9860 1570 9910 1580
rect 9990 1570 9990 1580
rect 2140 1560 2380 1570
rect 2680 1560 2990 1570
rect 4280 1560 4310 1570
rect 5260 1560 5270 1570
rect 5570 1560 5580 1570
rect 5640 1560 5660 1570
rect 5690 1560 5710 1570
rect 7000 1560 7160 1570
rect 7990 1560 8310 1570
rect 8580 1560 8600 1570
rect 8620 1560 8660 1570
rect 9070 1560 9720 1570
rect 9810 1560 9820 1570
rect 9860 1560 9910 1570
rect 2140 1550 2440 1560
rect 2520 1550 2960 1560
rect 4280 1550 4320 1560
rect 5570 1550 5580 1560
rect 5640 1550 5670 1560
rect 5700 1550 5720 1560
rect 7000 1550 7180 1560
rect 8000 1550 8300 1560
rect 8590 1550 8670 1560
rect 9070 1550 9710 1560
rect 9850 1550 9900 1560
rect 2160 1540 2950 1550
rect 4270 1540 4320 1550
rect 5280 1540 5300 1550
rect 5310 1540 5320 1550
rect 5570 1540 5580 1550
rect 5610 1540 5630 1550
rect 5660 1540 5680 1550
rect 5710 1540 5720 1550
rect 6980 1540 6990 1550
rect 7000 1540 7180 1550
rect 8000 1540 8300 1550
rect 8580 1540 8660 1550
rect 9060 1540 9580 1550
rect 9600 1540 9710 1550
rect 9850 1540 9900 1550
rect 2170 1530 2940 1540
rect 4270 1530 4330 1540
rect 5280 1530 5320 1540
rect 5560 1530 5580 1540
rect 5610 1530 5630 1540
rect 5660 1530 5680 1540
rect 5710 1530 5720 1540
rect 6980 1530 7170 1540
rect 8000 1530 8300 1540
rect 8620 1530 8670 1540
rect 9060 1530 9470 1540
rect 9540 1530 9710 1540
rect 9840 1530 9890 1540
rect 9910 1530 9930 1540
rect 9960 1530 9980 1540
rect 2180 1520 2930 1530
rect 4260 1520 4330 1530
rect 5290 1520 5310 1530
rect 5560 1520 5580 1530
rect 5610 1520 5630 1530
rect 5660 1520 5680 1530
rect 5710 1520 5720 1530
rect 6990 1520 7170 1530
rect 7190 1520 7220 1530
rect 8010 1520 8300 1530
rect 8650 1520 8670 1530
rect 9070 1520 9490 1530
rect 9510 1520 9710 1530
rect 9830 1520 9890 1530
rect 9910 1520 9930 1530
rect 9960 1520 9980 1530
rect 2190 1510 2920 1520
rect 4250 1510 4340 1520
rect 5560 1510 5580 1520
rect 5610 1510 5620 1520
rect 5660 1510 5680 1520
rect 5710 1510 5720 1520
rect 6990 1510 7210 1520
rect 8020 1510 8290 1520
rect 8650 1510 8670 1520
rect 9060 1510 9180 1520
rect 9210 1510 9490 1520
rect 9510 1510 9700 1520
rect 9830 1510 9880 1520
rect 9910 1510 9930 1520
rect 2210 1500 2920 1510
rect 4250 1500 4340 1510
rect 5460 1500 5490 1510
rect 5560 1500 5580 1510
rect 5610 1500 5620 1510
rect 5660 1500 5680 1510
rect 5700 1500 5720 1510
rect 6980 1500 7200 1510
rect 8020 1500 8290 1510
rect 8640 1500 8680 1510
rect 9060 1500 9130 1510
rect 9200 1500 9230 1510
rect 9240 1500 9360 1510
rect 9370 1500 9410 1510
rect 9430 1500 9490 1510
rect 9500 1500 9590 1510
rect 9600 1500 9710 1510
rect 9830 1500 9880 1510
rect 9910 1500 9930 1510
rect 9940 1500 9960 1510
rect 2210 1490 2910 1500
rect 4250 1490 4350 1500
rect 5460 1490 5500 1500
rect 5560 1490 5580 1500
rect 5610 1490 5620 1500
rect 5670 1490 5690 1500
rect 5700 1490 5720 1500
rect 6960 1490 6970 1500
rect 6980 1490 7190 1500
rect 7200 1490 7220 1500
rect 8000 1490 8290 1500
rect 8640 1490 8670 1500
rect 8680 1490 8690 1500
rect 9070 1490 9130 1500
rect 9200 1490 9220 1500
rect 9240 1490 9350 1500
rect 9370 1490 9720 1500
rect 9820 1490 9870 1500
rect 9940 1490 9990 1500
rect 2220 1480 2900 1490
rect 4140 1480 4150 1490
rect 4260 1480 4350 1490
rect 5480 1480 5490 1490
rect 5560 1480 5580 1490
rect 5610 1480 5620 1490
rect 5680 1480 5690 1490
rect 5700 1480 5710 1490
rect 6960 1480 7230 1490
rect 7240 1480 7250 1490
rect 7990 1480 8270 1490
rect 8610 1480 8670 1490
rect 8680 1480 8720 1490
rect 9070 1480 9130 1490
rect 9190 1480 9210 1490
rect 9240 1480 9340 1490
rect 9370 1480 9570 1490
rect 9580 1480 9720 1490
rect 9810 1480 9860 1490
rect 9930 1480 9990 1490
rect 2220 1470 2890 1480
rect 4260 1470 4350 1480
rect 5560 1470 5580 1480
rect 5610 1470 5620 1480
rect 6960 1470 7260 1480
rect 8000 1470 8270 1480
rect 8590 1470 8690 1480
rect 8700 1470 8720 1480
rect 9070 1470 9130 1480
rect 9180 1470 9210 1480
rect 9230 1470 9570 1480
rect 9580 1470 9590 1480
rect 9640 1470 9710 1480
rect 9810 1470 9860 1480
rect 9880 1470 9910 1480
rect 9920 1470 9990 1480
rect 2230 1460 2880 1470
rect 4150 1460 4160 1470
rect 4270 1460 4360 1470
rect 5450 1460 5460 1470
rect 5500 1460 5510 1470
rect 5560 1460 5570 1470
rect 5610 1460 5620 1470
rect 6930 1460 7250 1470
rect 8010 1460 8270 1470
rect 8590 1460 8750 1470
rect 9070 1460 9090 1470
rect 9100 1460 9130 1470
rect 9170 1460 9520 1470
rect 9530 1460 9580 1470
rect 9650 1460 9710 1470
rect 9800 1460 9990 1470
rect 2240 1450 2870 1460
rect 4270 1450 4360 1460
rect 5450 1450 5460 1460
rect 5500 1450 5510 1460
rect 5560 1450 5570 1460
rect 5610 1450 5620 1460
rect 6930 1450 7230 1460
rect 8010 1450 8260 1460
rect 8590 1450 8700 1460
rect 8710 1450 8720 1460
rect 9070 1450 9080 1460
rect 9110 1450 9130 1460
rect 9160 1450 9580 1460
rect 9650 1450 9710 1460
rect 9790 1450 9950 1460
rect 9960 1450 9990 1460
rect 2240 1440 2850 1450
rect 4280 1440 4370 1450
rect 5450 1440 5470 1450
rect 5500 1440 5510 1450
rect 5550 1440 5570 1450
rect 5610 1440 5620 1450
rect 6920 1440 7230 1450
rect 7250 1440 7260 1450
rect 8010 1440 8260 1450
rect 8590 1440 8620 1450
rect 8630 1440 8690 1450
rect 9110 1440 9130 1450
rect 9150 1440 9340 1450
rect 9350 1440 9360 1450
rect 9380 1440 9390 1450
rect 9410 1440 9580 1450
rect 9590 1440 9600 1450
rect 9640 1440 9700 1450
rect 9790 1440 9950 1450
rect 9970 1440 9990 1450
rect 2250 1430 2850 1440
rect 4290 1430 4370 1440
rect 5450 1430 5470 1440
rect 5500 1430 5510 1440
rect 5550 1430 5570 1440
rect 5610 1430 5620 1440
rect 6880 1430 6900 1440
rect 6910 1430 7260 1440
rect 8010 1430 8240 1440
rect 8580 1430 8610 1440
rect 8640 1430 8700 1440
rect 9070 1430 9080 1440
rect 9110 1430 9350 1440
rect 9370 1430 9510 1440
rect 9560 1430 9580 1440
rect 9590 1430 9610 1440
rect 9650 1430 9700 1440
rect 9780 1430 9840 1440
rect 9850 1430 9990 1440
rect 2260 1420 2840 1430
rect 4160 1420 4170 1430
rect 4290 1420 4370 1430
rect 5450 1420 5470 1430
rect 5500 1420 5520 1430
rect 5540 1420 5560 1430
rect 5600 1420 5620 1430
rect 6860 1420 7270 1430
rect 8010 1420 8230 1430
rect 8590 1420 8610 1430
rect 8680 1420 8690 1430
rect 9070 1420 9080 1430
rect 9110 1420 9350 1430
rect 9370 1420 9490 1430
rect 9560 1420 9580 1430
rect 9590 1420 9610 1430
rect 9650 1420 9700 1430
rect 9770 1420 9830 1430
rect 9850 1420 9990 1430
rect 2270 1410 2830 1420
rect 4160 1410 4170 1420
rect 4290 1410 4380 1420
rect 5460 1410 5480 1420
rect 5510 1410 5550 1420
rect 5600 1410 5610 1420
rect 6860 1410 7270 1420
rect 7990 1410 8060 1420
rect 8070 1410 8220 1420
rect 8600 1410 8620 1420
rect 9110 1410 9240 1420
rect 9250 1410 9410 1420
rect 9420 1410 9490 1420
rect 9510 1410 9530 1420
rect 9550 1410 9620 1420
rect 9650 1410 9690 1420
rect 9770 1410 9930 1420
rect 9950 1410 9970 1420
rect 9990 1410 9990 1420
rect 2290 1400 2820 1410
rect 4310 1400 4380 1410
rect 5460 1400 5480 1410
rect 5590 1400 5610 1410
rect 6860 1400 7270 1410
rect 7990 1400 8040 1410
rect 8050 1400 8210 1410
rect 9110 1400 9230 1410
rect 9250 1400 9290 1410
rect 9310 1400 9590 1410
rect 9600 1400 9620 1410
rect 9640 1400 9690 1410
rect 9760 1400 9870 1410
rect 9880 1400 9930 1410
rect 9950 1400 9960 1410
rect 9990 1400 9990 1410
rect 2300 1390 2810 1400
rect 4320 1390 4380 1400
rect 5470 1390 5490 1400
rect 5590 1390 5610 1400
rect 6850 1390 7260 1400
rect 8010 1390 8170 1400
rect 8180 1390 8200 1400
rect 9110 1390 9220 1400
rect 9270 1390 9280 1400
rect 9310 1390 9590 1400
rect 9600 1390 9620 1400
rect 9640 1390 9690 1400
rect 9760 1390 9810 1400
rect 9830 1390 9860 1400
rect 9870 1390 9930 1400
rect 2310 1380 2800 1390
rect 4330 1380 4390 1390
rect 5470 1380 5490 1390
rect 5580 1380 5600 1390
rect 6850 1380 7270 1390
rect 8010 1380 8190 1390
rect 9110 1380 9210 1390
rect 9300 1380 9540 1390
rect 9560 1380 9620 1390
rect 9650 1380 9680 1390
rect 9750 1380 9810 1390
rect 9830 1380 9920 1390
rect 2320 1370 2780 1380
rect 4330 1370 4390 1380
rect 5510 1370 5520 1380
rect 5570 1370 5590 1380
rect 6860 1370 7270 1380
rect 8010 1370 8170 1380
rect 9110 1370 9200 1380
rect 9290 1370 9520 1380
rect 9550 1370 9570 1380
rect 9610 1370 9680 1380
rect 9750 1370 9800 1380
rect 9830 1370 9870 1380
rect 9920 1370 9930 1380
rect 9950 1370 9960 1380
rect 2340 1360 2770 1370
rect 4340 1360 4400 1370
rect 5500 1360 5580 1370
rect 6850 1360 7260 1370
rect 8010 1360 8160 1370
rect 9110 1360 9200 1370
rect 9270 1360 9310 1370
rect 9330 1360 9460 1370
rect 9470 1360 9590 1370
rect 9620 1360 9680 1370
rect 9740 1360 9800 1370
rect 9830 1360 9900 1370
rect 9920 1360 9960 1370
rect 2370 1350 2760 1360
rect 3570 1350 3600 1360
rect 4340 1350 4400 1360
rect 5510 1350 5580 1360
rect 6850 1350 7260 1360
rect 8020 1350 8150 1360
rect 9120 1350 9190 1360
rect 9270 1350 9590 1360
rect 9610 1350 9670 1360
rect 9740 1350 9790 1360
rect 9830 1350 9960 1360
rect 2390 1340 2730 1350
rect 3550 1340 3630 1350
rect 4340 1340 4400 1350
rect 6850 1340 7270 1350
rect 7280 1340 7290 1350
rect 8040 1340 8130 1350
rect 9120 1340 9180 1350
rect 9270 1340 9600 1350
rect 9620 1340 9640 1350
rect 9740 1340 9790 1350
rect 9840 1340 9950 1350
rect 2410 1330 2720 1340
rect 3530 1330 3640 1340
rect 4330 1330 4400 1340
rect 6850 1330 7290 1340
rect 8050 1330 8110 1340
rect 9120 1330 9170 1340
rect 9270 1330 9480 1340
rect 9490 1330 9620 1340
rect 9630 1330 9640 1340
rect 9730 1330 9770 1340
rect 9840 1330 9960 1340
rect 2440 1320 2700 1330
rect 3530 1320 3650 1330
rect 4290 1320 4410 1330
rect 6850 1320 7300 1330
rect 8010 1320 8030 1330
rect 8060 1320 8080 1330
rect 9120 1320 9160 1330
rect 9270 1320 9380 1330
rect 9400 1320 9450 1330
rect 9470 1320 9640 1330
rect 9720 1320 9760 1330
rect 9840 1320 9990 1330
rect 2530 1310 2660 1320
rect 3520 1310 3670 1320
rect 4290 1310 4410 1320
rect 6850 1310 7280 1320
rect 7290 1310 7310 1320
rect 8020 1310 8030 1320
rect 9120 1310 9150 1320
rect 9270 1310 9640 1320
rect 9710 1310 9760 1320
rect 9840 1310 9920 1320
rect 9940 1310 9990 1320
rect 3510 1300 3680 1310
rect 4290 1300 4420 1310
rect 6850 1300 7310 1310
rect 9120 1300 9140 1310
rect 9260 1300 9670 1310
rect 9710 1300 9760 1310
rect 9850 1300 9980 1310
rect 3510 1290 3690 1300
rect 4250 1290 4260 1300
rect 4290 1290 4420 1300
rect 6850 1290 7290 1300
rect 7300 1290 7310 1300
rect 9120 1290 9130 1300
rect 9260 1290 9580 1300
rect 9600 1290 9610 1300
rect 9620 1290 9670 1300
rect 9700 1290 9760 1300
rect 9860 1290 9960 1300
rect 3510 1280 3700 1290
rect 4240 1280 4270 1290
rect 4290 1280 4420 1290
rect 6850 1280 7290 1290
rect 9270 1280 9480 1290
rect 9500 1280 9660 1290
rect 9700 1280 9750 1290
rect 9840 1280 9950 1290
rect 3510 1270 3720 1280
rect 4210 1270 4420 1280
rect 6850 1270 7300 1280
rect 9120 1270 9130 1280
rect 9310 1270 9460 1280
rect 9470 1270 9480 1280
rect 9500 1270 9650 1280
rect 9700 1270 9750 1280
rect 9840 1270 9890 1280
rect 9910 1270 9950 1280
rect 3510 1260 3730 1270
rect 4210 1260 4430 1270
rect 5430 1260 5440 1270
rect 6850 1260 7290 1270
rect 9120 1260 9130 1270
rect 9330 1260 9400 1270
rect 9450 1260 9490 1270
rect 9500 1260 9650 1270
rect 9690 1260 9740 1270
rect 9840 1260 9880 1270
rect 9900 1260 9940 1270
rect 3610 1250 3620 1260
rect 3650 1250 3740 1260
rect 4210 1250 4430 1260
rect 5340 1250 5350 1260
rect 5370 1250 5380 1260
rect 6850 1250 7300 1260
rect 9120 1250 9130 1260
rect 9320 1250 9490 1260
rect 9510 1250 9590 1260
rect 9610 1250 9630 1260
rect 9680 1250 9730 1260
rect 9840 1250 9970 1260
rect 3670 1240 3750 1250
rect 4210 1240 4430 1250
rect 5210 1240 5220 1250
rect 5240 1240 5250 1250
rect 5270 1240 5280 1250
rect 5300 1240 5310 1250
rect 5320 1240 5330 1250
rect 5340 1240 5350 1250
rect 5370 1240 5380 1250
rect 5400 1240 5410 1250
rect 6850 1240 7300 1250
rect 9120 1240 9140 1250
rect 9320 1240 9600 1250
rect 9680 1240 9720 1250
rect 9830 1240 9910 1250
rect 9940 1240 9970 1250
rect 3680 1230 3760 1240
rect 4210 1230 4430 1240
rect 5110 1230 5130 1240
rect 5190 1230 5200 1240
rect 5210 1230 5220 1240
rect 5240 1230 5250 1240
rect 5270 1230 5280 1240
rect 5290 1230 5300 1240
rect 5320 1230 5330 1240
rect 5340 1230 5350 1240
rect 5370 1230 5380 1240
rect 6860 1230 7300 1240
rect 9120 1230 9130 1240
rect 9280 1230 9490 1240
rect 9520 1230 9610 1240
rect 9670 1230 9720 1240
rect 9820 1230 9900 1240
rect 3690 1220 3780 1230
rect 4210 1220 4440 1230
rect 5060 1220 5070 1230
rect 5190 1220 5200 1230
rect 5210 1220 5220 1230
rect 5240 1220 5260 1230
rect 5270 1220 5310 1230
rect 5330 1220 5350 1230
rect 5380 1220 5390 1230
rect 6850 1220 7300 1230
rect 9120 1220 9130 1230
rect 9280 1220 9490 1230
rect 9530 1220 9610 1230
rect 9670 1220 9720 1230
rect 9820 1220 9950 1230
rect 3700 1210 3800 1220
rect 4210 1210 4440 1220
rect 5000 1210 5010 1220
rect 5150 1210 5160 1220
rect 5190 1210 5210 1220
rect 5250 1210 5260 1220
rect 5280 1210 5310 1220
rect 5330 1210 5350 1220
rect 5400 1210 5410 1220
rect 5430 1210 5450 1220
rect 6860 1210 7300 1220
rect 9120 1210 9140 1220
rect 9280 1210 9310 1220
rect 9330 1210 9500 1220
rect 9530 1210 9620 1220
rect 9660 1210 9710 1220
rect 9830 1210 9880 1220
rect 9910 1210 9960 1220
rect 3720 1200 3810 1210
rect 4220 1200 4440 1210
rect 5000 1200 5010 1210
rect 5060 1200 5070 1210
rect 5200 1200 5210 1210
rect 5250 1200 5260 1210
rect 5290 1200 5300 1210
rect 6860 1200 7300 1210
rect 9120 1200 9140 1210
rect 9280 1200 9310 1210
rect 9320 1200 9510 1210
rect 9540 1200 9570 1210
rect 9590 1200 9600 1210
rect 9660 1200 9710 1210
rect 9830 1200 9850 1210
rect 9860 1200 9890 1210
rect 9930 1200 9940 1210
rect 3730 1190 3830 1200
rect 4220 1190 4450 1200
rect 4810 1190 4820 1200
rect 4870 1190 4880 1200
rect 4990 1190 5010 1200
rect 5110 1190 5120 1200
rect 6850 1190 7300 1200
rect 9120 1190 9140 1200
rect 9330 1190 9500 1200
rect 9540 1190 9610 1200
rect 9650 1190 9700 1200
rect 9830 1190 9840 1200
rect 9850 1190 9940 1200
rect 3750 1180 3840 1190
rect 4220 1180 4450 1190
rect 4770 1180 4780 1190
rect 4800 1180 4810 1190
rect 4990 1180 5020 1190
rect 5060 1180 5070 1190
rect 5110 1180 5120 1190
rect 6860 1180 7300 1190
rect 9120 1180 9140 1190
rect 9280 1180 9310 1190
rect 9380 1180 9500 1190
rect 9540 1180 9600 1190
rect 9650 1180 9700 1190
rect 9820 1180 9970 1190
rect 9980 1180 9990 1190
rect 3750 1170 3860 1180
rect 4220 1170 4450 1180
rect 4670 1170 4680 1180
rect 4710 1170 4720 1180
rect 4820 1170 4830 1180
rect 4990 1170 5000 1180
rect 5010 1170 5020 1180
rect 5030 1170 5040 1180
rect 6750 1170 6760 1180
rect 6860 1170 7300 1180
rect 9120 1170 9140 1180
rect 9280 1170 9320 1180
rect 9370 1170 9500 1180
rect 9550 1170 9600 1180
rect 9640 1170 9690 1180
rect 9820 1170 9990 1180
rect 3750 1160 3870 1170
rect 4220 1160 4450 1170
rect 4770 1160 4780 1170
rect 6710 1160 6750 1170
rect 6860 1160 7300 1170
rect 9120 1160 9140 1170
rect 9280 1160 9330 1170
rect 9370 1160 9510 1170
rect 9550 1160 9590 1170
rect 9640 1160 9680 1170
rect 9820 1160 9840 1170
rect 9870 1160 9990 1170
rect 3760 1150 3880 1160
rect 4230 1150 4450 1160
rect 4880 1150 4890 1160
rect 6690 1150 6770 1160
rect 6860 1150 7300 1160
rect 8090 1150 8100 1160
rect 9120 1150 9150 1160
rect 9290 1150 9330 1160
rect 9380 1150 9520 1160
rect 9560 1150 9590 1160
rect 9630 1150 9710 1160
rect 9830 1150 9850 1160
rect 9860 1150 9990 1160
rect 3750 1140 3900 1150
rect 4230 1140 4460 1150
rect 4700 1140 4710 1150
rect 4770 1140 4780 1150
rect 4800 1140 4810 1150
rect 6670 1140 6780 1150
rect 6850 1140 7310 1150
rect 8090 1140 8100 1150
rect 9120 1140 9150 1150
rect 9290 1140 9320 1150
rect 9390 1140 9520 1150
rect 9560 1140 9580 1150
rect 9620 1140 9710 1150
rect 9840 1140 9850 1150
rect 9860 1140 9890 1150
rect 9940 1140 9980 1150
rect 3750 1130 3910 1140
rect 4240 1130 4460 1140
rect 6650 1130 6770 1140
rect 6860 1130 7310 1140
rect 8070 1130 8100 1140
rect 9120 1130 9150 1140
rect 9290 1130 9340 1140
rect 9390 1130 9580 1140
rect 9620 1130 9710 1140
rect 9830 1130 9880 1140
rect 9940 1130 9990 1140
rect 3760 1120 3920 1130
rect 4240 1120 4460 1130
rect 4640 1120 4650 1130
rect 6630 1120 6780 1130
rect 6860 1120 7310 1130
rect 8070 1120 8100 1130
rect 9120 1120 9150 1130
rect 9290 1120 9350 1130
rect 9390 1120 9550 1130
rect 9560 1120 9570 1130
rect 9610 1120 9720 1130
rect 9820 1120 9870 1130
rect 9920 1120 9990 1130
rect 3770 1110 3940 1120
rect 4230 1110 4460 1120
rect 6620 1110 6780 1120
rect 6860 1110 7300 1120
rect 8060 1110 8090 1120
rect 9120 1110 9150 1120
rect 9290 1110 9350 1120
rect 9390 1110 9540 1120
rect 9610 1110 9720 1120
rect 9840 1110 9870 1120
rect 9910 1110 9990 1120
rect 3780 1100 3950 1110
rect 4230 1100 4470 1110
rect 6610 1100 6780 1110
rect 6860 1100 7300 1110
rect 8060 1100 8090 1110
rect 9120 1100 9150 1110
rect 9300 1100 9360 1110
rect 9410 1100 9530 1110
rect 9610 1100 9650 1110
rect 9670 1100 9720 1110
rect 9840 1100 9860 1110
rect 9910 1100 9990 1110
rect 3840 1090 3970 1100
rect 4230 1090 4470 1100
rect 6580 1090 6780 1100
rect 6850 1090 7310 1100
rect 8070 1090 8090 1100
rect 9120 1090 9150 1100
rect 9250 1090 9270 1100
rect 9300 1090 9360 1100
rect 9420 1090 9540 1100
rect 9590 1090 9640 1100
rect 9660 1090 9720 1100
rect 9830 1090 9850 1100
rect 9930 1090 9940 1100
rect 9950 1090 9990 1100
rect 3850 1080 3980 1090
rect 4230 1080 4470 1090
rect 6580 1080 6780 1090
rect 6860 1080 7310 1090
rect 8060 1080 8090 1090
rect 9120 1080 9150 1090
rect 9190 1080 9270 1090
rect 9300 1080 9360 1090
rect 9420 1080 9550 1090
rect 9590 1080 9630 1090
rect 9650 1080 9720 1090
rect 9830 1080 9850 1090
rect 3860 1070 4000 1080
rect 4230 1070 4480 1080
rect 6580 1070 6780 1080
rect 6860 1070 7300 1080
rect 8070 1070 8080 1080
rect 9140 1070 9160 1080
rect 9170 1070 9260 1080
rect 9300 1070 9360 1080
rect 9420 1070 9540 1080
rect 9580 1070 9720 1080
rect 9920 1070 9940 1080
rect 3670 1060 3680 1070
rect 3870 1060 4020 1070
rect 4230 1060 4480 1070
rect 6560 1060 6780 1070
rect 6860 1060 7300 1070
rect 8060 1060 8080 1070
rect 9140 1060 9260 1070
rect 9310 1060 9360 1070
rect 9420 1060 9530 1070
rect 9580 1060 9720 1070
rect 9860 1060 9880 1070
rect 9920 1060 9950 1070
rect 3680 1050 3690 1060
rect 3870 1050 4030 1060
rect 4230 1050 4480 1060
rect 6560 1050 6780 1060
rect 6850 1050 7300 1060
rect 8050 1050 8070 1060
rect 9140 1050 9250 1060
rect 9310 1050 9350 1060
rect 9420 1050 9530 1060
rect 9570 1050 9620 1060
rect 9630 1050 9720 1060
rect 9850 1050 9890 1060
rect 9930 1050 9940 1060
rect 3870 1040 4040 1050
rect 4230 1040 4550 1050
rect 6560 1040 6780 1050
rect 6860 1040 7320 1050
rect 8050 1040 8070 1050
rect 9110 1040 9120 1050
rect 9140 1040 9240 1050
rect 9310 1040 9360 1050
rect 9420 1040 9530 1050
rect 9570 1040 9710 1050
rect 9830 1040 9850 1050
rect 9870 1040 9900 1050
rect 3870 1030 4060 1040
rect 4230 1030 4580 1040
rect 6550 1030 6790 1040
rect 6870 1030 7320 1040
rect 8050 1030 8070 1040
rect 9140 1030 9240 1040
rect 9310 1030 9330 1040
rect 9340 1030 9380 1040
rect 9430 1030 9520 1040
rect 9560 1030 9710 1040
rect 9830 1030 9850 1040
rect 9870 1030 9910 1040
rect 9990 1030 9990 1040
rect 3870 1020 4070 1030
rect 4220 1020 4620 1030
rect 6540 1020 6790 1030
rect 6860 1020 7320 1030
rect 8050 1020 8070 1030
rect 9140 1020 9240 1030
rect 9260 1020 9380 1030
rect 9430 1020 9510 1030
rect 9560 1020 9720 1030
rect 9830 1020 9850 1030
rect 9870 1020 9930 1030
rect 9970 1020 9990 1030
rect 3870 1010 4090 1020
rect 4220 1010 4650 1020
rect 6540 1010 6790 1020
rect 6860 1010 7310 1020
rect 9150 1010 9220 1020
rect 9250 1010 9380 1020
rect 9430 1010 9510 1020
rect 9550 1010 9740 1020
rect 9830 1010 9930 1020
rect 9960 1010 9990 1020
rect 3870 1000 4110 1010
rect 4220 1000 4670 1010
rect 6540 1000 6790 1010
rect 6860 1000 7310 1010
rect 9150 1000 9220 1010
rect 9240 1000 9400 1010
rect 9430 1000 9500 1010
rect 9540 1000 9650 1010
rect 9660 1000 9740 1010
rect 9830 1000 9920 1010
rect 9960 1000 9990 1010
rect 3890 990 4120 1000
rect 4210 990 4700 1000
rect 6540 990 6790 1000
rect 6870 990 7310 1000
rect 9150 990 9220 1000
rect 9260 990 9410 1000
rect 9430 990 9490 1000
rect 9540 990 9730 1000
rect 9830 990 9950 1000
rect 9970 990 9990 1000
rect 3890 980 4140 990
rect 4200 980 4720 990
rect 6540 980 6790 990
rect 6860 980 7310 990
rect 9160 980 9220 990
rect 9250 980 9410 990
rect 9420 980 9490 990
rect 9540 980 9690 990
rect 9700 980 9730 990
rect 9830 980 9870 990
rect 9900 980 9990 990
rect 3880 970 4170 980
rect 4190 970 4740 980
rect 6540 970 6790 980
rect 6860 970 7310 980
rect 9160 970 9480 980
rect 9530 970 9720 980
rect 9730 970 9760 980
rect 9790 970 9810 980
rect 9840 970 9870 980
rect 9920 970 9950 980
rect 9960 970 9990 980
rect 3870 960 4760 970
rect 6540 960 6800 970
rect 6860 960 7310 970
rect 9160 960 9200 970
rect 9220 960 9480 970
rect 9520 960 9750 970
rect 9780 960 9810 970
rect 9850 960 9990 970
rect 3870 950 4780 960
rect 5460 950 5480 960
rect 5500 950 5510 960
rect 5530 950 5540 960
rect 5800 950 5810 960
rect 6540 950 6800 960
rect 6860 950 7310 960
rect 9160 950 9210 960
rect 9260 950 9470 960
rect 9520 950 9750 960
rect 9760 950 9850 960
rect 9860 950 9990 960
rect 3870 940 4800 950
rect 5370 940 5380 950
rect 5410 940 5420 950
rect 5460 940 5470 950
rect 5500 940 5510 950
rect 5530 940 5540 950
rect 5570 940 5580 950
rect 5640 940 5650 950
rect 6560 940 6800 950
rect 6880 940 7320 950
rect 9160 940 9190 950
rect 9200 940 9210 950
rect 9260 940 9470 950
rect 9520 940 9990 950
rect 3870 930 4810 940
rect 5370 930 5380 940
rect 5420 930 5430 940
rect 5620 930 5630 940
rect 6550 930 6810 940
rect 6880 930 7320 940
rect 9170 930 9190 940
rect 9260 930 9460 940
rect 9510 930 9800 940
rect 9810 930 9990 940
rect 710 920 720 930
rect 3880 920 4820 930
rect 5370 920 5380 930
rect 5430 920 5440 930
rect 5530 920 5540 930
rect 5550 920 5560 930
rect 6560 920 6810 930
rect 6880 920 7310 930
rect 9170 920 9210 930
rect 9240 920 9460 930
rect 9500 920 9990 930
rect 700 910 710 920
rect 3890 910 4630 920
rect 4640 910 4830 920
rect 5370 910 5390 920
rect 5430 910 5440 920
rect 5530 910 5540 920
rect 6560 910 6810 920
rect 6890 910 7320 920
rect 9170 910 9450 920
rect 9500 910 9660 920
rect 9670 910 9990 920
rect 700 900 710 910
rect 3820 900 3830 910
rect 3900 900 3980 910
rect 4040 900 4620 910
rect 4640 900 4840 910
rect 5430 900 5440 910
rect 5480 900 5490 910
rect 5530 900 5540 910
rect 6560 900 6810 910
rect 6870 900 7310 910
rect 9170 900 9450 910
rect 9490 900 9540 910
rect 9550 900 9990 910
rect 700 890 710 900
rect 3830 890 3840 900
rect 3920 890 3930 900
rect 4050 890 4620 900
rect 4630 890 4850 900
rect 5340 890 5350 900
rect 5380 890 5390 900
rect 5440 890 5450 900
rect 5530 890 5540 900
rect 5610 890 5620 900
rect 6570 890 6810 900
rect 6880 890 7300 900
rect 9170 890 9440 900
rect 9480 890 9540 900
rect 9550 890 9990 900
rect 690 880 700 890
rect 3840 880 3850 890
rect 4050 880 4610 890
rect 4620 880 4850 890
rect 5340 880 5350 890
rect 5380 880 5390 890
rect 5440 880 5450 890
rect 5470 880 5480 890
rect 6570 880 6810 890
rect 6880 880 7290 890
rect 9180 880 9430 890
rect 9480 880 9530 890
rect 9560 880 9990 890
rect 3850 870 3860 880
rect 4050 870 4570 880
rect 4610 870 4860 880
rect 5350 870 5360 880
rect 5390 870 5400 880
rect 6570 870 6820 880
rect 6890 870 7290 880
rect 9180 870 9430 880
rect 9480 870 9520 880
rect 9590 870 9990 880
rect 680 860 690 870
rect 3860 860 3870 870
rect 4050 860 4240 870
rect 4260 860 4560 870
rect 4600 860 4860 870
rect 6570 860 6820 870
rect 6890 860 7290 870
rect 9190 860 9420 870
rect 9470 860 9520 870
rect 9540 860 9550 870
rect 9590 860 9820 870
rect 9830 860 9990 870
rect 2450 850 2470 860
rect 2530 850 2540 860
rect 2550 850 2560 860
rect 4050 850 4240 860
rect 4270 850 4560 860
rect 4590 850 4870 860
rect 6570 850 6830 860
rect 6890 850 7290 860
rect 9190 850 9420 860
rect 9460 850 9800 860
rect 9830 850 9990 860
rect 2430 840 2490 850
rect 2520 840 2570 850
rect 3880 840 3890 850
rect 4050 840 4250 850
rect 4280 840 4570 850
rect 4590 840 4880 850
rect 6580 840 6830 850
rect 6890 840 7290 850
rect 9190 840 9410 850
rect 9460 840 9780 850
rect 9800 840 9850 850
rect 9890 840 9990 850
rect 670 830 680 840
rect 2420 830 2490 840
rect 2540 830 2580 840
rect 4050 830 4250 840
rect 4290 830 4330 840
rect 4340 830 4570 840
rect 4580 830 4880 840
rect 6580 830 6830 840
rect 6890 830 7290 840
rect 9200 830 9410 840
rect 9450 830 9780 840
rect 9800 830 9850 840
rect 9880 830 9990 840
rect 670 820 690 830
rect 2370 820 2380 830
rect 2420 820 2470 830
rect 2480 820 2500 830
rect 2520 820 2570 830
rect 3900 820 3910 830
rect 4050 820 4270 830
rect 4300 820 4320 830
rect 4340 820 4890 830
rect 6580 820 6840 830
rect 6890 820 7280 830
rect 9200 820 9400 830
rect 9450 820 9830 830
rect 9880 820 9910 830
rect 9920 820 9990 830
rect 670 810 680 820
rect 2370 810 2390 820
rect 2410 810 2450 820
rect 2460 810 2470 820
rect 2500 810 2560 820
rect 4040 810 4270 820
rect 4340 810 4890 820
rect 6580 810 6840 820
rect 6890 810 7280 820
rect 9200 810 9290 820
rect 9300 810 9390 820
rect 9440 810 9810 820
rect 9860 810 9880 820
rect 9940 810 9990 820
rect 660 800 670 810
rect 2390 800 2430 810
rect 2470 800 2560 810
rect 4040 800 4280 810
rect 4350 800 4900 810
rect 6580 800 6840 810
rect 6890 800 7280 810
rect 9200 800 9290 810
rect 9320 800 9390 810
rect 9430 800 9880 810
rect 9910 800 9930 810
rect 9950 800 9990 810
rect 660 790 670 800
rect 2360 790 2370 800
rect 2380 790 2420 800
rect 2470 790 2550 800
rect 4030 790 4290 800
rect 4350 790 4900 800
rect 6590 790 6840 800
rect 6890 790 7280 800
rect 9200 790 9290 800
rect 9320 790 9380 800
rect 9430 790 9940 800
rect 9950 790 9990 800
rect 2360 780 2430 790
rect 2470 780 2540 790
rect 4030 780 4300 790
rect 4350 780 4900 790
rect 6590 780 6840 790
rect 6900 780 7280 790
rect 9210 780 9300 790
rect 9330 780 9380 790
rect 9420 780 9990 790
rect 660 770 670 780
rect 2340 770 2430 780
rect 2460 770 2520 780
rect 4030 770 4310 780
rect 4350 770 4910 780
rect 6590 770 6840 780
rect 6900 770 7280 780
rect 9210 770 9240 780
rect 9250 770 9370 780
rect 9420 770 9610 780
rect 9620 770 9840 780
rect 9850 770 9990 780
rect 650 760 670 770
rect 2320 760 2330 770
rect 2340 760 2430 770
rect 2460 760 2500 770
rect 3710 760 3760 770
rect 3800 760 3810 770
rect 4030 760 4320 770
rect 4350 760 4910 770
rect 6590 760 6840 770
rect 6900 760 7280 770
rect 9210 760 9240 770
rect 9260 760 9360 770
rect 9410 760 9460 770
rect 9510 760 9610 770
rect 9630 760 9990 770
rect 650 750 660 760
rect 2310 750 2440 760
rect 2450 750 2480 760
rect 3600 750 3660 760
rect 3710 750 3870 760
rect 4000 750 4020 760
rect 4040 750 4330 760
rect 4350 750 4530 760
rect 4540 750 4800 760
rect 4810 750 4910 760
rect 6590 750 6840 760
rect 6900 750 7280 760
rect 9210 750 9240 760
rect 9250 750 9360 760
rect 9410 750 9460 760
rect 9490 750 9620 760
rect 9630 750 9990 760
rect 640 740 660 750
rect 2290 740 2470 750
rect 3560 740 3890 750
rect 4010 740 4020 750
rect 4060 740 4340 750
rect 4350 740 4530 750
rect 4540 740 4790 750
rect 4810 740 4910 750
rect 6600 740 6840 750
rect 6900 740 7280 750
rect 9230 740 9350 750
rect 9400 740 9450 750
rect 9480 740 9990 750
rect 640 730 660 740
rect 2270 730 2450 740
rect 3520 730 3900 740
rect 4080 730 4110 740
rect 4130 730 4140 740
rect 4160 730 4170 740
rect 4180 730 4520 740
rect 4540 730 4780 740
rect 4810 730 4910 740
rect 6600 730 6840 740
rect 6910 730 7270 740
rect 9220 730 9290 740
rect 9310 730 9350 740
rect 9390 730 9450 740
rect 9460 730 9680 740
rect 9730 730 9990 740
rect 640 720 660 730
rect 2180 720 2220 730
rect 2240 720 2440 730
rect 3490 720 3910 730
rect 4220 720 4770 730
rect 4800 720 4910 730
rect 6610 720 6840 730
rect 6910 720 7270 730
rect 9300 720 9340 730
rect 9390 720 9670 730
rect 9690 720 9990 730
rect 630 710 650 720
rect 2190 710 2200 720
rect 2210 710 2230 720
rect 2240 710 2390 720
rect 2410 710 2420 720
rect 3410 710 3920 720
rect 4230 710 4730 720
rect 4820 710 4920 720
rect 6620 710 6840 720
rect 6920 710 7270 720
rect 9260 710 9340 720
rect 9390 710 9510 720
rect 9520 710 9530 720
rect 9560 710 9990 720
rect 630 700 650 710
rect 2200 700 2380 710
rect 2390 700 2400 710
rect 3390 700 3940 710
rect 4210 700 4710 710
rect 4830 700 4910 710
rect 6620 700 6840 710
rect 6920 700 7260 710
rect 9100 700 9110 710
rect 9220 700 9330 710
rect 9380 700 9990 710
rect 620 690 640 700
rect 2220 690 2320 700
rect 2330 690 2360 700
rect 2370 690 2380 700
rect 3360 690 4040 700
rect 4200 690 4710 700
rect 4840 690 4890 700
rect 6630 690 6850 700
rect 6920 690 7240 700
rect 9210 690 9330 700
rect 9370 690 9990 700
rect 620 680 640 690
rect 2260 680 2300 690
rect 2330 680 2350 690
rect 2360 680 2370 690
rect 3350 680 4050 690
rect 4190 680 4710 690
rect 4850 680 4880 690
rect 6640 680 6850 690
rect 6940 680 7250 690
rect 9220 680 9320 690
rect 9360 680 9680 690
rect 9710 680 9990 690
rect 2250 670 2300 680
rect 2330 670 2340 680
rect 3330 670 4050 680
rect 4180 670 4710 680
rect 4890 670 4920 680
rect 6640 670 6850 680
rect 6940 670 7240 680
rect 9220 670 9310 680
rect 9360 670 9610 680
rect 9630 670 9680 680
rect 9720 670 9990 680
rect 2260 660 2280 670
rect 2290 660 2300 670
rect 2310 660 2330 670
rect 3310 660 4060 670
rect 4170 660 4710 670
rect 4870 660 4920 670
rect 6650 660 6850 670
rect 6940 660 7230 670
rect 9230 660 9310 670
rect 9350 660 9590 670
rect 9640 660 9690 670
rect 9720 660 9990 670
rect 2270 650 2280 660
rect 3300 650 4070 660
rect 4160 650 4560 660
rect 4570 650 4700 660
rect 4860 650 4920 660
rect 6660 650 6850 660
rect 6940 650 7230 660
rect 9220 650 9310 660
rect 9350 650 9590 660
rect 9650 650 9680 660
rect 9730 650 9990 660
rect 3290 640 4080 650
rect 4130 640 4560 650
rect 4570 640 4690 650
rect 4850 640 4930 650
rect 6660 640 6850 650
rect 6950 640 6960 650
rect 6970 640 7220 650
rect 9180 640 9300 650
rect 9340 640 9590 650
rect 9660 640 9670 650
rect 9690 640 9720 650
rect 9740 640 9940 650
rect 9960 640 9990 650
rect 3270 630 4080 640
rect 4120 630 4550 640
rect 4570 630 4680 640
rect 4830 630 4930 640
rect 6680 630 6860 640
rect 6960 630 7210 640
rect 9200 630 9290 640
rect 9340 630 9590 640
rect 9690 630 9910 640
rect 9920 630 9940 640
rect 9960 630 9990 640
rect 3260 620 4050 630
rect 4110 620 4550 630
rect 4570 620 4670 630
rect 4820 620 4930 630
rect 6680 620 6860 630
rect 6960 620 7220 630
rect 9220 620 9290 630
rect 9330 620 9590 630
rect 9610 620 9620 630
rect 9690 620 9940 630
rect 9980 620 9990 630
rect 3240 610 4040 620
rect 4080 610 4550 620
rect 4570 610 4670 620
rect 4800 610 4930 620
rect 6690 610 6860 620
rect 6970 610 7220 620
rect 9230 610 9280 620
rect 9320 610 9620 620
rect 9660 610 9670 620
rect 9690 610 9960 620
rect 9990 610 9990 620
rect 540 600 560 610
rect 3160 600 3170 610
rect 3220 600 4040 610
rect 4080 600 4540 610
rect 4570 600 4670 610
rect 4800 600 4940 610
rect 6700 600 6860 610
rect 6980 600 7210 610
rect 9140 600 9160 610
rect 9170 600 9180 610
rect 9240 600 9280 610
rect 9320 600 9690 610
rect 9710 600 9990 610
rect 460 590 580 600
rect 3140 590 4050 600
rect 4090 590 4530 600
rect 4570 590 4660 600
rect 4790 590 4940 600
rect 6710 590 6870 600
rect 6990 590 7200 600
rect 9120 590 9140 600
rect 9240 590 9270 600
rect 9310 590 9670 600
rect 9730 590 9910 600
rect 9930 590 9980 600
rect 9990 590 9990 600
rect 430 580 600 590
rect 3130 580 4060 590
rect 4090 580 4510 590
rect 4570 580 4660 590
rect 4790 580 4880 590
rect 4890 580 4940 590
rect 6710 580 6870 590
rect 6990 580 7180 590
rect 7190 580 7200 590
rect 9100 580 9120 590
rect 9240 580 9260 590
rect 9310 580 9620 590
rect 9640 580 9670 590
rect 9700 580 9990 590
rect 390 570 590 580
rect 3120 570 4070 580
rect 4090 570 4370 580
rect 4390 570 4460 580
rect 4570 570 4650 580
rect 4800 570 4870 580
rect 4890 570 4940 580
rect 6710 570 6870 580
rect 7020 570 7160 580
rect 7190 570 7200 580
rect 9240 570 9260 580
rect 9300 570 9630 580
rect 9660 570 9960 580
rect 9970 570 9990 580
rect 370 560 600 570
rect 3110 560 4350 570
rect 4560 560 4640 570
rect 4800 560 4860 570
rect 4900 560 4940 570
rect 6720 560 6870 570
rect 7030 560 7160 570
rect 9240 560 9250 570
rect 9300 560 9650 570
rect 9660 560 9780 570
rect 9790 560 9930 570
rect 9940 560 9950 570
rect 9960 560 9990 570
rect 360 550 550 560
rect 560 550 580 560
rect 1400 550 1440 560
rect 3030 550 3080 560
rect 3100 550 4330 560
rect 4570 550 4630 560
rect 4810 550 4840 560
rect 4900 550 4950 560
rect 6730 550 6880 560
rect 7030 550 7140 560
rect 9230 550 9250 560
rect 9290 550 9940 560
rect 9960 550 9990 560
rect 360 540 540 550
rect 1390 540 1440 550
rect 3010 540 4250 550
rect 4580 540 4600 550
rect 4800 540 4840 550
rect 4900 540 4950 550
rect 6740 540 6880 550
rect 7030 540 7130 550
rect 9220 540 9240 550
rect 9290 540 9960 550
rect 350 530 530 540
rect 1310 530 1330 540
rect 1370 530 1440 540
rect 2990 530 4240 540
rect 4790 530 4850 540
rect 4900 530 4950 540
rect 6750 530 6880 540
rect 7030 530 7120 540
rect 9220 530 9230 540
rect 9280 530 9960 540
rect 370 520 510 530
rect 1260 520 1460 530
rect 2980 520 4220 530
rect 4790 520 4860 530
rect 4900 520 4950 530
rect 6750 520 6880 530
rect 7080 520 7130 530
rect 9270 520 9940 530
rect 370 510 490 520
rect 1260 510 1490 520
rect 2970 510 4220 520
rect 4790 510 4870 520
rect 4900 510 4950 520
rect 6750 510 6890 520
rect 7110 510 7120 520
rect 9270 510 9920 520
rect 380 500 470 510
rect 1250 500 1490 510
rect 2940 500 4210 510
rect 4790 500 4870 510
rect 4900 500 4960 510
rect 6770 500 6880 510
rect 9260 500 9910 510
rect 390 490 460 500
rect 1200 490 1480 500
rect 2900 490 4200 500
rect 4790 490 4860 500
rect 4900 490 4960 500
rect 6760 490 6890 500
rect 9260 490 9860 500
rect 9890 490 9900 500
rect 9950 490 9980 500
rect 400 480 440 490
rect 1180 480 1480 490
rect 2870 480 4190 490
rect 4800 480 4860 490
rect 4900 480 4960 490
rect 6770 480 6900 490
rect 9250 480 9860 490
rect 9940 480 9990 490
rect 1170 470 1480 480
rect 1520 470 1530 480
rect 2840 470 4180 480
rect 4790 470 4860 480
rect 4910 470 4960 480
rect 6790 470 6810 480
rect 6830 470 6890 480
rect 9190 470 9200 480
rect 9250 470 9850 480
rect 9940 470 9990 480
rect 1160 460 1480 470
rect 1510 460 1540 470
rect 2800 460 4180 470
rect 4790 460 4870 470
rect 4910 460 4960 470
rect 6800 460 6810 470
rect 6840 460 6900 470
rect 9180 460 9190 470
rect 9250 460 9300 470
rect 9320 460 9850 470
rect 9880 460 9910 470
rect 9930 460 9990 470
rect 160 450 240 460
rect 1150 450 1470 460
rect 1510 450 1540 460
rect 2080 450 2190 460
rect 2740 450 4170 460
rect 4780 450 4880 460
rect 4920 450 4960 460
rect 6870 450 6900 460
rect 9170 450 9190 460
rect 9240 450 9290 460
rect 9320 450 9370 460
rect 9410 450 9860 460
rect 9880 450 9990 460
rect 140 440 270 450
rect 1140 440 1470 450
rect 1510 440 1540 450
rect 2030 440 2250 450
rect 2690 440 4170 450
rect 4780 440 4880 450
rect 4920 440 4960 450
rect 6870 440 6890 450
rect 9170 440 9180 450
rect 9230 440 9290 450
rect 9340 440 9860 450
rect 9880 440 9990 450
rect 120 430 280 440
rect 1130 430 1470 440
rect 1510 430 1550 440
rect 1980 430 2280 440
rect 2650 430 4160 440
rect 4770 430 4890 440
rect 4910 430 4970 440
rect 6860 430 6880 440
rect 9160 430 9180 440
rect 9220 430 9280 440
rect 9350 430 9990 440
rect 110 420 280 430
rect 1130 420 1470 430
rect 1500 420 1690 430
rect 1860 420 2310 430
rect 2600 420 4160 430
rect 4770 420 4900 430
rect 4910 420 4970 430
rect 9160 420 9170 430
rect 9220 420 9290 430
rect 9380 420 9990 430
rect 100 410 290 420
rect 1120 410 1470 420
rect 1500 410 2340 420
rect 2530 410 4150 420
rect 4760 410 4970 420
rect 9160 410 9170 420
rect 9210 410 9290 420
rect 9300 410 9320 420
rect 9400 410 9990 420
rect 100 400 300 410
rect 1110 400 1470 410
rect 1500 400 2420 410
rect 2460 400 4150 410
rect 4760 400 4970 410
rect 9140 400 9160 410
rect 9200 400 9270 410
rect 9290 400 9310 410
rect 9400 400 9980 410
rect 9990 400 9990 410
rect 90 390 300 400
rect 1110 390 1470 400
rect 1500 390 4140 400
rect 4760 390 4970 400
rect 9140 390 9150 400
rect 9200 390 9260 400
rect 9410 390 9990 400
rect 80 380 300 390
rect 1100 380 1230 390
rect 1250 380 1470 390
rect 1490 380 4140 390
rect 4750 380 4970 390
rect 9130 380 9150 390
rect 9200 380 9250 390
rect 9420 380 9990 390
rect 70 370 300 380
rect 1090 370 1230 380
rect 1260 370 1470 380
rect 1490 370 4140 380
rect 4760 370 4920 380
rect 4930 370 4970 380
rect 9120 370 9140 380
rect 9190 370 9250 380
rect 9430 370 9700 380
rect 9710 370 9990 380
rect 70 360 290 370
rect 1080 360 1220 370
rect 1250 360 1470 370
rect 1480 360 4140 370
rect 4760 360 4910 370
rect 4940 360 4970 370
rect 9120 360 9140 370
rect 9180 360 9240 370
rect 9430 360 9970 370
rect 9990 360 9990 370
rect 60 350 290 360
rect 1080 350 4130 360
rect 4760 350 4900 360
rect 4960 350 4970 360
rect 9110 350 9130 360
rect 9180 350 9230 360
rect 9440 350 9970 360
rect 9990 350 9990 360
rect 60 340 280 350
rect 1070 340 4120 350
rect 4770 340 4900 350
rect 9110 340 9130 350
rect 9170 340 9220 350
rect 9430 340 9940 350
rect 50 330 100 340
rect 110 330 270 340
rect 1060 330 4110 340
rect 4770 330 4820 340
rect 4830 330 4850 340
rect 4860 330 4880 340
rect 4960 330 4970 340
rect 9100 330 9120 340
rect 9160 330 9220 340
rect 9420 330 9490 340
rect 9510 330 9980 340
rect 9990 330 9990 340
rect 50 320 100 330
rect 120 320 260 330
rect 1050 320 4090 330
rect 4800 320 4810 330
rect 4960 320 4970 330
rect 9090 320 9120 330
rect 9160 320 9210 330
rect 9420 320 9490 330
rect 9530 320 9990 330
rect 40 310 70 320
rect 130 310 240 320
rect 1050 310 4080 320
rect 4950 310 4970 320
rect 9090 310 9110 320
rect 9160 310 9210 320
rect 9420 310 9990 320
rect 40 300 70 310
rect 140 300 230 310
rect 1040 300 1270 310
rect 1290 300 4070 310
rect 4960 300 4970 310
rect 9080 300 9110 310
rect 9150 300 9210 310
rect 9430 300 9720 310
rect 9740 300 9750 310
rect 9760 300 9990 310
rect 30 290 70 300
rect 150 290 210 300
rect 510 290 550 300
rect 1040 290 1260 300
rect 1310 290 4070 300
rect 4950 290 4960 300
rect 4970 290 4980 300
rect 9070 290 9100 300
rect 9140 290 9210 300
rect 9440 290 9500 300
rect 9520 290 9560 300
rect 9580 290 9690 300
rect 9760 290 9810 300
rect 9820 290 9990 300
rect 30 280 60 290
rect 520 280 560 290
rect 1040 280 1250 290
rect 1310 280 4070 290
rect 4950 280 4980 290
rect 9070 280 9090 290
rect 9130 280 9200 290
rect 9450 280 9500 290
rect 9520 280 9550 290
rect 9580 280 9620 290
rect 9640 280 9810 290
rect 9820 280 9990 290
rect 30 270 50 280
rect 520 270 560 280
rect 1040 270 1240 280
rect 1300 270 4070 280
rect 4220 270 4230 280
rect 4950 270 4980 280
rect 9060 270 9090 280
rect 9130 270 9190 280
rect 9470 270 9500 280
rect 9530 270 9560 280
rect 9590 270 9810 280
rect 9820 270 9990 280
rect 520 260 550 270
rect 1030 260 1230 270
rect 1290 260 4080 270
rect 4940 260 4990 270
rect 9060 260 9080 270
rect 9120 260 9190 270
rect 9310 260 9330 270
rect 9480 260 9520 270
rect 9540 260 9550 270
rect 9580 260 9790 270
rect 9800 260 9820 270
rect 9840 260 9980 270
rect 520 250 550 260
rect 1030 250 1230 260
rect 1280 250 4090 260
rect 4940 250 4990 260
rect 9050 250 9080 260
rect 9120 250 9190 260
rect 9300 250 9340 260
rect 9390 250 9410 260
rect 9440 250 9460 260
rect 9480 250 9530 260
rect 9550 250 9590 260
rect 9600 250 9820 260
rect 9850 250 9990 260
rect 520 240 550 250
rect 1030 240 1220 250
rect 1270 240 4090 250
rect 4950 240 4990 250
rect 9040 240 9070 250
rect 9110 240 9170 250
rect 9300 240 9330 250
rect 9390 240 9400 250
rect 9450 240 9490 250
rect 9500 240 9590 250
rect 9610 240 9790 250
rect 9820 240 9830 250
rect 9850 240 9990 250
rect 530 230 540 240
rect 1030 230 1220 240
rect 1230 230 4100 240
rect 4950 230 4990 240
rect 9040 230 9070 240
rect 9110 230 9160 240
rect 9400 230 9420 240
rect 9460 230 9470 240
rect 9510 230 9780 240
rect 9850 230 9990 240
rect 530 220 540 230
rect 1030 220 4100 230
rect 4940 220 4990 230
rect 8880 220 8890 230
rect 9030 220 9060 230
rect 9100 220 9160 230
rect 9410 220 9430 230
rect 9520 220 9780 230
rect 9860 220 9990 230
rect 520 210 540 220
rect 1030 210 4110 220
rect 4940 210 5000 220
rect 8880 210 8890 220
rect 9030 210 9060 220
rect 9100 210 9160 220
rect 9320 210 9350 220
rect 9410 210 9780 220
rect 9850 210 9930 220
rect 9960 210 9990 220
rect 1020 200 4120 210
rect 4920 200 4930 210
rect 4950 200 5000 210
rect 8880 200 8910 210
rect 9020 200 9050 210
rect 9090 200 9150 210
rect 9160 200 9180 210
rect 9310 200 9680 210
rect 9690 200 9780 210
rect 9850 200 9940 210
rect 9970 200 9990 210
rect 1020 190 4130 200
rect 4930 190 5000 200
rect 8870 190 8910 200
rect 9010 190 9040 200
rect 9080 190 9140 200
rect 9300 190 9680 200
rect 9700 190 9740 200
rect 9850 190 9920 200
rect 9990 190 9990 200
rect 1020 180 4140 190
rect 4930 180 5000 190
rect 8860 180 8880 190
rect 8890 180 8900 190
rect 9010 180 9040 190
rect 9080 180 9130 190
rect 9310 180 9690 190
rect 9700 180 9730 190
rect 9870 180 9890 190
rect 1020 170 4150 180
rect 4940 170 5000 180
rect 9000 170 9030 180
rect 9080 170 9130 180
rect 9330 170 9710 180
rect 9960 170 9970 180
rect 1020 160 4160 170
rect 4940 160 5000 170
rect 9010 160 9030 170
rect 9080 160 9130 170
rect 9160 160 9180 170
rect 9340 160 9550 170
rect 9560 160 9690 170
rect 9950 160 9970 170
rect 1010 150 4170 160
rect 4980 150 5010 160
rect 8840 150 8870 160
rect 9080 150 9130 160
rect 9340 150 9550 160
rect 9570 150 9600 160
rect 9610 150 9700 160
rect 1010 140 4180 150
rect 4980 140 5010 150
rect 8840 140 8900 150
rect 9090 140 9130 150
rect 9350 140 9560 150
rect 9630 140 9650 150
rect 9660 140 9710 150
rect 9990 140 9990 150
rect 1010 130 4200 140
rect 4980 130 5010 140
rect 8840 130 8920 140
rect 9110 130 9140 140
rect 9350 130 9600 140
rect 9620 130 9710 140
rect 9980 130 9990 140
rect 1020 120 4210 130
rect 4980 120 5020 130
rect 8830 120 8930 130
rect 9110 120 9150 130
rect 9350 120 9370 130
rect 9380 120 9710 130
rect 9990 120 9990 130
rect 1020 110 4220 120
rect 4970 110 5020 120
rect 8830 110 8930 120
rect 9100 110 9140 120
rect 9420 110 9470 120
rect 9490 110 9730 120
rect 1020 100 4230 110
rect 4970 100 5030 110
rect 8840 100 8930 110
rect 9100 100 9140 110
rect 9430 100 9480 110
rect 9500 100 9570 110
rect 9590 100 9640 110
rect 9650 100 9730 110
rect 9870 100 9880 110
rect 9920 100 9940 110
rect 1020 90 4240 100
rect 4970 90 5030 100
rect 8810 90 8940 100
rect 9090 90 9140 100
rect 9440 90 9560 100
rect 9590 90 9730 100
rect 9920 90 9950 100
rect 1030 80 4250 90
rect 4970 80 5030 90
rect 8790 80 8930 90
rect 9090 80 9140 90
rect 9450 80 9560 90
rect 9600 80 9730 90
rect 9910 80 9950 90
rect 0 70 20 80
rect 1030 70 4270 80
rect 4980 70 5040 80
rect 8780 70 8900 80
rect 9090 70 9140 80
rect 9460 70 9550 80
rect 9610 70 9660 80
rect 9700 70 9740 80
rect 9930 70 9940 80
rect 0 60 20 70
rect 1030 60 4280 70
rect 4980 60 5040 70
rect 8780 60 8900 70
rect 8920 60 8930 70
rect 9010 60 9030 70
rect 9060 60 9070 70
rect 9090 60 9150 70
rect 9480 60 9540 70
rect 9560 60 9580 70
rect 9610 60 9660 70
rect 9720 60 9740 70
rect 9930 60 9950 70
rect 0 50 20 60
rect 1030 50 4300 60
rect 4980 50 5040 60
rect 8770 50 8900 60
rect 8940 50 8950 60
rect 9010 50 9070 60
rect 9100 50 9160 60
rect 9500 50 9530 60
rect 9570 50 9580 60
rect 9640 50 9660 60
rect 9720 50 9740 60
rect 9940 50 9950 60
rect 0 40 20 50
rect 1030 40 4310 50
rect 4980 40 5050 50
rect 8760 40 8920 50
rect 9020 40 9080 50
rect 9100 40 9160 50
rect 9640 40 9670 50
rect 9720 40 9740 50
rect 9940 40 9970 50
rect 0 30 20 40
rect 1020 30 4330 40
rect 4980 30 5050 40
rect 8750 30 8930 40
rect 9030 30 9080 40
rect 9100 30 9170 40
rect 9610 30 9620 40
rect 9630 30 9670 40
rect 9720 30 9770 40
rect 9940 30 9980 40
rect 0 20 20 30
rect 1020 20 1290 30
rect 1310 20 4340 30
rect 4980 20 5050 30
rect 8730 20 8920 30
rect 9040 20 9090 30
rect 9110 20 9160 30
rect 9530 20 9580 30
rect 9630 20 9660 30
rect 9720 20 9770 30
rect 9940 20 9990 30
rect 0 10 10 20
rect 1020 10 1280 20
rect 1320 10 4350 20
rect 4980 10 5050 20
rect 8580 10 8610 20
rect 8730 10 8910 20
rect 9040 10 9090 20
rect 9120 10 9170 20
rect 9490 10 9590 20
rect 9640 10 9660 20
rect 9720 10 9780 20
rect 9950 10 9960 20
rect 9980 10 9990 20
rect 1020 0 1280 10
rect 1320 0 4370 10
rect 4980 0 5060 10
rect 8610 0 8670 10
rect 8720 0 8790 10
rect 8800 0 8900 10
rect 9030 0 9090 10
rect 9120 0 9180 10
rect 9480 0 9600 10
rect 9740 0 9780 10
rect 9940 0 9980 10
rect 9990 0 9990 10
<< end >>
