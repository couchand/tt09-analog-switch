magic
tech sky130A
timestamp 1730992266
<< locali >>
rect 2280 7490 3320 7500
rect 3560 7490 3640 7500
rect 2280 7480 3320 7490
rect 3560 7480 3640 7490
rect 2280 7470 3320 7480
rect 3560 7470 3640 7480
rect 2280 7460 3320 7470
rect 3560 7460 3640 7470
rect 2200 7450 3320 7460
rect 3600 7450 3640 7460
rect 9800 7450 9920 7460
rect 2200 7440 3320 7450
rect 3600 7440 3640 7450
rect 9800 7440 9920 7450
rect 2200 7430 3320 7440
rect 3600 7430 3640 7440
rect 9800 7430 9920 7440
rect 2200 7420 3320 7430
rect 3600 7420 3640 7430
rect 9800 7420 9920 7430
rect 2160 7410 3320 7420
rect 9760 7410 9840 7420
rect 2160 7400 3320 7410
rect 9760 7400 9840 7410
rect 2160 7390 3320 7400
rect 9760 7390 9840 7400
rect 2160 7380 3320 7390
rect 9760 7380 9840 7390
rect 2120 7370 3320 7380
rect 2120 7360 3320 7370
rect 2120 7350 3320 7360
rect 2120 7340 3320 7350
rect 2080 7330 3320 7340
rect 2080 7320 3320 7330
rect 2080 7310 3320 7320
rect 2080 7300 3320 7310
rect 2080 7290 2520 7300
rect 2560 7290 3320 7300
rect 2080 7280 2520 7290
rect 2560 7280 3320 7290
rect 2080 7270 2520 7280
rect 2560 7270 3320 7280
rect 2080 7260 2520 7270
rect 2560 7260 3320 7270
rect 2040 7250 2440 7260
rect 2560 7250 3320 7260
rect 2040 7240 2440 7250
rect 2560 7240 3320 7250
rect 2040 7230 2440 7240
rect 2560 7230 3320 7240
rect 2040 7220 2440 7230
rect 2560 7220 3320 7230
rect 2040 7210 2120 7220
rect 2280 7210 2400 7220
rect 2440 7210 3320 7220
rect 2040 7200 2120 7210
rect 2280 7200 2400 7210
rect 2440 7200 3320 7210
rect 2040 7190 2120 7200
rect 2280 7190 2400 7200
rect 2440 7190 3320 7200
rect 2040 7180 2120 7190
rect 2280 7180 2400 7190
rect 2440 7180 3320 7190
rect 2000 7170 2080 7180
rect 2320 7170 3320 7180
rect 2000 7160 2080 7170
rect 2320 7160 3320 7170
rect 2000 7150 2080 7160
rect 2320 7150 3320 7160
rect 2000 7140 2080 7150
rect 2320 7140 3320 7150
rect 2000 7130 2040 7140
rect 2200 7130 3400 7140
rect 9880 7130 9920 7140
rect 2000 7120 2040 7130
rect 2200 7120 3400 7130
rect 9880 7120 9920 7130
rect 2000 7110 2040 7120
rect 2200 7110 3400 7120
rect 9880 7110 9920 7120
rect 2000 7100 2040 7110
rect 2200 7100 3400 7110
rect 9880 7100 9920 7110
rect 2160 7090 3400 7100
rect 9840 7090 9960 7100
rect 2160 7080 3400 7090
rect 9840 7080 9960 7090
rect 2160 7070 3400 7080
rect 9840 7070 9960 7080
rect 2160 7060 3400 7070
rect 9840 7060 9960 7070
rect 2120 7050 2200 7060
rect 3080 7050 3440 7060
rect 9800 7050 9920 7060
rect 2120 7040 2200 7050
rect 3080 7040 3440 7050
rect 9800 7040 9920 7050
rect 2120 7030 2200 7040
rect 3080 7030 3440 7040
rect 9800 7030 9920 7040
rect 2120 7020 2200 7030
rect 3080 7020 3440 7030
rect 9800 7020 9920 7030
rect 2040 7010 2160 7020
rect 3240 7010 3480 7020
rect 9720 7010 9760 7020
rect 2040 7000 2160 7010
rect 3240 7000 3480 7010
rect 9720 7000 9760 7010
rect 2040 6990 2160 7000
rect 3240 6990 3480 7000
rect 9720 6990 9760 7000
rect 2040 6980 2160 6990
rect 3240 6980 3480 6990
rect 9720 6980 9760 6990
rect 2000 6970 2160 6980
rect 3360 6970 3520 6980
rect 9680 6970 9720 6980
rect 9880 6970 9990 6980
rect 2000 6960 2160 6970
rect 3360 6960 3520 6970
rect 9680 6960 9720 6970
rect 9880 6960 9990 6970
rect 2000 6950 2160 6960
rect 3360 6950 3520 6960
rect 9680 6950 9720 6960
rect 9880 6950 9990 6960
rect 2000 6940 2160 6950
rect 3360 6940 3520 6950
rect 9680 6940 9720 6950
rect 9880 6940 9990 6950
rect 1960 6930 2200 6940
rect 3480 6930 3560 6940
rect 9840 6930 9990 6940
rect 1960 6920 2200 6930
rect 3480 6920 3560 6930
rect 9840 6920 9990 6930
rect 1960 6910 2200 6920
rect 3480 6910 3560 6920
rect 9840 6910 9990 6920
rect 1960 6900 2200 6910
rect 3480 6900 3560 6910
rect 9840 6900 9990 6910
rect 1920 6890 2240 6900
rect 3560 6890 3640 6900
rect 9880 6890 9990 6900
rect 1920 6880 2240 6890
rect 3560 6880 3640 6890
rect 9880 6880 9990 6890
rect 1920 6870 2240 6880
rect 3560 6870 3640 6880
rect 9880 6870 9990 6880
rect 1920 6860 2240 6870
rect 3560 6860 3640 6870
rect 9880 6860 9990 6870
rect 1920 6850 2280 6860
rect 3600 6850 3680 6860
rect 9880 6850 9920 6860
rect 1920 6840 2280 6850
rect 3600 6840 3680 6850
rect 9880 6840 9920 6850
rect 1920 6830 2280 6840
rect 3600 6830 3680 6840
rect 9880 6830 9920 6840
rect 1920 6820 2280 6830
rect 3600 6820 3680 6830
rect 9880 6820 9920 6830
rect 1920 6810 1960 6820
rect 2040 6810 2280 6820
rect 3680 6810 3720 6820
rect 9880 6810 9920 6820
rect 1920 6800 1960 6810
rect 2040 6800 2280 6810
rect 3680 6800 3720 6810
rect 9880 6800 9920 6810
rect 1920 6790 1960 6800
rect 2040 6790 2280 6800
rect 3680 6790 3720 6800
rect 9880 6790 9920 6800
rect 1920 6780 1960 6790
rect 2040 6780 2280 6790
rect 3680 6780 3720 6790
rect 9880 6780 9920 6790
rect 2040 6770 2240 6780
rect 2440 6770 2520 6780
rect 2600 6770 2640 6780
rect 3760 6770 3800 6780
rect 9840 6770 9960 6780
rect 2040 6760 2240 6770
rect 2440 6760 2520 6770
rect 2600 6760 2640 6770
rect 3760 6760 3800 6770
rect 9840 6760 9960 6770
rect 2040 6750 2240 6760
rect 2440 6750 2520 6760
rect 2600 6750 2640 6760
rect 3760 6750 3800 6760
rect 9840 6750 9960 6760
rect 2040 6740 2240 6750
rect 2440 6740 2520 6750
rect 2600 6740 2640 6750
rect 3760 6740 3800 6750
rect 9840 6740 9960 6750
rect 2000 6730 2200 6740
rect 2560 6730 3000 6740
rect 3800 6730 3840 6740
rect 9840 6730 9990 6740
rect 2000 6720 2200 6730
rect 2560 6720 3000 6730
rect 3800 6720 3840 6730
rect 9840 6720 9990 6730
rect 2000 6710 2200 6720
rect 2560 6710 3000 6720
rect 3800 6710 3840 6720
rect 9840 6710 9990 6720
rect 2000 6700 2200 6710
rect 2560 6700 3000 6710
rect 3800 6700 3840 6710
rect 9840 6700 9990 6710
rect 1960 6690 2200 6700
rect 2640 6690 3280 6700
rect 3840 6690 3880 6700
rect 9840 6690 9880 6700
rect 1960 6680 2200 6690
rect 2640 6680 3280 6690
rect 3840 6680 3880 6690
rect 9840 6680 9880 6690
rect 1960 6670 2200 6680
rect 2640 6670 3280 6680
rect 3840 6670 3880 6680
rect 9840 6670 9880 6680
rect 1960 6660 2200 6670
rect 2640 6660 3280 6670
rect 3840 6660 3880 6670
rect 9840 6660 9880 6670
rect 1920 6650 2200 6660
rect 2680 6650 3480 6660
rect 3880 6650 3920 6660
rect 1920 6640 2200 6650
rect 2680 6640 3480 6650
rect 3880 6640 3920 6650
rect 1920 6630 2200 6640
rect 2680 6630 3480 6640
rect 3880 6630 3920 6640
rect 1920 6620 2200 6630
rect 2680 6620 3480 6630
rect 3880 6620 3920 6630
rect 1800 6610 2120 6620
rect 2680 6610 3600 6620
rect 1800 6600 2120 6610
rect 2680 6600 3600 6610
rect 1800 6590 2120 6600
rect 2680 6590 3600 6600
rect 1800 6580 2120 6590
rect 2680 6580 3600 6590
rect 1840 6570 2000 6580
rect 2680 6570 3720 6580
rect 1840 6560 2000 6570
rect 2680 6560 3720 6570
rect 1840 6550 2000 6560
rect 2680 6550 3720 6560
rect 1840 6540 2000 6550
rect 2680 6540 3720 6550
rect 1520 6530 1560 6540
rect 1640 6530 1720 6540
rect 1880 6530 2040 6540
rect 2640 6530 3800 6540
rect 1520 6520 1560 6530
rect 1640 6520 1720 6530
rect 1880 6520 2040 6530
rect 2640 6520 3800 6530
rect 1520 6510 1560 6520
rect 1640 6510 1720 6520
rect 1880 6510 2040 6520
rect 2640 6510 3800 6520
rect 1520 6500 1560 6510
rect 1640 6500 1720 6510
rect 1880 6500 2040 6510
rect 2640 6500 3800 6510
rect 1400 6490 1520 6500
rect 1600 6490 1640 6500
rect 1960 6490 2080 6500
rect 2600 6490 3880 6500
rect 1400 6480 1520 6490
rect 1600 6480 1640 6490
rect 1960 6480 2080 6490
rect 2600 6480 3880 6490
rect 1400 6470 1520 6480
rect 1600 6470 1640 6480
rect 1960 6470 2080 6480
rect 2600 6470 3880 6480
rect 1400 6460 1520 6470
rect 1600 6460 1640 6470
rect 1960 6460 2080 6470
rect 2600 6460 3880 6470
rect 1400 6450 1440 6460
rect 1480 6450 1560 6460
rect 2400 6450 2480 6460
rect 2560 6450 3920 6460
rect 9840 6450 9920 6460
rect 1400 6440 1440 6450
rect 1480 6440 1560 6450
rect 2400 6440 2480 6450
rect 2560 6440 3920 6450
rect 9840 6440 9920 6450
rect 1400 6430 1440 6440
rect 1480 6430 1560 6440
rect 2400 6430 2480 6440
rect 2560 6430 3920 6440
rect 9840 6430 9920 6440
rect 1400 6420 1440 6430
rect 1480 6420 1560 6430
rect 2400 6420 2480 6430
rect 2560 6420 3920 6430
rect 9840 6420 9920 6430
rect 1480 6410 1560 6420
rect 2400 6410 4000 6420
rect 9800 6410 9920 6420
rect 1480 6400 1560 6410
rect 2400 6400 4000 6410
rect 9800 6400 9920 6410
rect 1480 6390 1560 6400
rect 2400 6390 4000 6400
rect 9800 6390 9920 6400
rect 1480 6380 1560 6390
rect 2400 6380 4000 6390
rect 9800 6380 9920 6390
rect 1480 6370 1560 6380
rect 1760 6370 1800 6380
rect 2480 6370 4040 6380
rect 9880 6370 9920 6380
rect 1480 6360 1560 6370
rect 1760 6360 1800 6370
rect 2480 6360 4040 6370
rect 9880 6360 9920 6370
rect 1480 6350 1560 6360
rect 1760 6350 1800 6360
rect 2480 6350 4040 6360
rect 9880 6350 9920 6360
rect 1480 6340 1560 6350
rect 1760 6340 1800 6350
rect 2480 6340 4040 6350
rect 9880 6340 9920 6350
rect 1440 6330 1560 6340
rect 1720 6330 1800 6340
rect 2480 6330 4120 6340
rect 9720 6330 9760 6340
rect 9840 6330 9920 6340
rect 1440 6320 1560 6330
rect 1720 6320 1800 6330
rect 2480 6320 4120 6330
rect 9720 6320 9760 6330
rect 9840 6320 9920 6330
rect 1440 6310 1560 6320
rect 1720 6310 1800 6320
rect 2480 6310 4120 6320
rect 9720 6310 9760 6320
rect 9840 6310 9920 6320
rect 1440 6300 1560 6310
rect 1720 6300 1800 6310
rect 2480 6300 4120 6310
rect 9720 6300 9760 6310
rect 9840 6300 9920 6310
rect 1440 6290 1520 6300
rect 1720 6290 1760 6300
rect 2480 6290 4160 6300
rect 5440 6290 5480 6300
rect 9680 6290 9800 6300
rect 1440 6280 1520 6290
rect 1720 6280 1760 6290
rect 2480 6280 4160 6290
rect 5440 6280 5480 6290
rect 9680 6280 9800 6290
rect 1440 6270 1520 6280
rect 1720 6270 1760 6280
rect 2480 6270 4160 6280
rect 5440 6270 5480 6280
rect 9680 6270 9800 6280
rect 1440 6260 1520 6270
rect 1720 6260 1760 6270
rect 2480 6260 4160 6270
rect 5440 6260 5480 6270
rect 9680 6260 9800 6270
rect 1440 6250 1560 6260
rect 1680 6250 1720 6260
rect 2480 6250 4200 6260
rect 5400 6250 5480 6260
rect 9680 6250 9800 6260
rect 1440 6240 1560 6250
rect 1680 6240 1720 6250
rect 2480 6240 4200 6250
rect 5400 6240 5480 6250
rect 9680 6240 9800 6250
rect 1440 6230 1560 6240
rect 1680 6230 1720 6240
rect 2480 6230 4200 6240
rect 5400 6230 5480 6240
rect 9680 6230 9800 6240
rect 1440 6220 1560 6230
rect 1680 6220 1720 6230
rect 2480 6220 4200 6230
rect 5400 6220 5480 6230
rect 9680 6220 9800 6230
rect 1440 6210 1560 6220
rect 2440 6210 4240 6220
rect 5360 6210 5440 6220
rect 9440 6210 9600 6220
rect 9720 6210 9760 6220
rect 1440 6200 1560 6210
rect 2440 6200 4240 6210
rect 5360 6200 5440 6210
rect 9440 6200 9600 6210
rect 9720 6200 9760 6210
rect 1440 6190 1560 6200
rect 2440 6190 4240 6200
rect 5360 6190 5440 6200
rect 9440 6190 9600 6200
rect 9720 6190 9760 6200
rect 1440 6180 1560 6190
rect 2440 6180 4240 6190
rect 5360 6180 5440 6190
rect 9440 6180 9600 6190
rect 9720 6180 9760 6190
rect 1440 6170 1600 6180
rect 2440 6170 4240 6180
rect 5320 6170 5400 6180
rect 9480 6170 9600 6180
rect 9720 6170 9800 6180
rect 1440 6160 1600 6170
rect 2440 6160 4240 6170
rect 5320 6160 5400 6170
rect 9480 6160 9600 6170
rect 9720 6160 9800 6170
rect 1440 6150 1600 6160
rect 2440 6150 4240 6160
rect 5320 6150 5400 6160
rect 9480 6150 9600 6160
rect 9720 6150 9800 6160
rect 1440 6140 1600 6150
rect 2440 6140 4240 6150
rect 5320 6140 5400 6150
rect 9480 6140 9600 6150
rect 9720 6140 9800 6150
rect 1440 6130 1600 6140
rect 2440 6130 3920 6140
rect 3960 6130 4280 6140
rect 5320 6130 5360 6140
rect 9280 6130 9320 6140
rect 9480 6130 9640 6140
rect 9720 6130 9800 6140
rect 1440 6120 1600 6130
rect 2440 6120 3920 6130
rect 3960 6120 4280 6130
rect 5320 6120 5360 6130
rect 9280 6120 9320 6130
rect 9480 6120 9640 6130
rect 9720 6120 9800 6130
rect 1440 6110 1600 6120
rect 2440 6110 3920 6120
rect 3960 6110 4280 6120
rect 5320 6110 5360 6120
rect 9280 6110 9320 6120
rect 9480 6110 9640 6120
rect 9720 6110 9800 6120
rect 1440 6100 1600 6110
rect 2440 6100 3920 6110
rect 3960 6100 4280 6110
rect 5320 6100 5360 6110
rect 9280 6100 9320 6110
rect 9480 6100 9640 6110
rect 9720 6100 9800 6110
rect 1440 6090 1600 6100
rect 2480 6090 3760 6100
rect 4000 6090 4280 6100
rect 5280 6090 5360 6100
rect 9280 6090 9320 6100
rect 9520 6090 9640 6100
rect 9720 6090 9840 6100
rect 1440 6080 1600 6090
rect 2480 6080 3760 6090
rect 4000 6080 4280 6090
rect 5280 6080 5360 6090
rect 9280 6080 9320 6090
rect 9520 6080 9640 6090
rect 9720 6080 9840 6090
rect 1440 6070 1600 6080
rect 2480 6070 3760 6080
rect 4000 6070 4280 6080
rect 5280 6070 5360 6080
rect 9280 6070 9320 6080
rect 9520 6070 9640 6080
rect 9720 6070 9840 6080
rect 1440 6060 1600 6070
rect 2480 6060 3760 6070
rect 4000 6060 4280 6070
rect 5280 6060 5360 6070
rect 9280 6060 9320 6070
rect 9520 6060 9640 6070
rect 9720 6060 9840 6070
rect 1360 6050 1600 6060
rect 2480 6050 3200 6060
rect 3280 6050 3760 6060
rect 4040 6050 4320 6060
rect 5240 6050 5360 6060
rect 9520 6050 9640 6060
rect 9720 6050 9840 6060
rect 1360 6040 1600 6050
rect 2480 6040 3200 6050
rect 3280 6040 3760 6050
rect 4040 6040 4320 6050
rect 5240 6040 5360 6050
rect 9520 6040 9640 6050
rect 9720 6040 9840 6050
rect 1360 6030 1600 6040
rect 2480 6030 3200 6040
rect 3280 6030 3760 6040
rect 4040 6030 4320 6040
rect 5240 6030 5360 6040
rect 9520 6030 9640 6040
rect 9720 6030 9840 6040
rect 1360 6020 1600 6030
rect 2480 6020 3200 6030
rect 3280 6020 3760 6030
rect 4040 6020 4320 6030
rect 5240 6020 5360 6030
rect 9520 6020 9640 6030
rect 9720 6020 9840 6030
rect 1360 6010 1600 6020
rect 2520 6010 3160 6020
rect 3280 6010 3760 6020
rect 4080 6010 4320 6020
rect 5240 6010 5320 6020
rect 9480 6010 9640 6020
rect 9720 6010 9840 6020
rect 1360 6000 1600 6010
rect 2520 6000 3160 6010
rect 3280 6000 3760 6010
rect 4080 6000 4320 6010
rect 5240 6000 5320 6010
rect 9480 6000 9640 6010
rect 9720 6000 9840 6010
rect 1360 5990 1600 6000
rect 2520 5990 3160 6000
rect 3280 5990 3760 6000
rect 4080 5990 4320 6000
rect 5240 5990 5320 6000
rect 9480 5990 9640 6000
rect 9720 5990 9840 6000
rect 1360 5980 1600 5990
rect 2520 5980 3160 5990
rect 3280 5980 3760 5990
rect 4080 5980 4320 5990
rect 5240 5980 5320 5990
rect 9480 5980 9640 5990
rect 9720 5980 9840 5990
rect 1200 5970 1240 5980
rect 1280 5970 1640 5980
rect 2560 5970 3120 5980
rect 3280 5970 3760 5980
rect 4160 5970 4320 5980
rect 5200 5970 5320 5980
rect 9520 5970 9680 5980
rect 9760 5970 9880 5980
rect 1200 5960 1240 5970
rect 1280 5960 1640 5970
rect 2560 5960 3120 5970
rect 3280 5960 3760 5970
rect 4160 5960 4320 5970
rect 5200 5960 5320 5970
rect 9520 5960 9680 5970
rect 9760 5960 9880 5970
rect 1200 5950 1240 5960
rect 1280 5950 1640 5960
rect 2560 5950 3120 5960
rect 3280 5950 3760 5960
rect 4160 5950 4320 5960
rect 5200 5950 5320 5960
rect 9520 5950 9680 5960
rect 9760 5950 9880 5960
rect 1200 5940 1240 5950
rect 1280 5940 1640 5950
rect 2560 5940 3120 5950
rect 3280 5940 3760 5950
rect 4160 5940 4320 5950
rect 5200 5940 5320 5950
rect 9520 5940 9680 5950
rect 9760 5940 9880 5950
rect 1080 5930 1160 5940
rect 1200 5930 1680 5940
rect 2600 5930 3080 5940
rect 3280 5930 3760 5940
rect 4240 5930 4280 5940
rect 5160 5930 5320 5940
rect 9520 5930 9680 5940
rect 9760 5930 9880 5940
rect 1080 5920 1160 5930
rect 1200 5920 1680 5930
rect 2600 5920 3080 5930
rect 3280 5920 3760 5930
rect 4240 5920 4280 5930
rect 5160 5920 5320 5930
rect 9520 5920 9680 5930
rect 9760 5920 9880 5930
rect 1080 5910 1160 5920
rect 1200 5910 1680 5920
rect 2600 5910 3080 5920
rect 3280 5910 3760 5920
rect 4240 5910 4280 5920
rect 5160 5910 5320 5920
rect 9520 5910 9680 5920
rect 9760 5910 9880 5920
rect 1080 5900 1160 5910
rect 1200 5900 1680 5910
rect 2600 5900 3080 5910
rect 3280 5900 3760 5910
rect 4240 5900 4280 5910
rect 5160 5900 5320 5910
rect 9520 5900 9680 5910
rect 9760 5900 9880 5910
rect 1120 5890 1720 5900
rect 2680 5890 3000 5900
rect 3280 5890 3720 5900
rect 5160 5890 5320 5900
rect 6840 5890 6920 5900
rect 9440 5890 9720 5900
rect 9760 5890 9880 5900
rect 1120 5880 1720 5890
rect 2680 5880 3000 5890
rect 3280 5880 3720 5890
rect 5160 5880 5320 5890
rect 6840 5880 6920 5890
rect 9440 5880 9720 5890
rect 9760 5880 9880 5890
rect 1120 5870 1720 5880
rect 2680 5870 3000 5880
rect 3280 5870 3720 5880
rect 5160 5870 5320 5880
rect 6840 5870 6920 5880
rect 9440 5870 9720 5880
rect 9760 5870 9880 5880
rect 1120 5860 1720 5870
rect 2680 5860 3000 5870
rect 3280 5860 3720 5870
rect 5160 5860 5320 5870
rect 6840 5860 6920 5870
rect 9440 5860 9720 5870
rect 9760 5860 9880 5870
rect 1000 5850 1840 5860
rect 2720 5850 2840 5860
rect 3280 5850 3720 5860
rect 5120 5850 5280 5860
rect 6840 5850 6920 5860
rect 9360 5850 9880 5860
rect 1000 5840 1840 5850
rect 2720 5840 2840 5850
rect 3280 5840 3720 5850
rect 5120 5840 5280 5850
rect 6840 5840 6920 5850
rect 9360 5840 9880 5850
rect 1000 5830 1840 5840
rect 2720 5830 2840 5840
rect 3280 5830 3720 5840
rect 5120 5830 5280 5840
rect 6840 5830 6920 5840
rect 9360 5830 9880 5840
rect 1000 5820 1840 5830
rect 2720 5820 2840 5830
rect 3280 5820 3720 5830
rect 5120 5820 5280 5830
rect 6840 5820 6920 5830
rect 9360 5820 9880 5830
rect 920 5810 1840 5820
rect 3320 5810 3720 5820
rect 5120 5810 5280 5820
rect 6880 5810 6920 5820
rect 9280 5810 9920 5820
rect 920 5800 1840 5810
rect 3320 5800 3720 5810
rect 5120 5800 5280 5810
rect 6880 5800 6920 5810
rect 9280 5800 9920 5810
rect 920 5790 1840 5800
rect 3320 5790 3720 5800
rect 5120 5790 5280 5800
rect 6880 5790 6920 5800
rect 9280 5790 9920 5800
rect 920 5780 1840 5790
rect 3320 5780 3720 5790
rect 5120 5780 5280 5790
rect 6880 5780 6920 5790
rect 9280 5780 9920 5790
rect 920 5770 1840 5780
rect 3320 5770 3720 5780
rect 5120 5770 5280 5780
rect 9080 5770 9160 5780
rect 9200 5770 9920 5780
rect 920 5760 1840 5770
rect 3320 5760 3720 5770
rect 5120 5760 5280 5770
rect 9080 5760 9160 5770
rect 9200 5760 9920 5770
rect 920 5750 1840 5760
rect 3320 5750 3720 5760
rect 5120 5750 5280 5760
rect 9080 5750 9160 5760
rect 9200 5750 9920 5760
rect 920 5740 1840 5750
rect 3320 5740 3720 5750
rect 5120 5740 5280 5750
rect 9080 5740 9160 5750
rect 9200 5740 9920 5750
rect 880 5730 1160 5740
rect 1240 5730 1840 5740
rect 3320 5730 3720 5740
rect 3880 5730 3920 5740
rect 5120 5730 5280 5740
rect 8760 5730 8800 5740
rect 9040 5730 9920 5740
rect 880 5720 1160 5730
rect 1240 5720 1840 5730
rect 3320 5720 3720 5730
rect 3880 5720 3920 5730
rect 5120 5720 5280 5730
rect 8760 5720 8800 5730
rect 9040 5720 9920 5730
rect 880 5710 1160 5720
rect 1240 5710 1840 5720
rect 3320 5710 3720 5720
rect 3880 5710 3920 5720
rect 5120 5710 5280 5720
rect 8760 5710 8800 5720
rect 9040 5710 9920 5720
rect 880 5700 1160 5710
rect 1240 5700 1840 5710
rect 3320 5700 3720 5710
rect 3880 5700 3920 5710
rect 5120 5700 5280 5710
rect 8760 5700 8800 5710
rect 9040 5700 9920 5710
rect 840 5690 1080 5700
rect 1200 5690 1840 5700
rect 3320 5690 3680 5700
rect 5160 5690 5280 5700
rect 8760 5690 8920 5700
rect 9000 5690 9960 5700
rect 840 5680 1080 5690
rect 1200 5680 1840 5690
rect 3320 5680 3680 5690
rect 5160 5680 5280 5690
rect 8760 5680 8920 5690
rect 9000 5680 9960 5690
rect 840 5670 1080 5680
rect 1200 5670 1840 5680
rect 3320 5670 3680 5680
rect 5160 5670 5280 5680
rect 8760 5670 8920 5680
rect 9000 5670 9960 5680
rect 840 5660 1080 5670
rect 1200 5660 1840 5670
rect 3320 5660 3680 5670
rect 5160 5660 5280 5670
rect 8760 5660 8920 5670
rect 9000 5660 9960 5670
rect 840 5650 1840 5660
rect 3320 5650 3680 5660
rect 5160 5650 5240 5660
rect 6880 5650 6920 5660
rect 8560 5650 9960 5660
rect 840 5640 1840 5650
rect 3320 5640 3680 5650
rect 5160 5640 5240 5650
rect 6880 5640 6920 5650
rect 8560 5640 9960 5650
rect 840 5630 1840 5640
rect 3320 5630 3680 5640
rect 5160 5630 5240 5640
rect 6880 5630 6920 5640
rect 8560 5630 9960 5640
rect 840 5620 1840 5630
rect 3320 5620 3680 5630
rect 5160 5620 5240 5630
rect 6880 5620 6920 5630
rect 8560 5620 9960 5630
rect 760 5610 1840 5620
rect 3320 5610 3400 5620
rect 3480 5610 3640 5620
rect 3720 5610 3760 5620
rect 5120 5610 5240 5620
rect 8480 5610 8920 5620
rect 9080 5610 9960 5620
rect 760 5600 1840 5610
rect 3320 5600 3400 5610
rect 3480 5600 3640 5610
rect 3720 5600 3760 5610
rect 5120 5600 5240 5610
rect 8480 5600 8920 5610
rect 9080 5600 9960 5610
rect 760 5590 1840 5600
rect 3320 5590 3400 5600
rect 3480 5590 3640 5600
rect 3720 5590 3760 5600
rect 5120 5590 5240 5600
rect 8480 5590 8920 5600
rect 9080 5590 9960 5600
rect 760 5580 1840 5590
rect 3320 5580 3400 5590
rect 3480 5580 3640 5590
rect 3720 5580 3760 5590
rect 5120 5580 5240 5590
rect 8480 5580 8920 5590
rect 9080 5580 9960 5590
rect 680 5570 1880 5580
rect 3320 5570 3440 5580
rect 3520 5570 3640 5580
rect 5120 5570 5240 5580
rect 5720 5570 5840 5580
rect 8400 5570 8840 5580
rect 9120 5570 9990 5580
rect 680 5560 1880 5570
rect 3320 5560 3440 5570
rect 3520 5560 3640 5570
rect 5120 5560 5240 5570
rect 5720 5560 5840 5570
rect 8400 5560 8840 5570
rect 9120 5560 9990 5570
rect 680 5550 1880 5560
rect 3320 5550 3440 5560
rect 3520 5550 3640 5560
rect 5120 5550 5240 5560
rect 5720 5550 5840 5560
rect 8400 5550 8840 5560
rect 9120 5550 9990 5560
rect 680 5540 1880 5550
rect 3320 5540 3440 5550
rect 3520 5540 3640 5550
rect 5120 5540 5240 5550
rect 5720 5540 5840 5550
rect 8400 5540 8840 5550
rect 9120 5540 9990 5550
rect 680 5530 920 5540
rect 960 5530 1880 5540
rect 3320 5530 3480 5540
rect 3520 5530 3640 5540
rect 5160 5530 5240 5540
rect 6280 5530 6440 5540
rect 8200 5530 8680 5540
rect 9120 5530 9990 5540
rect 680 5520 920 5530
rect 960 5520 1880 5530
rect 3320 5520 3480 5530
rect 3520 5520 3640 5530
rect 5160 5520 5240 5530
rect 6280 5520 6440 5530
rect 8200 5520 8680 5530
rect 9120 5520 9990 5530
rect 680 5510 920 5520
rect 960 5510 1880 5520
rect 3320 5510 3480 5520
rect 3520 5510 3640 5520
rect 5160 5510 5240 5520
rect 6280 5510 6440 5520
rect 8200 5510 8680 5520
rect 9120 5510 9990 5520
rect 680 5500 920 5510
rect 960 5500 1880 5510
rect 3320 5500 3480 5510
rect 3520 5500 3640 5510
rect 5160 5500 5240 5510
rect 6280 5500 6440 5510
rect 8200 5500 8680 5510
rect 9120 5500 9990 5510
rect 640 5490 920 5500
rect 1000 5490 1880 5500
rect 3320 5490 3560 5500
rect 5160 5490 5240 5500
rect 6240 5490 6360 5500
rect 8160 5490 8520 5500
rect 9160 5490 9990 5500
rect 640 5480 920 5490
rect 1000 5480 1880 5490
rect 3320 5480 3560 5490
rect 5160 5480 5240 5490
rect 6240 5480 6360 5490
rect 8160 5480 8520 5490
rect 9160 5480 9990 5490
rect 640 5470 920 5480
rect 1000 5470 1880 5480
rect 3320 5470 3560 5480
rect 5160 5470 5240 5480
rect 6240 5470 6360 5480
rect 8160 5470 8520 5480
rect 9160 5470 9990 5480
rect 640 5460 920 5470
rect 1000 5460 1880 5470
rect 3320 5460 3560 5470
rect 5160 5460 5240 5470
rect 6240 5460 6360 5470
rect 8160 5460 8520 5470
rect 9160 5460 9990 5470
rect 600 5450 1920 5460
rect 2440 5450 2560 5460
rect 3320 5450 3560 5460
rect 5160 5450 5240 5460
rect 5720 5450 5800 5460
rect 6240 5450 6360 5460
rect 8160 5450 8400 5460
rect 9120 5450 9520 5460
rect 9600 5450 9990 5460
rect 600 5440 1920 5450
rect 2440 5440 2560 5450
rect 3320 5440 3560 5450
rect 5160 5440 5240 5450
rect 5720 5440 5800 5450
rect 6240 5440 6360 5450
rect 8160 5440 8400 5450
rect 9120 5440 9520 5450
rect 9600 5440 9990 5450
rect 600 5430 1920 5440
rect 2440 5430 2560 5440
rect 3320 5430 3560 5440
rect 5160 5430 5240 5440
rect 5720 5430 5800 5440
rect 6240 5430 6360 5440
rect 8160 5430 8400 5440
rect 9120 5430 9520 5440
rect 9600 5430 9990 5440
rect 600 5420 1920 5430
rect 2440 5420 2560 5430
rect 3320 5420 3560 5430
rect 5160 5420 5240 5430
rect 5720 5420 5800 5430
rect 6240 5420 6360 5430
rect 8160 5420 8400 5430
rect 9120 5420 9520 5430
rect 9600 5420 9990 5430
rect 600 5410 1920 5420
rect 2440 5410 2560 5420
rect 3240 5410 3560 5420
rect 5120 5410 5200 5420
rect 5560 5410 5840 5420
rect 6240 5410 6560 5420
rect 8160 5410 8280 5420
rect 9120 5410 9400 5420
rect 9440 5410 9480 5420
rect 9600 5410 9990 5420
rect 600 5400 1920 5410
rect 2440 5400 2560 5410
rect 3240 5400 3560 5410
rect 5120 5400 5200 5410
rect 5560 5400 5840 5410
rect 6240 5400 6560 5410
rect 8160 5400 8280 5410
rect 9120 5400 9400 5410
rect 9440 5400 9480 5410
rect 9600 5400 9990 5410
rect 600 5390 1920 5400
rect 2440 5390 2560 5400
rect 3240 5390 3560 5400
rect 5120 5390 5200 5400
rect 5560 5390 5840 5400
rect 6240 5390 6560 5400
rect 8160 5390 8280 5400
rect 9120 5390 9400 5400
rect 9440 5390 9480 5400
rect 9600 5390 9990 5400
rect 600 5380 1920 5390
rect 2440 5380 2560 5390
rect 3240 5380 3560 5390
rect 5120 5380 5200 5390
rect 5560 5380 5840 5390
rect 6240 5380 6560 5390
rect 8160 5380 8280 5390
rect 9120 5380 9400 5390
rect 9440 5380 9480 5390
rect 9600 5380 9990 5390
rect 560 5370 1920 5380
rect 2440 5370 2480 5380
rect 2520 5370 2560 5380
rect 3040 5370 3480 5380
rect 3520 5370 3560 5380
rect 5120 5370 5200 5380
rect 5760 5370 5840 5380
rect 6200 5370 6360 5380
rect 6400 5370 6640 5380
rect 7800 5370 7840 5380
rect 8960 5370 9240 5380
rect 9600 5370 9990 5380
rect 560 5360 1920 5370
rect 2440 5360 2480 5370
rect 2520 5360 2560 5370
rect 3040 5360 3480 5370
rect 3520 5360 3560 5370
rect 5120 5360 5200 5370
rect 5760 5360 5840 5370
rect 6200 5360 6360 5370
rect 6400 5360 6640 5370
rect 7800 5360 7840 5370
rect 8960 5360 9240 5370
rect 9600 5360 9990 5370
rect 560 5350 1920 5360
rect 2440 5350 2480 5360
rect 2520 5350 2560 5360
rect 3040 5350 3480 5360
rect 3520 5350 3560 5360
rect 5120 5350 5200 5360
rect 5760 5350 5840 5360
rect 6200 5350 6360 5360
rect 6400 5350 6640 5360
rect 7800 5350 7840 5360
rect 8960 5350 9240 5360
rect 9600 5350 9990 5360
rect 560 5340 1920 5350
rect 2440 5340 2480 5350
rect 2520 5340 2560 5350
rect 3040 5340 3480 5350
rect 3520 5340 3560 5350
rect 5120 5340 5200 5350
rect 5760 5340 5840 5350
rect 6200 5340 6360 5350
rect 6400 5340 6640 5350
rect 7800 5340 7840 5350
rect 8960 5340 9240 5350
rect 9600 5340 9990 5350
rect 600 5330 1920 5340
rect 3040 5330 3520 5340
rect 7720 5330 7840 5340
rect 8800 5330 9120 5340
rect 9160 5330 9240 5340
rect 9480 5330 9520 5340
rect 9640 5330 9990 5340
rect 600 5320 1920 5330
rect 3040 5320 3520 5330
rect 7720 5320 7840 5330
rect 8800 5320 9120 5330
rect 9160 5320 9240 5330
rect 9480 5320 9520 5330
rect 9640 5320 9990 5330
rect 600 5310 1920 5320
rect 3040 5310 3520 5320
rect 7720 5310 7840 5320
rect 8800 5310 9120 5320
rect 9160 5310 9240 5320
rect 9480 5310 9520 5320
rect 9640 5310 9990 5320
rect 600 5300 1920 5310
rect 3040 5300 3520 5310
rect 7720 5300 7840 5310
rect 8800 5300 9120 5310
rect 9160 5300 9240 5310
rect 9480 5300 9520 5310
rect 9640 5300 9990 5310
rect 640 5290 1920 5300
rect 3000 5290 3520 5300
rect 7640 5290 7840 5300
rect 8680 5290 8920 5300
rect 8960 5290 9040 5300
rect 9200 5290 9240 5300
rect 9480 5290 9520 5300
rect 9640 5290 9840 5300
rect 640 5280 1920 5290
rect 3000 5280 3520 5290
rect 7640 5280 7840 5290
rect 8680 5280 8920 5290
rect 8960 5280 9040 5290
rect 9200 5280 9240 5290
rect 9480 5280 9520 5290
rect 9640 5280 9840 5290
rect 640 5270 1920 5280
rect 3000 5270 3520 5280
rect 7640 5270 7840 5280
rect 8680 5270 8920 5280
rect 8960 5270 9040 5280
rect 9200 5270 9240 5280
rect 9480 5270 9520 5280
rect 9640 5270 9840 5280
rect 640 5260 1920 5270
rect 3000 5260 3520 5270
rect 7640 5260 7840 5270
rect 8680 5260 8920 5270
rect 8960 5260 9040 5270
rect 9200 5260 9240 5270
rect 9480 5260 9520 5270
rect 9640 5260 9840 5270
rect 640 5250 1960 5260
rect 2960 5250 3480 5260
rect 7480 5250 7560 5260
rect 7680 5250 7840 5260
rect 8520 5250 8800 5260
rect 9000 5250 9040 5260
rect 9200 5250 9280 5260
rect 9400 5250 9440 5260
rect 9480 5250 9720 5260
rect 640 5240 1960 5250
rect 2960 5240 3480 5250
rect 7480 5240 7560 5250
rect 7680 5240 7840 5250
rect 8520 5240 8800 5250
rect 9000 5240 9040 5250
rect 9200 5240 9280 5250
rect 9400 5240 9440 5250
rect 9480 5240 9720 5250
rect 640 5230 1960 5240
rect 2960 5230 3480 5240
rect 7480 5230 7560 5240
rect 7680 5230 7840 5240
rect 8520 5230 8800 5240
rect 9000 5230 9040 5240
rect 9200 5230 9280 5240
rect 9400 5230 9440 5240
rect 9480 5230 9720 5240
rect 640 5220 1960 5230
rect 2960 5220 3480 5230
rect 7480 5220 7560 5230
rect 7680 5220 7840 5230
rect 8520 5220 8800 5230
rect 9000 5220 9040 5230
rect 9200 5220 9280 5230
rect 9400 5220 9440 5230
rect 9480 5220 9720 5230
rect 720 5210 1960 5220
rect 3000 5210 3480 5220
rect 7440 5210 7520 5220
rect 7680 5210 7840 5220
rect 8360 5210 8640 5220
rect 9200 5210 9280 5220
rect 9400 5210 9520 5220
rect 9600 5210 9680 5220
rect 720 5200 1960 5210
rect 3000 5200 3480 5210
rect 7440 5200 7520 5210
rect 7680 5200 7840 5210
rect 8360 5200 8640 5210
rect 9200 5200 9280 5210
rect 9400 5200 9520 5210
rect 9600 5200 9680 5210
rect 720 5190 1960 5200
rect 3000 5190 3480 5200
rect 7440 5190 7520 5200
rect 7680 5190 7840 5200
rect 8360 5190 8640 5200
rect 9200 5190 9280 5200
rect 9400 5190 9520 5200
rect 9600 5190 9680 5200
rect 720 5180 1960 5190
rect 3000 5180 3480 5190
rect 7440 5180 7520 5190
rect 7680 5180 7840 5190
rect 8360 5180 8640 5190
rect 9200 5180 9280 5190
rect 9400 5180 9520 5190
rect 9600 5180 9680 5190
rect 720 5170 1800 5180
rect 1880 5170 1960 5180
rect 3040 5170 3440 5180
rect 7440 5170 7560 5180
rect 7600 5170 7880 5180
rect 8280 5170 8600 5180
rect 9120 5170 9160 5180
rect 9200 5170 9360 5180
rect 9640 5170 9680 5180
rect 9760 5170 9800 5180
rect 9920 5170 9960 5180
rect 720 5160 1800 5170
rect 1880 5160 1960 5170
rect 3040 5160 3440 5170
rect 7440 5160 7560 5170
rect 7600 5160 7880 5170
rect 8280 5160 8600 5170
rect 9120 5160 9160 5170
rect 9200 5160 9360 5170
rect 9640 5160 9680 5170
rect 9760 5160 9800 5170
rect 9920 5160 9960 5170
rect 720 5150 1800 5160
rect 1880 5150 1960 5160
rect 3040 5150 3440 5160
rect 7440 5150 7560 5160
rect 7600 5150 7880 5160
rect 8280 5150 8600 5160
rect 9120 5150 9160 5160
rect 9200 5150 9360 5160
rect 9640 5150 9680 5160
rect 9760 5150 9800 5160
rect 9920 5150 9960 5160
rect 720 5140 1800 5150
rect 1880 5140 1960 5150
rect 3040 5140 3440 5150
rect 7440 5140 7560 5150
rect 7600 5140 7880 5150
rect 8280 5140 8600 5150
rect 9120 5140 9160 5150
rect 9200 5140 9360 5150
rect 9640 5140 9680 5150
rect 9760 5140 9800 5150
rect 9920 5140 9960 5150
rect 760 5130 1800 5140
rect 1880 5130 1960 5140
rect 3040 5130 3400 5140
rect 7440 5130 7880 5140
rect 8240 5130 8400 5140
rect 8520 5130 8640 5140
rect 8720 5130 8760 5140
rect 9040 5130 9240 5140
rect 9640 5130 9720 5140
rect 9920 5130 9990 5140
rect 760 5120 1800 5130
rect 1880 5120 1960 5130
rect 3040 5120 3400 5130
rect 7440 5120 7880 5130
rect 8240 5120 8400 5130
rect 8520 5120 8640 5130
rect 8720 5120 8760 5130
rect 9040 5120 9240 5130
rect 9640 5120 9720 5130
rect 9920 5120 9990 5130
rect 760 5110 1800 5120
rect 1880 5110 1960 5120
rect 3040 5110 3400 5120
rect 7440 5110 7880 5120
rect 8240 5110 8400 5120
rect 8520 5110 8640 5120
rect 8720 5110 8760 5120
rect 9040 5110 9240 5120
rect 9640 5110 9720 5120
rect 9920 5110 9990 5120
rect 760 5100 1800 5110
rect 1880 5100 1960 5110
rect 3040 5100 3400 5110
rect 7440 5100 7880 5110
rect 8240 5100 8400 5110
rect 8520 5100 8640 5110
rect 8720 5100 8760 5110
rect 9040 5100 9240 5110
rect 9640 5100 9720 5110
rect 9920 5100 9990 5110
rect 640 5090 680 5100
rect 760 5090 1760 5100
rect 1880 5090 1960 5100
rect 2960 5090 3400 5100
rect 7440 5090 7880 5100
rect 8040 5090 8120 5100
rect 8520 5090 8640 5100
rect 8720 5090 8760 5100
rect 8920 5090 9080 5100
rect 9320 5090 9360 5100
rect 9480 5090 9520 5100
rect 9640 5090 9720 5100
rect 9840 5090 9990 5100
rect 640 5080 680 5090
rect 760 5080 1760 5090
rect 1880 5080 1960 5090
rect 2960 5080 3400 5090
rect 7440 5080 7880 5090
rect 8040 5080 8120 5090
rect 8520 5080 8640 5090
rect 8720 5080 8760 5090
rect 8920 5080 9080 5090
rect 9320 5080 9360 5090
rect 9480 5080 9520 5090
rect 9640 5080 9720 5090
rect 9840 5080 9990 5090
rect 640 5070 680 5080
rect 760 5070 1760 5080
rect 1880 5070 1960 5080
rect 2960 5070 3400 5080
rect 7440 5070 7880 5080
rect 8040 5070 8120 5080
rect 8520 5070 8640 5080
rect 8720 5070 8760 5080
rect 8920 5070 9080 5080
rect 9320 5070 9360 5080
rect 9480 5070 9520 5080
rect 9640 5070 9720 5080
rect 9840 5070 9990 5080
rect 640 5060 680 5070
rect 760 5060 1760 5070
rect 1880 5060 1960 5070
rect 2960 5060 3400 5070
rect 7440 5060 7880 5070
rect 8040 5060 8120 5070
rect 8520 5060 8640 5070
rect 8720 5060 8760 5070
rect 8920 5060 9080 5070
rect 9320 5060 9360 5070
rect 9480 5060 9520 5070
rect 9640 5060 9720 5070
rect 9840 5060 9990 5070
rect 640 5050 1760 5060
rect 1880 5050 2000 5060
rect 3040 5050 3360 5060
rect 7480 5050 7880 5060
rect 8520 5050 8680 5060
rect 8720 5050 8960 5060
rect 9200 5050 9280 5060
rect 9320 5050 9360 5060
rect 9640 5050 9990 5060
rect 640 5040 1760 5050
rect 1880 5040 2000 5050
rect 3040 5040 3360 5050
rect 7480 5040 7880 5050
rect 8520 5040 8680 5050
rect 8720 5040 8960 5050
rect 9200 5040 9280 5050
rect 9320 5040 9360 5050
rect 9640 5040 9990 5050
rect 640 5030 1760 5040
rect 1880 5030 2000 5040
rect 3040 5030 3360 5040
rect 7480 5030 7880 5040
rect 8520 5030 8680 5040
rect 8720 5030 8960 5040
rect 9200 5030 9280 5040
rect 9320 5030 9360 5040
rect 9640 5030 9990 5040
rect 640 5020 1760 5030
rect 1880 5020 2000 5030
rect 3040 5020 3360 5030
rect 7480 5020 7880 5030
rect 8520 5020 8680 5030
rect 8720 5020 8960 5030
rect 9200 5020 9280 5030
rect 9320 5020 9360 5030
rect 9640 5020 9990 5030
rect 480 5010 1760 5020
rect 1840 5010 2000 5020
rect 3040 5010 3320 5020
rect 7360 5010 7880 5020
rect 8560 5010 8760 5020
rect 8840 5010 8880 5020
rect 9080 5010 9120 5020
rect 9200 5010 9280 5020
rect 9360 5010 9400 5020
rect 9520 5010 9990 5020
rect 480 5000 1760 5010
rect 1840 5000 2000 5010
rect 3040 5000 3320 5010
rect 7360 5000 7880 5010
rect 8560 5000 8760 5010
rect 8840 5000 8880 5010
rect 9080 5000 9120 5010
rect 9200 5000 9280 5010
rect 9360 5000 9400 5010
rect 9520 5000 9990 5010
rect 480 4990 1760 5000
rect 1840 4990 2000 5000
rect 3040 4990 3320 5000
rect 7360 4990 7880 5000
rect 8560 4990 8760 5000
rect 8840 4990 8880 5000
rect 9080 4990 9120 5000
rect 9200 4990 9280 5000
rect 9360 4990 9400 5000
rect 9520 4990 9990 5000
rect 480 4980 1760 4990
rect 1840 4980 2000 4990
rect 3040 4980 3320 4990
rect 7360 4980 7880 4990
rect 8560 4980 8760 4990
rect 8840 4980 8880 4990
rect 9080 4980 9120 4990
rect 9200 4980 9280 4990
rect 9360 4980 9400 4990
rect 9520 4980 9990 4990
rect 560 4970 2080 4980
rect 2960 4970 3320 4980
rect 7360 4970 7800 4980
rect 8480 4970 8600 4980
rect 9360 4970 9520 4980
rect 9720 4970 9990 4980
rect 560 4960 2080 4970
rect 2960 4960 3320 4970
rect 7360 4960 7800 4970
rect 8480 4960 8600 4970
rect 9360 4960 9520 4970
rect 9720 4960 9990 4970
rect 560 4950 2080 4960
rect 2960 4950 3320 4960
rect 7360 4950 7800 4960
rect 8480 4950 8600 4960
rect 9360 4950 9520 4960
rect 9720 4950 9990 4960
rect 560 4940 2080 4950
rect 2960 4940 3320 4950
rect 7360 4940 7800 4950
rect 8480 4940 8600 4950
rect 9360 4940 9520 4950
rect 9720 4940 9990 4950
rect 720 4930 1040 4940
rect 1080 4930 2160 4940
rect 2880 4930 3280 4940
rect 4200 4930 4360 4940
rect 4400 4930 4440 4940
rect 7360 4930 7680 4940
rect 8280 4930 8480 4940
rect 9320 4930 9440 4940
rect 9720 4930 9990 4940
rect 720 4920 1040 4930
rect 1080 4920 2160 4930
rect 2880 4920 3280 4930
rect 4200 4920 4360 4930
rect 4400 4920 4440 4930
rect 7360 4920 7680 4930
rect 8280 4920 8480 4930
rect 9320 4920 9440 4930
rect 9720 4920 9990 4930
rect 720 4910 1040 4920
rect 1080 4910 2160 4920
rect 2880 4910 3280 4920
rect 4200 4910 4360 4920
rect 4400 4910 4440 4920
rect 7360 4910 7680 4920
rect 8280 4910 8480 4920
rect 9320 4910 9440 4920
rect 9720 4910 9990 4920
rect 720 4900 1040 4910
rect 1080 4900 2160 4910
rect 2880 4900 3280 4910
rect 4200 4900 4360 4910
rect 4400 4900 4440 4910
rect 7360 4900 7680 4910
rect 8280 4900 8480 4910
rect 9320 4900 9440 4910
rect 9720 4900 9990 4910
rect 760 4890 1040 4900
rect 1080 4890 2200 4900
rect 2800 4890 3160 4900
rect 3200 4890 3280 4900
rect 4080 4890 4160 4900
rect 4200 4890 4480 4900
rect 4680 4890 4720 4900
rect 6200 4890 6280 4900
rect 7400 4890 7680 4900
rect 8160 4890 8320 4900
rect 8360 4890 8440 4900
rect 8960 4890 9000 4900
rect 9040 4890 9080 4900
rect 9720 4890 9990 4900
rect 760 4880 1040 4890
rect 1080 4880 2200 4890
rect 2800 4880 3160 4890
rect 3200 4880 3280 4890
rect 4080 4880 4160 4890
rect 4200 4880 4480 4890
rect 4680 4880 4720 4890
rect 6200 4880 6280 4890
rect 7400 4880 7680 4890
rect 8160 4880 8320 4890
rect 8360 4880 8440 4890
rect 8960 4880 9000 4890
rect 9040 4880 9080 4890
rect 9720 4880 9990 4890
rect 760 4870 1040 4880
rect 1080 4870 2200 4880
rect 2800 4870 3160 4880
rect 3200 4870 3280 4880
rect 4080 4870 4160 4880
rect 4200 4870 4480 4880
rect 4680 4870 4720 4880
rect 6200 4870 6280 4880
rect 7400 4870 7680 4880
rect 8160 4870 8320 4880
rect 8360 4870 8440 4880
rect 8960 4870 9000 4880
rect 9040 4870 9080 4880
rect 9720 4870 9990 4880
rect 760 4860 1040 4870
rect 1080 4860 2200 4870
rect 2800 4860 3160 4870
rect 3200 4860 3280 4870
rect 4080 4860 4160 4870
rect 4200 4860 4480 4870
rect 4680 4860 4720 4870
rect 6200 4860 6280 4870
rect 7400 4860 7680 4870
rect 8160 4860 8320 4870
rect 8360 4860 8440 4870
rect 8960 4860 9000 4870
rect 9040 4860 9080 4870
rect 9720 4860 9990 4870
rect 800 4850 1040 4860
rect 1120 4850 2320 4860
rect 2800 4850 3080 4860
rect 3160 4850 3240 4860
rect 3280 4850 3320 4860
rect 3880 4850 3920 4860
rect 4000 4850 4880 4860
rect 7400 4850 7680 4860
rect 8080 4850 8200 4860
rect 8400 4850 8440 4860
rect 8800 4850 8840 4860
rect 8880 4850 9040 4860
rect 9760 4850 9990 4860
rect 800 4840 1040 4850
rect 1120 4840 2320 4850
rect 2800 4840 3080 4850
rect 3160 4840 3240 4850
rect 3280 4840 3320 4850
rect 3880 4840 3920 4850
rect 4000 4840 4880 4850
rect 7400 4840 7680 4850
rect 8080 4840 8200 4850
rect 8400 4840 8440 4850
rect 8800 4840 8840 4850
rect 8880 4840 9040 4850
rect 9760 4840 9990 4850
rect 800 4830 1040 4840
rect 1120 4830 2320 4840
rect 2800 4830 3080 4840
rect 3160 4830 3240 4840
rect 3280 4830 3320 4840
rect 3880 4830 3920 4840
rect 4000 4830 4880 4840
rect 7400 4830 7680 4840
rect 8080 4830 8200 4840
rect 8400 4830 8440 4840
rect 8800 4830 8840 4840
rect 8880 4830 9040 4840
rect 9760 4830 9990 4840
rect 800 4820 1040 4830
rect 1120 4820 2320 4830
rect 2800 4820 3080 4830
rect 3160 4820 3240 4830
rect 3280 4820 3320 4830
rect 3880 4820 3920 4830
rect 4000 4820 4880 4830
rect 7400 4820 7680 4830
rect 8080 4820 8200 4830
rect 8400 4820 8440 4830
rect 8800 4820 8840 4830
rect 8880 4820 9040 4830
rect 9760 4820 9990 4830
rect 480 4810 560 4820
rect 880 4810 1040 4820
rect 1120 4810 2360 4820
rect 2920 4810 3040 4820
rect 3160 4810 3200 4820
rect 3280 4810 3320 4820
rect 3640 4810 3720 4820
rect 3800 4810 3880 4820
rect 3960 4810 4920 4820
rect 5560 4810 5600 4820
rect 7360 4810 7680 4820
rect 7920 4810 7960 4820
rect 8400 4810 8480 4820
rect 8560 4810 8600 4820
rect 8760 4810 8920 4820
rect 8960 4810 9000 4820
rect 9360 4810 9400 4820
rect 9520 4810 9560 4820
rect 9720 4810 9990 4820
rect 480 4800 560 4810
rect 880 4800 1040 4810
rect 1120 4800 2360 4810
rect 2920 4800 3040 4810
rect 3160 4800 3200 4810
rect 3280 4800 3320 4810
rect 3640 4800 3720 4810
rect 3800 4800 3880 4810
rect 3960 4800 4920 4810
rect 5560 4800 5600 4810
rect 7360 4800 7680 4810
rect 7920 4800 7960 4810
rect 8400 4800 8480 4810
rect 8560 4800 8600 4810
rect 8760 4800 8920 4810
rect 8960 4800 9000 4810
rect 9360 4800 9400 4810
rect 9520 4800 9560 4810
rect 9720 4800 9990 4810
rect 480 4790 560 4800
rect 880 4790 1040 4800
rect 1120 4790 2360 4800
rect 2920 4790 3040 4800
rect 3160 4790 3200 4800
rect 3280 4790 3320 4800
rect 3640 4790 3720 4800
rect 3800 4790 3880 4800
rect 3960 4790 4920 4800
rect 5560 4790 5600 4800
rect 7360 4790 7680 4800
rect 7920 4790 7960 4800
rect 8400 4790 8480 4800
rect 8560 4790 8600 4800
rect 8760 4790 8920 4800
rect 8960 4790 9000 4800
rect 9360 4790 9400 4800
rect 9520 4790 9560 4800
rect 9720 4790 9990 4800
rect 480 4780 560 4790
rect 880 4780 1040 4790
rect 1120 4780 2360 4790
rect 2920 4780 3040 4790
rect 3160 4780 3200 4790
rect 3280 4780 3320 4790
rect 3640 4780 3720 4790
rect 3800 4780 3880 4790
rect 3960 4780 4920 4790
rect 5560 4780 5600 4790
rect 7360 4780 7680 4790
rect 7920 4780 7960 4790
rect 8400 4780 8480 4790
rect 8560 4780 8600 4790
rect 8760 4780 8920 4790
rect 8960 4780 9000 4790
rect 9360 4780 9400 4790
rect 9520 4780 9560 4790
rect 9720 4780 9990 4790
rect 360 4770 480 4780
rect 1000 4770 1040 4780
rect 1160 4770 2360 4780
rect 3120 4770 3240 4780
rect 3600 4770 3840 4780
rect 3880 4770 5040 4780
rect 5520 4770 5560 4780
rect 7400 4770 7880 4780
rect 8400 4770 8480 4780
rect 8560 4770 8800 4780
rect 9360 4770 9400 4780
rect 9520 4770 9880 4780
rect 360 4760 480 4770
rect 1000 4760 1040 4770
rect 1160 4760 2360 4770
rect 3120 4760 3240 4770
rect 3600 4760 3840 4770
rect 3880 4760 5040 4770
rect 5520 4760 5560 4770
rect 7400 4760 7880 4770
rect 8400 4760 8480 4770
rect 8560 4760 8800 4770
rect 9360 4760 9400 4770
rect 9520 4760 9880 4770
rect 360 4750 480 4760
rect 1000 4750 1040 4760
rect 1160 4750 2360 4760
rect 3120 4750 3240 4760
rect 3600 4750 3840 4760
rect 3880 4750 5040 4760
rect 5520 4750 5560 4760
rect 7400 4750 7880 4760
rect 8400 4750 8480 4760
rect 8560 4750 8800 4760
rect 9360 4750 9400 4760
rect 9520 4750 9880 4760
rect 360 4740 480 4750
rect 1000 4740 1040 4750
rect 1160 4740 2360 4750
rect 3120 4740 3240 4750
rect 3600 4740 3840 4750
rect 3880 4740 5040 4750
rect 5520 4740 5560 4750
rect 7400 4740 7880 4750
rect 8400 4740 8480 4750
rect 8560 4740 8800 4750
rect 9360 4740 9400 4750
rect 9520 4740 9880 4750
rect 440 4730 600 4740
rect 1040 4730 1080 4740
rect 1160 4730 2400 4740
rect 3120 4730 3240 4740
rect 3600 4730 3760 4740
rect 3800 4730 5080 4740
rect 5520 4730 5560 4740
rect 7440 4730 7720 4740
rect 8400 4730 8600 4740
rect 8680 4730 8760 4740
rect 9360 4730 9800 4740
rect 440 4720 600 4730
rect 1040 4720 1080 4730
rect 1160 4720 2400 4730
rect 3120 4720 3240 4730
rect 3600 4720 3760 4730
rect 3800 4720 5080 4730
rect 5520 4720 5560 4730
rect 7440 4720 7720 4730
rect 8400 4720 8600 4730
rect 8680 4720 8760 4730
rect 9360 4720 9800 4730
rect 440 4710 600 4720
rect 1040 4710 1080 4720
rect 1160 4710 2400 4720
rect 3120 4710 3240 4720
rect 3600 4710 3760 4720
rect 3800 4710 5080 4720
rect 5520 4710 5560 4720
rect 7440 4710 7720 4720
rect 8400 4710 8600 4720
rect 8680 4710 8760 4720
rect 9360 4710 9800 4720
rect 440 4700 600 4710
rect 1040 4700 1080 4710
rect 1160 4700 2400 4710
rect 3120 4700 3240 4710
rect 3600 4700 3760 4710
rect 3800 4700 5080 4710
rect 5520 4700 5560 4710
rect 7440 4700 7720 4710
rect 8400 4700 8600 4710
rect 8680 4700 8760 4710
rect 9360 4700 9800 4710
rect 520 4690 760 4700
rect 1040 4690 1120 4700
rect 1200 4690 2440 4700
rect 3200 4690 3240 4700
rect 3560 4690 5080 4700
rect 5520 4690 5560 4700
rect 7400 4690 7600 4700
rect 8280 4690 8480 4700
rect 8680 4690 8760 4700
rect 9280 4690 9800 4700
rect 520 4680 760 4690
rect 1040 4680 1120 4690
rect 1200 4680 2440 4690
rect 3200 4680 3240 4690
rect 3560 4680 5080 4690
rect 5520 4680 5560 4690
rect 7400 4680 7600 4690
rect 8280 4680 8480 4690
rect 8680 4680 8760 4690
rect 9280 4680 9800 4690
rect 520 4670 760 4680
rect 1040 4670 1120 4680
rect 1200 4670 2440 4680
rect 3200 4670 3240 4680
rect 3560 4670 5080 4680
rect 5520 4670 5560 4680
rect 7400 4670 7600 4680
rect 8280 4670 8480 4680
rect 8680 4670 8760 4680
rect 9280 4670 9800 4680
rect 520 4660 760 4670
rect 1040 4660 1120 4670
rect 1200 4660 2440 4670
rect 3200 4660 3240 4670
rect 3560 4660 5080 4670
rect 5520 4660 5560 4670
rect 7400 4660 7600 4670
rect 8280 4660 8480 4670
rect 8680 4660 8760 4670
rect 9280 4660 9800 4670
rect 600 4650 840 4660
rect 1200 4650 2560 4660
rect 3200 4650 3280 4660
rect 3480 4650 5120 4660
rect 5560 4650 5720 4660
rect 6520 4650 6560 4660
rect 7400 4650 7480 4660
rect 7840 4650 7880 4660
rect 8120 4650 8280 4660
rect 8400 4650 8480 4660
rect 8560 4650 8600 4660
rect 8680 4650 8760 4660
rect 9280 4650 9760 4660
rect 600 4640 840 4650
rect 1200 4640 2560 4650
rect 3200 4640 3280 4650
rect 3480 4640 5120 4650
rect 5560 4640 5720 4650
rect 6520 4640 6560 4650
rect 7400 4640 7480 4650
rect 7840 4640 7880 4650
rect 8120 4640 8280 4650
rect 8400 4640 8480 4650
rect 8560 4640 8600 4650
rect 8680 4640 8760 4650
rect 9280 4640 9760 4650
rect 600 4630 840 4640
rect 1200 4630 2560 4640
rect 3200 4630 3280 4640
rect 3480 4630 5120 4640
rect 5560 4630 5720 4640
rect 6520 4630 6560 4640
rect 7400 4630 7480 4640
rect 7840 4630 7880 4640
rect 8120 4630 8280 4640
rect 8400 4630 8480 4640
rect 8560 4630 8600 4640
rect 8680 4630 8760 4640
rect 9280 4630 9760 4640
rect 600 4620 840 4630
rect 1200 4620 2560 4630
rect 3200 4620 3280 4630
rect 3480 4620 5120 4630
rect 5560 4620 5720 4630
rect 6520 4620 6560 4630
rect 7400 4620 7480 4630
rect 7840 4620 7880 4630
rect 8120 4620 8280 4630
rect 8400 4620 8480 4630
rect 8560 4620 8600 4630
rect 8680 4620 8760 4630
rect 9280 4620 9760 4630
rect 680 4610 880 4620
rect 1240 4610 2840 4620
rect 3040 4610 3120 4620
rect 3480 4610 5200 4620
rect 5680 4610 5760 4620
rect 6280 4610 6520 4620
rect 7400 4610 7480 4620
rect 7960 4610 8080 4620
rect 8400 4610 8480 4620
rect 8680 4610 8800 4620
rect 8920 4610 8960 4620
rect 9280 4610 9720 4620
rect 680 4600 880 4610
rect 1240 4600 2840 4610
rect 3040 4600 3120 4610
rect 3480 4600 5200 4610
rect 5680 4600 5760 4610
rect 6280 4600 6520 4610
rect 7400 4600 7480 4610
rect 7960 4600 8080 4610
rect 8400 4600 8480 4610
rect 8680 4600 8800 4610
rect 8920 4600 8960 4610
rect 9280 4600 9720 4610
rect 680 4590 880 4600
rect 1240 4590 2840 4600
rect 3040 4590 3120 4600
rect 3480 4590 5200 4600
rect 5680 4590 5760 4600
rect 6280 4590 6520 4600
rect 7400 4590 7480 4600
rect 7960 4590 8080 4600
rect 8400 4590 8480 4600
rect 8680 4590 8800 4600
rect 8920 4590 8960 4600
rect 9280 4590 9720 4600
rect 680 4580 880 4590
rect 1240 4580 2840 4590
rect 3040 4580 3120 4590
rect 3480 4580 5200 4590
rect 5680 4580 5760 4590
rect 6280 4580 6520 4590
rect 7400 4580 7480 4590
rect 7960 4580 8080 4590
rect 8400 4580 8480 4590
rect 8680 4580 8800 4590
rect 8920 4580 8960 4590
rect 9280 4580 9720 4590
rect 720 4570 920 4580
rect 1240 4570 3040 4580
rect 3080 4570 3120 4580
rect 3480 4570 5200 4580
rect 5680 4570 5760 4580
rect 6320 4570 6480 4580
rect 7400 4570 7480 4580
rect 7800 4570 8000 4580
rect 8400 4570 8480 4580
rect 8680 4570 8920 4580
rect 9240 4570 9680 4580
rect 720 4560 920 4570
rect 1240 4560 3040 4570
rect 3080 4560 3120 4570
rect 3480 4560 5200 4570
rect 5680 4560 5760 4570
rect 6320 4560 6480 4570
rect 7400 4560 7480 4570
rect 7800 4560 8000 4570
rect 8400 4560 8480 4570
rect 8680 4560 8920 4570
rect 9240 4560 9680 4570
rect 720 4550 920 4560
rect 1240 4550 3040 4560
rect 3080 4550 3120 4560
rect 3480 4550 5200 4560
rect 5680 4550 5760 4560
rect 6320 4550 6480 4560
rect 7400 4550 7480 4560
rect 7800 4550 8000 4560
rect 8400 4550 8480 4560
rect 8680 4550 8920 4560
rect 9240 4550 9680 4560
rect 720 4540 920 4550
rect 1240 4540 3040 4550
rect 3080 4540 3120 4550
rect 3480 4540 5200 4550
rect 5680 4540 5760 4550
rect 6320 4540 6480 4550
rect 7400 4540 7480 4550
rect 7800 4540 8000 4550
rect 8400 4540 8480 4550
rect 8680 4540 8920 4550
rect 9240 4540 9680 4550
rect 760 4530 960 4540
rect 1160 4530 2960 4540
rect 3080 4530 3200 4540
rect 3440 4530 3880 4540
rect 3920 4530 5240 4540
rect 5720 4530 5760 4540
rect 6320 4530 6400 4540
rect 7440 4530 7480 4540
rect 7560 4530 7600 4540
rect 7680 4530 7800 4540
rect 8400 4530 8480 4540
rect 8520 4530 8920 4540
rect 9240 4530 9640 4540
rect 760 4520 960 4530
rect 1160 4520 2960 4530
rect 3080 4520 3200 4530
rect 3440 4520 3880 4530
rect 3920 4520 5240 4530
rect 5720 4520 5760 4530
rect 6320 4520 6400 4530
rect 7440 4520 7480 4530
rect 7560 4520 7600 4530
rect 7680 4520 7800 4530
rect 8400 4520 8480 4530
rect 8520 4520 8920 4530
rect 9240 4520 9640 4530
rect 760 4510 960 4520
rect 1160 4510 2960 4520
rect 3080 4510 3200 4520
rect 3440 4510 3880 4520
rect 3920 4510 5240 4520
rect 5720 4510 5760 4520
rect 6320 4510 6400 4520
rect 7440 4510 7480 4520
rect 7560 4510 7600 4520
rect 7680 4510 7800 4520
rect 8400 4510 8480 4520
rect 8520 4510 8920 4520
rect 9240 4510 9640 4520
rect 760 4500 960 4510
rect 1160 4500 2960 4510
rect 3080 4500 3200 4510
rect 3440 4500 3880 4510
rect 3920 4500 5240 4510
rect 5720 4500 5760 4510
rect 6320 4500 6400 4510
rect 7440 4500 7480 4510
rect 7560 4500 7600 4510
rect 7680 4500 7800 4510
rect 8400 4500 8480 4510
rect 8520 4500 8920 4510
rect 9240 4500 9640 4510
rect 640 4490 1000 4500
rect 1200 4490 3000 4500
rect 3120 4490 3240 4500
rect 3400 4490 3840 4500
rect 3960 4490 5280 4500
rect 6280 4490 6360 4500
rect 7440 4490 7760 4500
rect 8400 4490 8920 4500
rect 9240 4490 9600 4500
rect 640 4480 1000 4490
rect 1200 4480 3000 4490
rect 3120 4480 3240 4490
rect 3400 4480 3840 4490
rect 3960 4480 5280 4490
rect 6280 4480 6360 4490
rect 7440 4480 7760 4490
rect 8400 4480 8920 4490
rect 9240 4480 9600 4490
rect 640 4470 1000 4480
rect 1200 4470 3000 4480
rect 3120 4470 3240 4480
rect 3400 4470 3840 4480
rect 3960 4470 5280 4480
rect 6280 4470 6360 4480
rect 7440 4470 7760 4480
rect 8400 4470 8920 4480
rect 9240 4470 9600 4480
rect 640 4460 1000 4470
rect 1200 4460 3000 4470
rect 3120 4460 3240 4470
rect 3400 4460 3840 4470
rect 3960 4460 5280 4470
rect 6280 4460 6360 4470
rect 7440 4460 7760 4470
rect 8400 4460 8920 4470
rect 9240 4460 9600 4470
rect 480 4450 520 4460
rect 600 4450 1040 4460
rect 1160 4450 2800 4460
rect 2880 4450 2960 4460
rect 3400 4450 3840 4460
rect 3960 4450 4600 4460
rect 4680 4450 5280 4460
rect 6240 4450 6320 4460
rect 7440 4450 7760 4460
rect 8280 4450 8840 4460
rect 9240 4450 9560 4460
rect 9960 4450 9990 4460
rect 480 4440 520 4450
rect 600 4440 1040 4450
rect 1160 4440 2800 4450
rect 2880 4440 2960 4450
rect 3400 4440 3840 4450
rect 3960 4440 4600 4450
rect 4680 4440 5280 4450
rect 6240 4440 6320 4450
rect 7440 4440 7760 4450
rect 8280 4440 8840 4450
rect 9240 4440 9560 4450
rect 9960 4440 9990 4450
rect 480 4430 520 4440
rect 600 4430 1040 4440
rect 1160 4430 2800 4440
rect 2880 4430 2960 4440
rect 3400 4430 3840 4440
rect 3960 4430 4600 4440
rect 4680 4430 5280 4440
rect 6240 4430 6320 4440
rect 7440 4430 7760 4440
rect 8280 4430 8840 4440
rect 9240 4430 9560 4440
rect 9960 4430 9990 4440
rect 480 4420 520 4430
rect 600 4420 1040 4430
rect 1160 4420 2800 4430
rect 2880 4420 2960 4430
rect 3400 4420 3840 4430
rect 3960 4420 4600 4430
rect 4680 4420 5280 4430
rect 6240 4420 6320 4430
rect 7440 4420 7760 4430
rect 8280 4420 8840 4430
rect 9240 4420 9560 4430
rect 9960 4420 9990 4430
rect 280 4410 320 4420
rect 400 4410 2640 4420
rect 2680 4410 2800 4420
rect 2880 4410 2960 4420
rect 3400 4410 3800 4420
rect 3960 4410 4240 4420
rect 4320 4410 4600 4420
rect 4760 4410 4800 4420
rect 4880 4410 5280 4420
rect 7440 4410 7800 4420
rect 8080 4410 8120 4420
rect 8160 4410 8640 4420
rect 8720 4410 8840 4420
rect 9200 4410 9520 4420
rect 9920 4410 9990 4420
rect 280 4400 320 4410
rect 400 4400 2640 4410
rect 2680 4400 2800 4410
rect 2880 4400 2960 4410
rect 3400 4400 3800 4410
rect 3960 4400 4240 4410
rect 4320 4400 4600 4410
rect 4760 4400 4800 4410
rect 4880 4400 5280 4410
rect 7440 4400 7800 4410
rect 8080 4400 8120 4410
rect 8160 4400 8640 4410
rect 8720 4400 8840 4410
rect 9200 4400 9520 4410
rect 9920 4400 9990 4410
rect 280 4390 320 4400
rect 400 4390 2640 4400
rect 2680 4390 2800 4400
rect 2880 4390 2960 4400
rect 3400 4390 3800 4400
rect 3960 4390 4240 4400
rect 4320 4390 4600 4400
rect 4760 4390 4800 4400
rect 4880 4390 5280 4400
rect 7440 4390 7800 4400
rect 8080 4390 8120 4400
rect 8160 4390 8640 4400
rect 8720 4390 8840 4400
rect 9200 4390 9520 4400
rect 9920 4390 9990 4400
rect 280 4380 320 4390
rect 400 4380 2640 4390
rect 2680 4380 2800 4390
rect 2880 4380 2960 4390
rect 3400 4380 3800 4390
rect 3960 4380 4240 4390
rect 4320 4380 4600 4390
rect 4760 4380 4800 4390
rect 4880 4380 5280 4390
rect 7440 4380 7800 4390
rect 8080 4380 8120 4390
rect 8160 4380 8640 4390
rect 8720 4380 8840 4390
rect 9200 4380 9520 4390
rect 9920 4380 9990 4390
rect 240 4370 2800 4380
rect 2880 4370 2920 4380
rect 3120 4370 3160 4380
rect 3360 4370 3840 4380
rect 3920 4370 4280 4380
rect 4320 4370 4560 4380
rect 4920 4370 5320 4380
rect 7440 4370 7800 4380
rect 7880 4370 8120 4380
rect 8200 4370 8480 4380
rect 8760 4370 8840 4380
rect 9200 4370 9480 4380
rect 240 4360 2800 4370
rect 2880 4360 2920 4370
rect 3120 4360 3160 4370
rect 3360 4360 3840 4370
rect 3920 4360 4280 4370
rect 4320 4360 4560 4370
rect 4920 4360 5320 4370
rect 7440 4360 7800 4370
rect 7880 4360 8120 4370
rect 8200 4360 8480 4370
rect 8760 4360 8840 4370
rect 9200 4360 9480 4370
rect 240 4350 2800 4360
rect 2880 4350 2920 4360
rect 3120 4350 3160 4360
rect 3360 4350 3840 4360
rect 3920 4350 4280 4360
rect 4320 4350 4560 4360
rect 4920 4350 5320 4360
rect 7440 4350 7800 4360
rect 7880 4350 8120 4360
rect 8200 4350 8480 4360
rect 8760 4350 8840 4360
rect 9200 4350 9480 4360
rect 240 4340 2800 4350
rect 2880 4340 2920 4350
rect 3120 4340 3160 4350
rect 3360 4340 3840 4350
rect 3920 4340 4280 4350
rect 4320 4340 4560 4350
rect 4920 4340 5320 4350
rect 7440 4340 7800 4350
rect 7880 4340 8120 4350
rect 8200 4340 8480 4350
rect 8760 4340 8840 4350
rect 9200 4340 9480 4350
rect 240 4330 2800 4340
rect 2880 4330 2920 4340
rect 3040 4330 3080 4340
rect 3320 4330 4160 4340
rect 4280 4330 4520 4340
rect 4960 4330 5320 4340
rect 7400 4330 8160 4340
rect 8200 4330 8440 4340
rect 8760 4330 8840 4340
rect 9200 4330 9440 4340
rect 240 4320 2800 4330
rect 2880 4320 2920 4330
rect 3040 4320 3080 4330
rect 3320 4320 4160 4330
rect 4280 4320 4520 4330
rect 4960 4320 5320 4330
rect 7400 4320 8160 4330
rect 8200 4320 8440 4330
rect 8760 4320 8840 4330
rect 9200 4320 9440 4330
rect 240 4310 2800 4320
rect 2880 4310 2920 4320
rect 3040 4310 3080 4320
rect 3320 4310 4160 4320
rect 4280 4310 4520 4320
rect 4960 4310 5320 4320
rect 7400 4310 8160 4320
rect 8200 4310 8440 4320
rect 8760 4310 8840 4320
rect 9200 4310 9440 4320
rect 240 4300 2800 4310
rect 2880 4300 2920 4310
rect 3040 4300 3080 4310
rect 3320 4300 4160 4310
rect 4280 4300 4520 4310
rect 4960 4300 5320 4310
rect 7400 4300 8160 4310
rect 8200 4300 8440 4310
rect 8760 4300 8840 4310
rect 9200 4300 9440 4310
rect 80 4290 2800 4300
rect 3320 4290 4120 4300
rect 4320 4290 4520 4300
rect 5000 4290 5320 4300
rect 7240 4290 8160 4300
rect 8200 4290 8440 4300
rect 8760 4290 8840 4300
rect 9200 4290 9400 4300
rect 80 4280 2800 4290
rect 3320 4280 4120 4290
rect 4320 4280 4520 4290
rect 5000 4280 5320 4290
rect 7240 4280 8160 4290
rect 8200 4280 8440 4290
rect 8760 4280 8840 4290
rect 9200 4280 9400 4290
rect 80 4270 2800 4280
rect 3320 4270 4120 4280
rect 4320 4270 4520 4280
rect 5000 4270 5320 4280
rect 7240 4270 8160 4280
rect 8200 4270 8440 4280
rect 8760 4270 8840 4280
rect 9200 4270 9400 4280
rect 80 4260 2800 4270
rect 3320 4260 4120 4270
rect 4320 4260 4520 4270
rect 5000 4260 5320 4270
rect 7240 4260 8160 4270
rect 8200 4260 8440 4270
rect 8760 4260 8840 4270
rect 9200 4260 9400 4270
rect 120 4250 2800 4260
rect 3280 4250 4120 4260
rect 4360 4250 4480 4260
rect 5000 4250 5360 4260
rect 7480 4250 8160 4260
rect 8200 4250 8440 4260
rect 8560 4250 8840 4260
rect 9200 4250 9360 4260
rect 120 4240 2800 4250
rect 3280 4240 4120 4250
rect 4360 4240 4480 4250
rect 5000 4240 5360 4250
rect 7480 4240 8160 4250
rect 8200 4240 8440 4250
rect 8560 4240 8840 4250
rect 9200 4240 9360 4250
rect 120 4230 2800 4240
rect 3280 4230 4120 4240
rect 4360 4230 4480 4240
rect 5000 4230 5360 4240
rect 7480 4230 8160 4240
rect 8200 4230 8440 4240
rect 8560 4230 8840 4240
rect 9200 4230 9360 4240
rect 120 4220 2800 4230
rect 3280 4220 4120 4230
rect 4360 4220 4480 4230
rect 5000 4220 5360 4230
rect 7480 4220 8160 4230
rect 8200 4220 8440 4230
rect 8560 4220 8840 4230
rect 9200 4220 9360 4230
rect 120 4210 2560 4220
rect 2600 4210 2760 4220
rect 2800 4210 2840 4220
rect 2960 4210 3000 4220
rect 3280 4210 4080 4220
rect 5040 4210 5360 4220
rect 7480 4210 8160 4220
rect 8200 4210 8800 4220
rect 120 4200 2560 4210
rect 2600 4200 2760 4210
rect 2800 4200 2840 4210
rect 2960 4200 3000 4210
rect 3280 4200 4080 4210
rect 5040 4200 5360 4210
rect 7480 4200 8160 4210
rect 8200 4200 8800 4210
rect 120 4190 2560 4200
rect 2600 4190 2760 4200
rect 2800 4190 2840 4200
rect 2960 4190 3000 4200
rect 3280 4190 4080 4200
rect 5040 4190 5360 4200
rect 7480 4190 8160 4200
rect 8200 4190 8800 4200
rect 120 4180 2560 4190
rect 2600 4180 2760 4190
rect 2800 4180 2840 4190
rect 2960 4180 3000 4190
rect 3280 4180 4080 4190
rect 5040 4180 5360 4190
rect 7480 4180 8160 4190
rect 8200 4180 8800 4190
rect 160 4170 2560 4180
rect 3280 4170 4080 4180
rect 5080 4170 5400 4180
rect 5520 4170 5560 4180
rect 7280 4170 7320 4180
rect 7480 4170 8800 4180
rect 160 4160 2560 4170
rect 3280 4160 4080 4170
rect 5080 4160 5400 4170
rect 5520 4160 5560 4170
rect 7280 4160 7320 4170
rect 7480 4160 8800 4170
rect 160 4150 2560 4160
rect 3280 4150 4080 4160
rect 5080 4150 5400 4160
rect 5520 4150 5560 4160
rect 7280 4150 7320 4160
rect 7480 4150 8800 4160
rect 160 4140 2560 4150
rect 3280 4140 4080 4150
rect 5080 4140 5400 4150
rect 5520 4140 5560 4150
rect 7280 4140 7320 4150
rect 7480 4140 8800 4150
rect 0 4130 80 4140
rect 160 4130 2600 4140
rect 2640 4130 2680 4140
rect 3280 4130 4040 4140
rect 4760 4130 4880 4140
rect 5120 4130 5440 4140
rect 5520 4130 5600 4140
rect 7280 4130 7400 4140
rect 7480 4130 8800 4140
rect 0 4120 80 4130
rect 160 4120 2600 4130
rect 2640 4120 2680 4130
rect 3280 4120 4040 4130
rect 4760 4120 4880 4130
rect 5120 4120 5440 4130
rect 5520 4120 5600 4130
rect 7280 4120 7400 4130
rect 7480 4120 8800 4130
rect 0 4110 80 4120
rect 160 4110 2600 4120
rect 2640 4110 2680 4120
rect 3280 4110 4040 4120
rect 4760 4110 4880 4120
rect 5120 4110 5440 4120
rect 5520 4110 5600 4120
rect 7280 4110 7400 4120
rect 7480 4110 8800 4120
rect 0 4100 80 4110
rect 160 4100 2600 4110
rect 2640 4100 2680 4110
rect 3280 4100 4040 4110
rect 4760 4100 4880 4110
rect 5120 4100 5440 4110
rect 5520 4100 5600 4110
rect 7280 4100 7400 4110
rect 7480 4100 8800 4110
rect 0 4090 120 4100
rect 160 4090 2600 4100
rect 3280 4090 4040 4100
rect 4680 4090 4800 4100
rect 5160 4090 5400 4100
rect 5520 4090 5640 4100
rect 7240 4090 7480 4100
rect 7640 4090 8760 4100
rect 0 4080 120 4090
rect 160 4080 2600 4090
rect 3280 4080 4040 4090
rect 4680 4080 4800 4090
rect 5160 4080 5400 4090
rect 5520 4080 5640 4090
rect 7240 4080 7480 4090
rect 7640 4080 8760 4090
rect 0 4070 120 4080
rect 160 4070 2600 4080
rect 3280 4070 4040 4080
rect 4680 4070 4800 4080
rect 5160 4070 5400 4080
rect 5520 4070 5640 4080
rect 7240 4070 7480 4080
rect 7640 4070 8760 4080
rect 0 4060 120 4070
rect 160 4060 2600 4070
rect 3280 4060 4040 4070
rect 4680 4060 4800 4070
rect 5160 4060 5400 4070
rect 5520 4060 5640 4070
rect 7240 4060 7480 4070
rect 7640 4060 8760 4070
rect 0 4050 2600 4060
rect 3280 4050 4000 4060
rect 4640 4050 4760 4060
rect 5160 4050 5400 4060
rect 5520 4050 5680 4060
rect 7240 4050 7600 4060
rect 7760 4050 8520 4060
rect 8680 4050 8760 4060
rect 0 4040 2600 4050
rect 3280 4040 4000 4050
rect 4640 4040 4760 4050
rect 5160 4040 5400 4050
rect 5520 4040 5680 4050
rect 7240 4040 7600 4050
rect 7760 4040 8520 4050
rect 8680 4040 8760 4050
rect 0 4030 2600 4040
rect 3280 4030 4000 4040
rect 4640 4030 4760 4040
rect 5160 4030 5400 4040
rect 5520 4030 5680 4040
rect 7240 4030 7600 4040
rect 7760 4030 8520 4040
rect 8680 4030 8760 4040
rect 0 4020 2600 4030
rect 3280 4020 4000 4030
rect 4640 4020 4760 4030
rect 5160 4020 5400 4030
rect 5520 4020 5680 4030
rect 7240 4020 7600 4030
rect 7760 4020 8520 4030
rect 8680 4020 8760 4030
rect 0 4010 2600 4020
rect 3280 4010 4000 4020
rect 5160 4010 5400 4020
rect 5520 4010 5720 4020
rect 7200 4010 7720 4020
rect 7840 4010 8320 4020
rect 0 4000 2600 4010
rect 3280 4000 4000 4010
rect 5160 4000 5400 4010
rect 5520 4000 5720 4010
rect 7200 4000 7720 4010
rect 7840 4000 8320 4010
rect 0 3990 2600 4000
rect 3280 3990 4000 4000
rect 5160 3990 5400 4000
rect 5520 3990 5720 4000
rect 7200 3990 7720 4000
rect 7840 3990 8320 4000
rect 0 3980 2600 3990
rect 3280 3980 4000 3990
rect 5160 3980 5400 3990
rect 5520 3980 5720 3990
rect 7200 3980 7720 3990
rect 7840 3980 8320 3990
rect 0 3970 2600 3980
rect 3280 3970 3920 3980
rect 5200 3970 5400 3980
rect 5520 3970 5800 3980
rect 7200 3970 7840 3980
rect 7960 3970 8120 3980
rect 0 3960 2600 3970
rect 3280 3960 3920 3970
rect 5200 3960 5400 3970
rect 5520 3960 5800 3970
rect 7200 3960 7840 3970
rect 7960 3960 8120 3970
rect 0 3950 2600 3960
rect 3280 3950 3920 3960
rect 5200 3950 5400 3960
rect 5520 3950 5800 3960
rect 7200 3950 7840 3960
rect 7960 3950 8120 3960
rect 0 3940 2600 3950
rect 3280 3940 3920 3950
rect 5200 3940 5400 3950
rect 5520 3940 5800 3950
rect 7200 3940 7840 3950
rect 7960 3940 8120 3950
rect 0 3930 2600 3940
rect 3280 3930 3880 3940
rect 5240 3930 5400 3940
rect 5480 3930 6040 3940
rect 7160 3930 7920 3940
rect 0 3920 2600 3930
rect 3280 3920 3880 3930
rect 5240 3920 5400 3930
rect 5480 3920 6040 3930
rect 7160 3920 7920 3930
rect 0 3910 2600 3920
rect 3280 3910 3880 3920
rect 5240 3910 5400 3920
rect 5480 3910 6040 3920
rect 7160 3910 7920 3920
rect 0 3900 2600 3910
rect 3280 3900 3880 3910
rect 5240 3900 5400 3910
rect 5480 3900 6040 3910
rect 7160 3900 7920 3910
rect 0 3890 2520 3900
rect 3280 3890 3880 3900
rect 5240 3890 6000 3900
rect 7160 3890 7960 3900
rect 8080 3890 8200 3900
rect 0 3880 2520 3890
rect 3280 3880 3880 3890
rect 5240 3880 6000 3890
rect 7160 3880 7960 3890
rect 8080 3880 8200 3890
rect 0 3870 2520 3880
rect 3280 3870 3880 3880
rect 5240 3870 6000 3880
rect 7160 3870 7960 3880
rect 8080 3870 8200 3880
rect 0 3860 2520 3870
rect 3280 3860 3880 3870
rect 5240 3860 6000 3870
rect 7160 3860 7960 3870
rect 8080 3860 8200 3870
rect 0 3850 2240 3860
rect 2280 3850 2400 3860
rect 2480 3850 2560 3860
rect 3280 3850 3840 3860
rect 4160 3850 4240 3860
rect 5280 3850 5960 3860
rect 7120 3850 8000 3860
rect 8120 3850 8160 3860
rect 9640 3850 9680 3860
rect 0 3840 2240 3850
rect 2280 3840 2400 3850
rect 2480 3840 2560 3850
rect 3280 3840 3840 3850
rect 4160 3840 4240 3850
rect 5280 3840 5960 3850
rect 7120 3840 8000 3850
rect 8120 3840 8160 3850
rect 9640 3840 9680 3850
rect 0 3830 2240 3840
rect 2280 3830 2400 3840
rect 2480 3830 2560 3840
rect 3280 3830 3840 3840
rect 4160 3830 4240 3840
rect 5280 3830 5960 3840
rect 7120 3830 8000 3840
rect 8120 3830 8160 3840
rect 9640 3830 9680 3840
rect 0 3820 2240 3830
rect 2280 3820 2400 3830
rect 2480 3820 2560 3830
rect 3280 3820 3840 3830
rect 4160 3820 4240 3830
rect 5280 3820 5960 3830
rect 7120 3820 8000 3830
rect 8120 3820 8160 3830
rect 9640 3820 9680 3830
rect 0 3810 2600 3820
rect 3280 3810 3840 3820
rect 4080 3810 4240 3820
rect 5280 3810 5960 3820
rect 7120 3810 8080 3820
rect 9640 3810 9680 3820
rect 0 3800 2600 3810
rect 3280 3800 3840 3810
rect 4080 3800 4240 3810
rect 5280 3800 5960 3810
rect 7120 3800 8080 3810
rect 9640 3800 9680 3810
rect 0 3790 2600 3800
rect 3280 3790 3840 3800
rect 4080 3790 4240 3800
rect 5280 3790 5960 3800
rect 7120 3790 8080 3800
rect 9640 3790 9680 3800
rect 0 3780 2600 3790
rect 3280 3780 3840 3790
rect 4080 3780 4240 3790
rect 5280 3780 5960 3790
rect 7120 3780 8080 3790
rect 9640 3780 9680 3790
rect 0 3770 1640 3780
rect 1720 3770 2560 3780
rect 2600 3770 2640 3780
rect 3320 3770 3880 3780
rect 4040 3770 4080 3780
rect 5320 3770 6000 3780
rect 7080 3770 8120 3780
rect 0 3760 1640 3770
rect 1720 3760 2560 3770
rect 2600 3760 2640 3770
rect 3320 3760 3880 3770
rect 4040 3760 4080 3770
rect 5320 3760 6000 3770
rect 7080 3760 8120 3770
rect 0 3750 1640 3760
rect 1720 3750 2560 3760
rect 2600 3750 2640 3760
rect 3320 3750 3880 3760
rect 4040 3750 4080 3760
rect 5320 3750 6000 3760
rect 7080 3750 8120 3760
rect 0 3740 1640 3750
rect 1720 3740 2560 3750
rect 2600 3740 2640 3750
rect 3320 3740 3880 3750
rect 4040 3740 4080 3750
rect 5320 3740 6000 3750
rect 7080 3740 8120 3750
rect 0 3730 1600 3740
rect 1720 3730 2760 3740
rect 3320 3730 3880 3740
rect 5320 3730 6040 3740
rect 7040 3730 8160 3740
rect 0 3720 1600 3730
rect 1720 3720 2760 3730
rect 3320 3720 3880 3730
rect 5320 3720 6040 3730
rect 7040 3720 8160 3730
rect 0 3710 1600 3720
rect 1720 3710 2760 3720
rect 3320 3710 3880 3720
rect 5320 3710 6040 3720
rect 7040 3710 8160 3720
rect 0 3700 1600 3710
rect 1720 3700 2760 3710
rect 3320 3700 3880 3710
rect 5320 3700 6040 3710
rect 7040 3700 8160 3710
rect 40 3690 1600 3700
rect 1720 3690 2880 3700
rect 2960 3690 3000 3700
rect 3360 3690 3880 3700
rect 5320 3690 6080 3700
rect 7040 3690 8200 3700
rect 40 3680 1600 3690
rect 1720 3680 2880 3690
rect 2960 3680 3000 3690
rect 3360 3680 3880 3690
rect 5320 3680 6080 3690
rect 7040 3680 8200 3690
rect 40 3670 1600 3680
rect 1720 3670 2880 3680
rect 2960 3670 3000 3680
rect 3360 3670 3880 3680
rect 5320 3670 6080 3680
rect 7040 3670 8200 3680
rect 40 3660 1600 3670
rect 1720 3660 2880 3670
rect 2960 3660 3000 3670
rect 3360 3660 3880 3670
rect 5320 3660 6080 3670
rect 7040 3660 8200 3670
rect 0 3650 1680 3660
rect 1720 3650 3080 3660
rect 3360 3650 3920 3660
rect 5360 3650 6160 3660
rect 7000 3650 8200 3660
rect 8440 3650 8480 3660
rect 0 3640 1680 3650
rect 1720 3640 3080 3650
rect 3360 3640 3920 3650
rect 5360 3640 6160 3650
rect 7000 3640 8200 3650
rect 8440 3640 8480 3650
rect 0 3630 1680 3640
rect 1720 3630 3080 3640
rect 3360 3630 3920 3640
rect 5360 3630 6160 3640
rect 7000 3630 8200 3640
rect 8440 3630 8480 3640
rect 0 3620 1680 3630
rect 1720 3620 3080 3630
rect 3360 3620 3920 3630
rect 5360 3620 6160 3630
rect 7000 3620 8200 3630
rect 8440 3620 8480 3630
rect 0 3610 1680 3620
rect 1720 3610 3200 3620
rect 3400 3610 3920 3620
rect 5360 3610 6160 3620
rect 6960 3610 8240 3620
rect 8440 3610 8480 3620
rect 0 3600 1680 3610
rect 1720 3600 3200 3610
rect 3400 3600 3920 3610
rect 5360 3600 6160 3610
rect 6960 3600 8240 3610
rect 8440 3600 8480 3610
rect 0 3590 1680 3600
rect 1720 3590 3200 3600
rect 3400 3590 3920 3600
rect 5360 3590 6160 3600
rect 6960 3590 8240 3600
rect 8440 3590 8480 3600
rect 0 3580 1680 3590
rect 1720 3580 3200 3590
rect 3400 3580 3920 3590
rect 5360 3580 6160 3590
rect 6960 3580 8240 3590
rect 8440 3580 8480 3590
rect 0 3570 1440 3580
rect 1480 3570 1680 3580
rect 1720 3570 3240 3580
rect 3400 3570 3880 3580
rect 5360 3570 6160 3580
rect 6920 3570 8280 3580
rect 0 3560 1440 3570
rect 1480 3560 1680 3570
rect 1720 3560 3240 3570
rect 3400 3560 3880 3570
rect 5360 3560 6160 3570
rect 6920 3560 8280 3570
rect 0 3550 1440 3560
rect 1480 3550 1680 3560
rect 1720 3550 3240 3560
rect 3400 3550 3880 3560
rect 5360 3550 6160 3560
rect 6920 3550 8280 3560
rect 0 3540 1440 3550
rect 1480 3540 1680 3550
rect 1720 3540 3240 3550
rect 3400 3540 3880 3550
rect 5360 3540 6160 3550
rect 6920 3540 8280 3550
rect 0 3530 1440 3540
rect 1480 3530 2520 3540
rect 2600 3530 3280 3540
rect 3440 3530 3920 3540
rect 5360 3530 6160 3540
rect 6880 3530 8320 3540
rect 0 3520 1440 3530
rect 1480 3520 2520 3530
rect 2600 3520 3280 3530
rect 3440 3520 3920 3530
rect 5360 3520 6160 3530
rect 6880 3520 8320 3530
rect 0 3510 1440 3520
rect 1480 3510 2520 3520
rect 2600 3510 3280 3520
rect 3440 3510 3920 3520
rect 5360 3510 6160 3520
rect 6880 3510 8320 3520
rect 0 3500 1440 3510
rect 1480 3500 2520 3510
rect 2600 3500 3280 3510
rect 3440 3500 3920 3510
rect 5360 3500 6160 3510
rect 6880 3500 8320 3510
rect 0 3490 1400 3500
rect 1480 3490 2360 3500
rect 2840 3490 3320 3500
rect 3440 3490 3920 3500
rect 5360 3490 6160 3500
rect 6880 3490 8360 3500
rect 0 3480 1400 3490
rect 1480 3480 2360 3490
rect 2840 3480 3320 3490
rect 3440 3480 3920 3490
rect 5360 3480 6160 3490
rect 6880 3480 8360 3490
rect 0 3470 1400 3480
rect 1480 3470 2360 3480
rect 2840 3470 3320 3480
rect 3440 3470 3920 3480
rect 5360 3470 6160 3480
rect 6880 3470 8360 3480
rect 0 3460 1400 3470
rect 1480 3460 2360 3470
rect 2840 3460 3320 3470
rect 3440 3460 3920 3470
rect 5360 3460 6160 3470
rect 6880 3460 8360 3470
rect 0 3450 1400 3460
rect 1440 3450 2240 3460
rect 2960 3450 3360 3460
rect 3440 3450 3920 3460
rect 4920 3450 5000 3460
rect 5360 3450 5840 3460
rect 6000 3450 6120 3460
rect 6840 3450 8440 3460
rect 0 3440 1400 3450
rect 1440 3440 2240 3450
rect 2960 3440 3360 3450
rect 3440 3440 3920 3450
rect 4920 3440 5000 3450
rect 5360 3440 5840 3450
rect 6000 3440 6120 3450
rect 6840 3440 8440 3450
rect 0 3430 1400 3440
rect 1440 3430 2240 3440
rect 2960 3430 3360 3440
rect 3440 3430 3920 3440
rect 4920 3430 5000 3440
rect 5360 3430 5840 3440
rect 6000 3430 6120 3440
rect 6840 3430 8440 3440
rect 0 3420 1400 3430
rect 1440 3420 2240 3430
rect 2960 3420 3360 3430
rect 3440 3420 3920 3430
rect 4920 3420 5000 3430
rect 5360 3420 5840 3430
rect 6000 3420 6120 3430
rect 6840 3420 8440 3430
rect 0 3410 1360 3420
rect 1440 3410 2200 3420
rect 3040 3410 3960 3420
rect 5360 3410 5680 3420
rect 5720 3410 5840 3420
rect 6080 3410 6120 3420
rect 6800 3410 8480 3420
rect 0 3400 1360 3410
rect 1440 3400 2200 3410
rect 3040 3400 3960 3410
rect 5360 3400 5680 3410
rect 5720 3400 5840 3410
rect 6080 3400 6120 3410
rect 6800 3400 8480 3410
rect 0 3390 1360 3400
rect 1440 3390 2200 3400
rect 3040 3390 3960 3400
rect 5360 3390 5680 3400
rect 5720 3390 5840 3400
rect 6080 3390 6120 3400
rect 6800 3390 8480 3400
rect 0 3380 1360 3390
rect 1440 3380 2200 3390
rect 3040 3380 3960 3390
rect 5360 3380 5680 3390
rect 5720 3380 5840 3390
rect 6080 3380 6120 3390
rect 6800 3380 8480 3390
rect 0 3370 1360 3380
rect 1440 3370 2120 3380
rect 3080 3370 3480 3380
rect 3600 3370 3960 3380
rect 4800 3370 4840 3380
rect 5360 3370 5640 3380
rect 5760 3370 5840 3380
rect 6080 3370 6120 3380
rect 6720 3370 8480 3380
rect 0 3360 1360 3370
rect 1440 3360 2120 3370
rect 3080 3360 3480 3370
rect 3600 3360 3960 3370
rect 4800 3360 4840 3370
rect 5360 3360 5640 3370
rect 5760 3360 5840 3370
rect 6080 3360 6120 3370
rect 6720 3360 8480 3370
rect 0 3350 1360 3360
rect 1440 3350 2120 3360
rect 3080 3350 3480 3360
rect 3600 3350 3960 3360
rect 4800 3350 4840 3360
rect 5360 3350 5640 3360
rect 5760 3350 5840 3360
rect 6080 3350 6120 3360
rect 6720 3350 8480 3360
rect 0 3340 1360 3350
rect 1440 3340 2120 3350
rect 3080 3340 3480 3350
rect 3600 3340 3960 3350
rect 4800 3340 4840 3350
rect 5360 3340 5640 3350
rect 5760 3340 5840 3350
rect 6080 3340 6120 3350
rect 6720 3340 8480 3350
rect 0 3330 1320 3340
rect 1400 3330 2080 3340
rect 3120 3330 3480 3340
rect 3600 3330 3960 3340
rect 5320 3330 5600 3340
rect 5800 3330 5840 3340
rect 6680 3330 8480 3340
rect 0 3320 1320 3330
rect 1400 3320 2080 3330
rect 3120 3320 3480 3330
rect 3600 3320 3960 3330
rect 5320 3320 5600 3330
rect 5800 3320 5840 3330
rect 6680 3320 8480 3330
rect 0 3310 1320 3320
rect 1400 3310 2080 3320
rect 3120 3310 3480 3320
rect 3600 3310 3960 3320
rect 5320 3310 5600 3320
rect 5800 3310 5840 3320
rect 6680 3310 8480 3320
rect 0 3300 1320 3310
rect 1400 3300 2080 3310
rect 3120 3300 3480 3310
rect 3600 3300 3960 3310
rect 5320 3300 5600 3310
rect 5800 3300 5840 3310
rect 6680 3300 8480 3310
rect 0 3290 1320 3300
rect 1400 3290 2080 3300
rect 3160 3290 3520 3300
rect 3600 3290 4000 3300
rect 4600 3290 4680 3300
rect 5320 3290 5600 3300
rect 6680 3290 8440 3300
rect 0 3280 1320 3290
rect 1400 3280 2080 3290
rect 3160 3280 3520 3290
rect 3600 3280 4000 3290
rect 4600 3280 4680 3290
rect 5320 3280 5600 3290
rect 6680 3280 8440 3290
rect 0 3270 1320 3280
rect 1400 3270 2080 3280
rect 3160 3270 3520 3280
rect 3600 3270 4000 3280
rect 4600 3270 4680 3280
rect 5320 3270 5600 3280
rect 6680 3270 8440 3280
rect 0 3260 1320 3270
rect 1400 3260 2080 3270
rect 3160 3260 3520 3270
rect 3600 3260 4000 3270
rect 4600 3260 4680 3270
rect 5320 3260 5600 3270
rect 6680 3260 8440 3270
rect 0 3250 1280 3260
rect 1400 3250 2040 3260
rect 3160 3250 3560 3260
rect 3640 3250 4040 3260
rect 4440 3250 4600 3260
rect 5320 3250 5640 3260
rect 6680 3250 8440 3260
rect 0 3240 1280 3250
rect 1400 3240 2040 3250
rect 3160 3240 3560 3250
rect 3640 3240 4040 3250
rect 4440 3240 4600 3250
rect 5320 3240 5640 3250
rect 6680 3240 8440 3250
rect 0 3230 1280 3240
rect 1400 3230 2040 3240
rect 3160 3230 3560 3240
rect 3640 3230 4040 3240
rect 4440 3230 4600 3240
rect 5320 3230 5640 3240
rect 6680 3230 8440 3240
rect 0 3220 1280 3230
rect 1400 3220 2040 3230
rect 3160 3220 3560 3230
rect 3640 3220 4040 3230
rect 4440 3220 4600 3230
rect 5320 3220 5640 3230
rect 6680 3220 8440 3230
rect 0 3210 1280 3220
rect 1360 3210 2040 3220
rect 3200 3210 3560 3220
rect 3600 3210 4040 3220
rect 4360 3210 4480 3220
rect 5320 3210 5680 3220
rect 6480 3210 6560 3220
rect 6680 3210 8400 3220
rect 9080 3210 9120 3220
rect 0 3200 1280 3210
rect 1360 3200 2040 3210
rect 3200 3200 3560 3210
rect 3600 3200 4040 3210
rect 4360 3200 4480 3210
rect 5320 3200 5680 3210
rect 6480 3200 6560 3210
rect 6680 3200 8400 3210
rect 9080 3200 9120 3210
rect 0 3190 1280 3200
rect 1360 3190 2040 3200
rect 3200 3190 3560 3200
rect 3600 3190 4040 3200
rect 4360 3190 4480 3200
rect 5320 3190 5680 3200
rect 6480 3190 6560 3200
rect 6680 3190 8400 3200
rect 9080 3190 9120 3200
rect 0 3180 1280 3190
rect 1360 3180 2040 3190
rect 3200 3180 3560 3190
rect 3600 3180 4040 3190
rect 4360 3180 4480 3190
rect 5320 3180 5680 3190
rect 6480 3180 6560 3190
rect 6680 3180 8400 3190
rect 9080 3180 9120 3190
rect 0 3170 1240 3180
rect 1360 3170 2040 3180
rect 3200 3170 4080 3180
rect 5280 3170 5720 3180
rect 6360 3170 6560 3180
rect 6640 3170 8400 3180
rect 9120 3170 9240 3180
rect 0 3160 1240 3170
rect 1360 3160 2040 3170
rect 3200 3160 4080 3170
rect 5280 3160 5720 3170
rect 6360 3160 6560 3170
rect 6640 3160 8400 3170
rect 9120 3160 9240 3170
rect 0 3150 1240 3160
rect 1360 3150 2040 3160
rect 3200 3150 4080 3160
rect 5280 3150 5720 3160
rect 6360 3150 6560 3160
rect 6640 3150 8400 3160
rect 9120 3150 9240 3160
rect 0 3140 1240 3150
rect 1360 3140 2040 3150
rect 3200 3140 4080 3150
rect 5280 3140 5720 3150
rect 6360 3140 6560 3150
rect 6640 3140 8400 3150
rect 9120 3140 9240 3150
rect 0 3130 1240 3140
rect 1360 3130 2000 3140
rect 3200 3130 3760 3140
rect 3920 3130 4080 3140
rect 5280 3130 5880 3140
rect 6120 3130 6560 3140
rect 6640 3130 8360 3140
rect 9120 3130 9200 3140
rect 0 3120 1240 3130
rect 1360 3120 2000 3130
rect 3200 3120 3760 3130
rect 3920 3120 4080 3130
rect 5280 3120 5880 3130
rect 6120 3120 6560 3130
rect 6640 3120 8360 3130
rect 9120 3120 9200 3130
rect 0 3110 1240 3120
rect 1360 3110 2000 3120
rect 3200 3110 3760 3120
rect 3920 3110 4080 3120
rect 5280 3110 5880 3120
rect 6120 3110 6560 3120
rect 6640 3110 8360 3120
rect 9120 3110 9200 3120
rect 0 3100 1240 3110
rect 1360 3100 2000 3110
rect 3200 3100 3760 3110
rect 3920 3100 4080 3110
rect 5280 3100 5880 3110
rect 6120 3100 6560 3110
rect 6640 3100 8360 3110
rect 9120 3100 9200 3110
rect 0 3090 1240 3100
rect 1320 3090 2000 3100
rect 3200 3090 3760 3100
rect 4040 3090 4120 3100
rect 5240 3090 6560 3100
rect 6640 3090 8360 3100
rect 9120 3090 9200 3100
rect 0 3080 1240 3090
rect 1320 3080 2000 3090
rect 3200 3080 3760 3090
rect 4040 3080 4120 3090
rect 5240 3080 6560 3090
rect 6640 3080 8360 3090
rect 9120 3080 9200 3090
rect 0 3070 1240 3080
rect 1320 3070 2000 3080
rect 3200 3070 3760 3080
rect 4040 3070 4120 3080
rect 5240 3070 6560 3080
rect 6640 3070 8360 3080
rect 9120 3070 9200 3080
rect 0 3060 1240 3070
rect 1320 3060 2000 3070
rect 3200 3060 3760 3070
rect 4040 3060 4120 3070
rect 5240 3060 6560 3070
rect 6640 3060 8360 3070
rect 9120 3060 9200 3070
rect 0 3050 1200 3060
rect 1320 3050 2000 3060
rect 3200 3050 3720 3060
rect 4040 3050 4120 3060
rect 4640 3050 4720 3060
rect 5240 3050 6560 3060
rect 6640 3050 8320 3060
rect 9080 3050 9240 3060
rect 0 3040 1200 3050
rect 1320 3040 2000 3050
rect 3200 3040 3720 3050
rect 4040 3040 4120 3050
rect 4640 3040 4720 3050
rect 5240 3040 6560 3050
rect 6640 3040 8320 3050
rect 9080 3040 9240 3050
rect 0 3030 1200 3040
rect 1320 3030 2000 3040
rect 3200 3030 3720 3040
rect 4040 3030 4120 3040
rect 4640 3030 4720 3040
rect 5240 3030 6560 3040
rect 6640 3030 8320 3040
rect 9080 3030 9240 3040
rect 0 3020 1200 3030
rect 1320 3020 2000 3030
rect 3200 3020 3720 3030
rect 4040 3020 4120 3030
rect 4640 3020 4720 3030
rect 5240 3020 6560 3030
rect 6640 3020 8320 3030
rect 9080 3020 9240 3030
rect 0 3010 1200 3020
rect 1320 3010 2000 3020
rect 3200 3010 3720 3020
rect 4120 3010 4160 3020
rect 5240 3010 6520 3020
rect 6600 3010 8320 3020
rect 9080 3010 9120 3020
rect 0 3000 1200 3010
rect 1320 3000 2000 3010
rect 3200 3000 3720 3010
rect 4120 3000 4160 3010
rect 5240 3000 6520 3010
rect 6600 3000 8320 3010
rect 9080 3000 9120 3010
rect 0 2990 1200 3000
rect 1320 2990 2000 3000
rect 3200 2990 3720 3000
rect 4120 2990 4160 3000
rect 5240 2990 6520 3000
rect 6600 2990 8320 3000
rect 9080 2990 9120 3000
rect 0 2980 1200 2990
rect 1320 2980 2000 2990
rect 3200 2980 3720 2990
rect 4120 2980 4160 2990
rect 5240 2980 6520 2990
rect 6600 2980 8320 2990
rect 9080 2980 9120 2990
rect 0 2970 1160 2980
rect 1280 2970 2000 2980
rect 3200 2970 3840 2980
rect 4200 2970 4240 2980
rect 5200 2970 6520 2980
rect 6600 2970 8280 2980
rect 0 2960 1160 2970
rect 1280 2960 2000 2970
rect 3200 2960 3840 2970
rect 4200 2960 4240 2970
rect 5200 2960 6520 2970
rect 6600 2960 8280 2970
rect 0 2950 1160 2960
rect 1280 2950 2000 2960
rect 3200 2950 3840 2960
rect 4200 2950 4240 2960
rect 5200 2950 6520 2960
rect 6600 2950 8280 2960
rect 0 2940 1160 2950
rect 1280 2940 2000 2950
rect 3200 2940 3840 2950
rect 4200 2940 4240 2950
rect 5200 2940 6520 2950
rect 6600 2940 8280 2950
rect 0 2930 1160 2940
rect 1280 2930 2000 2940
rect 3160 2930 3800 2940
rect 4240 2930 4280 2940
rect 5200 2930 6520 2940
rect 6600 2930 8280 2940
rect 0 2920 1160 2930
rect 1280 2920 2000 2930
rect 3160 2920 3800 2930
rect 4240 2920 4280 2930
rect 5200 2920 6520 2930
rect 6600 2920 8280 2930
rect 0 2910 1160 2920
rect 1280 2910 2000 2920
rect 3160 2910 3800 2920
rect 4240 2910 4280 2920
rect 5200 2910 6520 2920
rect 6600 2910 8280 2920
rect 0 2900 1160 2910
rect 1280 2900 2000 2910
rect 3160 2900 3800 2910
rect 4240 2900 4280 2910
rect 5200 2900 6520 2910
rect 6600 2900 8280 2910
rect 0 2890 1160 2900
rect 1240 2890 2000 2900
rect 3160 2890 3880 2900
rect 3920 2890 3960 2900
rect 4280 2890 4360 2900
rect 5160 2890 6520 2900
rect 6600 2890 7400 2900
rect 7520 2890 8240 2900
rect 0 2880 1160 2890
rect 1240 2880 2000 2890
rect 3160 2880 3880 2890
rect 3920 2880 3960 2890
rect 4280 2880 4360 2890
rect 5160 2880 6520 2890
rect 6600 2880 7400 2890
rect 7520 2880 8240 2890
rect 0 2870 1160 2880
rect 1240 2870 2000 2880
rect 3160 2870 3880 2880
rect 3920 2870 3960 2880
rect 4280 2870 4360 2880
rect 5160 2870 6520 2880
rect 6600 2870 7400 2880
rect 7520 2870 8240 2880
rect 0 2860 1160 2870
rect 1240 2860 2000 2870
rect 3160 2860 3880 2870
rect 3920 2860 3960 2870
rect 4280 2860 4360 2870
rect 5160 2860 6520 2870
rect 6600 2860 7400 2870
rect 7520 2860 8240 2870
rect 0 2850 1120 2860
rect 1240 2850 1960 2860
rect 3160 2850 3880 2860
rect 4280 2850 4440 2860
rect 5160 2850 6520 2860
rect 6560 2850 7200 2860
rect 7560 2850 8200 2860
rect 0 2840 1120 2850
rect 1240 2840 1960 2850
rect 3160 2840 3880 2850
rect 4280 2840 4440 2850
rect 5160 2840 6520 2850
rect 6560 2840 7200 2850
rect 7560 2840 8200 2850
rect 0 2830 1120 2840
rect 1240 2830 1960 2840
rect 3160 2830 3880 2840
rect 4280 2830 4440 2840
rect 5160 2830 6520 2840
rect 6560 2830 7200 2840
rect 7560 2830 8200 2840
rect 0 2820 1120 2830
rect 1240 2820 1960 2830
rect 3160 2820 3880 2830
rect 4280 2820 4440 2830
rect 5160 2820 6520 2830
rect 6560 2820 7200 2830
rect 7560 2820 8200 2830
rect 0 2810 1120 2820
rect 1240 2810 1960 2820
rect 3160 2810 3960 2820
rect 4280 2810 4480 2820
rect 5200 2810 5720 2820
rect 6120 2810 6520 2820
rect 6560 2810 7120 2820
rect 7600 2810 8160 2820
rect 0 2800 1120 2810
rect 1240 2800 1960 2810
rect 3160 2800 3960 2810
rect 4280 2800 4480 2810
rect 5200 2800 5720 2810
rect 6120 2800 6520 2810
rect 6560 2800 7120 2810
rect 7600 2800 8160 2810
rect 0 2790 1120 2800
rect 1240 2790 1960 2800
rect 3160 2790 3960 2800
rect 4280 2790 4480 2800
rect 5200 2790 5720 2800
rect 6120 2790 6520 2800
rect 6560 2790 7120 2800
rect 7600 2790 8160 2800
rect 0 2780 1120 2790
rect 1240 2780 1960 2790
rect 3160 2780 3960 2790
rect 4280 2780 4480 2790
rect 5200 2780 5720 2790
rect 6120 2780 6520 2790
rect 6560 2780 7120 2790
rect 7600 2780 8160 2790
rect 0 2770 1080 2780
rect 1200 2770 1960 2780
rect 3160 2770 3880 2780
rect 4280 2770 4560 2780
rect 5200 2770 5520 2780
rect 6160 2770 6520 2780
rect 6560 2770 7080 2780
rect 7640 2770 8120 2780
rect 8760 2770 8800 2780
rect 0 2760 1080 2770
rect 1200 2760 1960 2770
rect 3160 2760 3880 2770
rect 4280 2760 4560 2770
rect 5200 2760 5520 2770
rect 6160 2760 6520 2770
rect 6560 2760 7080 2770
rect 7640 2760 8120 2770
rect 8760 2760 8800 2770
rect 0 2750 1080 2760
rect 1200 2750 1960 2760
rect 3160 2750 3880 2760
rect 4280 2750 4560 2760
rect 5200 2750 5520 2760
rect 6160 2750 6520 2760
rect 6560 2750 7080 2760
rect 7640 2750 8120 2760
rect 8760 2750 8800 2760
rect 0 2740 1080 2750
rect 1200 2740 1960 2750
rect 3160 2740 3880 2750
rect 4280 2740 4560 2750
rect 5200 2740 5520 2750
rect 6160 2740 6520 2750
rect 6560 2740 7080 2750
rect 7640 2740 8120 2750
rect 8760 2740 8800 2750
rect 0 2730 1080 2740
rect 1160 2730 1960 2740
rect 3160 2730 3880 2740
rect 4280 2730 4680 2740
rect 5200 2730 5240 2740
rect 5360 2730 5480 2740
rect 6160 2730 6520 2740
rect 6560 2730 7000 2740
rect 7680 2730 8120 2740
rect 0 2720 1080 2730
rect 1160 2720 1960 2730
rect 3160 2720 3880 2730
rect 4280 2720 4680 2730
rect 5200 2720 5240 2730
rect 5360 2720 5480 2730
rect 6160 2720 6520 2730
rect 6560 2720 7000 2730
rect 7680 2720 8120 2730
rect 0 2710 1080 2720
rect 1160 2710 1960 2720
rect 3160 2710 3880 2720
rect 4280 2710 4680 2720
rect 5200 2710 5240 2720
rect 5360 2710 5480 2720
rect 6160 2710 6520 2720
rect 6560 2710 7000 2720
rect 7680 2710 8120 2720
rect 0 2700 1080 2710
rect 1160 2700 1960 2710
rect 3160 2700 3880 2710
rect 4280 2700 4680 2710
rect 5200 2700 5240 2710
rect 5360 2700 5480 2710
rect 6160 2700 6520 2710
rect 6560 2700 7000 2710
rect 7680 2700 8120 2710
rect 0 2690 1040 2700
rect 1120 2690 1960 2700
rect 3160 2690 3880 2700
rect 4280 2690 4840 2700
rect 5160 2690 5200 2700
rect 5400 2690 5440 2700
rect 6200 2690 6520 2700
rect 6560 2690 6920 2700
rect 7720 2690 8080 2700
rect 0 2680 1040 2690
rect 1120 2680 1960 2690
rect 3160 2680 3880 2690
rect 4280 2680 4840 2690
rect 5160 2680 5200 2690
rect 5400 2680 5440 2690
rect 6200 2680 6520 2690
rect 6560 2680 6920 2690
rect 7720 2680 8080 2690
rect 0 2670 1040 2680
rect 1120 2670 1960 2680
rect 3160 2670 3880 2680
rect 4280 2670 4840 2680
rect 5160 2670 5200 2680
rect 5400 2670 5440 2680
rect 6200 2670 6520 2680
rect 6560 2670 6920 2680
rect 7720 2670 8080 2680
rect 0 2660 1040 2670
rect 1120 2660 1960 2670
rect 3160 2660 3880 2670
rect 4280 2660 4840 2670
rect 5160 2660 5200 2670
rect 5400 2660 5440 2670
rect 6200 2660 6520 2670
rect 6560 2660 6920 2670
rect 7720 2660 8080 2670
rect 0 2650 1040 2660
rect 1120 2650 1960 2660
rect 3160 2650 3880 2660
rect 4280 2650 4800 2660
rect 5360 2650 5400 2660
rect 6240 2650 6880 2660
rect 7720 2650 8040 2660
rect 9120 2650 9160 2660
rect 0 2640 1040 2650
rect 1120 2640 1960 2650
rect 3160 2640 3880 2650
rect 4280 2640 4800 2650
rect 5360 2640 5400 2650
rect 6240 2640 6880 2650
rect 7720 2640 8040 2650
rect 9120 2640 9160 2650
rect 0 2630 1040 2640
rect 1120 2630 1960 2640
rect 3160 2630 3880 2640
rect 4280 2630 4800 2640
rect 5360 2630 5400 2640
rect 6240 2630 6880 2640
rect 7720 2630 8040 2640
rect 9120 2630 9160 2640
rect 0 2620 1040 2630
rect 1120 2620 1960 2630
rect 3160 2620 3880 2630
rect 4280 2620 4800 2630
rect 5360 2620 5400 2630
rect 6240 2620 6880 2630
rect 7720 2620 8040 2630
rect 9120 2620 9160 2630
rect 0 2610 1000 2620
rect 1080 2610 1920 2620
rect 2280 2610 2360 2620
rect 2880 2610 3040 2620
rect 3120 2610 3880 2620
rect 4280 2610 4720 2620
rect 6280 2610 6840 2620
rect 7760 2610 8000 2620
rect 0 2600 1000 2610
rect 1080 2600 1920 2610
rect 2280 2600 2360 2610
rect 2880 2600 3040 2610
rect 3120 2600 3880 2610
rect 4280 2600 4720 2610
rect 6280 2600 6840 2610
rect 7760 2600 8000 2610
rect 0 2590 1000 2600
rect 1080 2590 1920 2600
rect 2280 2590 2360 2600
rect 2880 2590 3040 2600
rect 3120 2590 3880 2600
rect 4280 2590 4720 2600
rect 6280 2590 6840 2600
rect 7760 2590 8000 2600
rect 0 2580 1000 2590
rect 1080 2580 1920 2590
rect 2280 2580 2360 2590
rect 2880 2580 3040 2590
rect 3120 2580 3880 2590
rect 4280 2580 4720 2590
rect 6280 2580 6840 2590
rect 7760 2580 8000 2590
rect 0 2570 1000 2580
rect 1080 2570 1920 2580
rect 2040 2570 2320 2580
rect 2360 2570 2400 2580
rect 2840 2570 2880 2580
rect 2920 2570 3880 2580
rect 4280 2570 4520 2580
rect 4800 2570 4840 2580
rect 4880 2570 4920 2580
rect 6280 2570 6800 2580
rect 7800 2570 7960 2580
rect 0 2560 1000 2570
rect 1080 2560 1920 2570
rect 2040 2560 2320 2570
rect 2360 2560 2400 2570
rect 2840 2560 2880 2570
rect 2920 2560 3880 2570
rect 4280 2560 4520 2570
rect 4800 2560 4840 2570
rect 4880 2560 4920 2570
rect 6280 2560 6800 2570
rect 7800 2560 7960 2570
rect 0 2550 1000 2560
rect 1080 2550 1920 2560
rect 2040 2550 2320 2560
rect 2360 2550 2400 2560
rect 2840 2550 2880 2560
rect 2920 2550 3880 2560
rect 4280 2550 4520 2560
rect 4800 2550 4840 2560
rect 4880 2550 4920 2560
rect 6280 2550 6800 2560
rect 7800 2550 7960 2560
rect 0 2540 1000 2550
rect 1080 2540 1920 2550
rect 2040 2540 2320 2550
rect 2360 2540 2400 2550
rect 2840 2540 2880 2550
rect 2920 2540 3880 2550
rect 4280 2540 4520 2550
rect 4800 2540 4840 2550
rect 4880 2540 4920 2550
rect 6280 2540 6800 2550
rect 7800 2540 7960 2550
rect 0 2530 960 2540
rect 1040 2530 1920 2540
rect 3200 2530 3920 2540
rect 4160 2530 4680 2540
rect 6320 2530 6760 2540
rect 7800 2530 7880 2540
rect 0 2520 960 2530
rect 1040 2520 1920 2530
rect 3200 2520 3920 2530
rect 4160 2520 4680 2530
rect 6320 2520 6760 2530
rect 7800 2520 7880 2530
rect 0 2510 960 2520
rect 1040 2510 1920 2520
rect 3200 2510 3920 2520
rect 4160 2510 4680 2520
rect 6320 2510 6760 2520
rect 7800 2510 7880 2520
rect 0 2500 960 2510
rect 1040 2500 1920 2510
rect 3200 2500 3920 2510
rect 4160 2500 4680 2510
rect 6320 2500 6760 2510
rect 7800 2500 7880 2510
rect 0 2490 960 2500
rect 1040 2490 1880 2500
rect 3240 2490 3960 2500
rect 4120 2490 4600 2500
rect 6360 2490 6760 2500
rect 0 2480 960 2490
rect 1040 2480 1880 2490
rect 3240 2480 3960 2490
rect 4120 2480 4600 2490
rect 6360 2480 6760 2490
rect 0 2470 960 2480
rect 1040 2470 1880 2480
rect 3240 2470 3960 2480
rect 4120 2470 4600 2480
rect 6360 2470 6760 2480
rect 0 2460 960 2470
rect 1040 2460 1880 2470
rect 3240 2460 3960 2470
rect 4120 2460 4600 2470
rect 6360 2460 6760 2470
rect 0 2450 920 2460
rect 1040 2450 1880 2460
rect 3280 2450 3960 2460
rect 4080 2450 4560 2460
rect 6360 2450 6720 2460
rect 0 2440 920 2450
rect 1040 2440 1880 2450
rect 3280 2440 3960 2450
rect 4080 2440 4560 2450
rect 6360 2440 6720 2450
rect 0 2430 920 2440
rect 1040 2430 1880 2440
rect 3280 2430 3960 2440
rect 4080 2430 4560 2440
rect 6360 2430 6720 2440
rect 0 2420 920 2430
rect 1040 2420 1880 2430
rect 3280 2420 3960 2430
rect 4080 2420 4560 2430
rect 6360 2420 6720 2430
rect 0 2410 920 2420
rect 1040 2410 1880 2420
rect 3280 2410 4560 2420
rect 6400 2410 6720 2420
rect 0 2400 920 2410
rect 1040 2400 1880 2410
rect 3280 2400 4560 2410
rect 6400 2400 6720 2410
rect 0 2390 920 2400
rect 1040 2390 1880 2400
rect 3280 2390 4560 2400
rect 6400 2390 6720 2400
rect 0 2380 920 2390
rect 1040 2380 1880 2390
rect 3280 2380 4560 2390
rect 6400 2380 6720 2390
rect 0 2370 880 2380
rect 1000 2370 1880 2380
rect 3320 2370 4520 2380
rect 6400 2370 6720 2380
rect 9160 2370 9200 2380
rect 0 2360 880 2370
rect 1000 2360 1880 2370
rect 3320 2360 4520 2370
rect 6400 2360 6720 2370
rect 9160 2360 9200 2370
rect 0 2350 880 2360
rect 1000 2350 1880 2360
rect 3320 2350 4520 2360
rect 6400 2350 6720 2360
rect 9160 2350 9200 2360
rect 0 2340 880 2350
rect 1000 2340 1880 2350
rect 3320 2340 4520 2350
rect 6400 2340 6720 2350
rect 9160 2340 9200 2350
rect 0 2330 880 2340
rect 1000 2330 1840 2340
rect 3320 2330 4480 2340
rect 6440 2330 6720 2340
rect 8400 2330 8440 2340
rect 9160 2330 9200 2340
rect 0 2320 880 2330
rect 1000 2320 1840 2330
rect 3320 2320 4480 2330
rect 6440 2320 6720 2330
rect 8400 2320 8440 2330
rect 9160 2320 9200 2330
rect 0 2310 880 2320
rect 1000 2310 1840 2320
rect 3320 2310 4480 2320
rect 6440 2310 6720 2320
rect 8400 2310 8440 2320
rect 9160 2310 9200 2320
rect 0 2300 880 2310
rect 1000 2300 1840 2310
rect 3320 2300 4480 2310
rect 6440 2300 6720 2310
rect 8400 2300 8440 2310
rect 9160 2300 9200 2310
rect 0 2290 840 2300
rect 1000 2290 1840 2300
rect 3320 2290 4080 2300
rect 6440 2290 6720 2300
rect 7520 2290 7560 2300
rect 8360 2290 8560 2300
rect 9160 2290 9200 2300
rect 9640 2290 9720 2300
rect 0 2280 840 2290
rect 1000 2280 1840 2290
rect 3320 2280 4080 2290
rect 6440 2280 6720 2290
rect 7520 2280 7560 2290
rect 8360 2280 8560 2290
rect 9160 2280 9200 2290
rect 9640 2280 9720 2290
rect 0 2270 840 2280
rect 1000 2270 1840 2280
rect 3320 2270 4080 2280
rect 6440 2270 6720 2280
rect 7520 2270 7560 2280
rect 8360 2270 8560 2280
rect 9160 2270 9200 2280
rect 9640 2270 9720 2280
rect 0 2260 840 2270
rect 1000 2260 1840 2270
rect 3320 2260 4080 2270
rect 6440 2260 6720 2270
rect 7520 2260 7560 2270
rect 8360 2260 8560 2270
rect 9160 2260 9200 2270
rect 9640 2260 9720 2270
rect 0 2250 840 2260
rect 1000 2250 1840 2260
rect 3360 2250 4320 2260
rect 6480 2250 6720 2260
rect 7160 2250 7200 2260
rect 7520 2250 7600 2260
rect 8360 2250 8600 2260
rect 9160 2250 9240 2260
rect 9640 2250 9680 2260
rect 0 2240 840 2250
rect 1000 2240 1840 2250
rect 3360 2240 4320 2250
rect 6480 2240 6720 2250
rect 7160 2240 7200 2250
rect 7520 2240 7600 2250
rect 8360 2240 8600 2250
rect 9160 2240 9240 2250
rect 9640 2240 9680 2250
rect 0 2230 840 2240
rect 1000 2230 1840 2240
rect 3360 2230 4320 2240
rect 6480 2230 6720 2240
rect 7160 2230 7200 2240
rect 7520 2230 7600 2240
rect 8360 2230 8600 2240
rect 9160 2230 9240 2240
rect 9640 2230 9680 2240
rect 0 2220 840 2230
rect 1000 2220 1840 2230
rect 3360 2220 4320 2230
rect 6480 2220 6720 2230
rect 7160 2220 7200 2230
rect 7520 2220 7600 2230
rect 8360 2220 8600 2230
rect 9160 2220 9240 2230
rect 9640 2220 9680 2230
rect 0 2210 800 2220
rect 1000 2210 1840 2220
rect 3360 2210 4360 2220
rect 6480 2210 6720 2220
rect 7000 2210 7280 2220
rect 7520 2210 7640 2220
rect 8360 2210 8840 2220
rect 9000 2210 9240 2220
rect 0 2200 800 2210
rect 1000 2200 1840 2210
rect 3360 2200 4360 2210
rect 6480 2200 6720 2210
rect 7000 2200 7280 2210
rect 7520 2200 7640 2210
rect 8360 2200 8840 2210
rect 9000 2200 9240 2210
rect 0 2190 800 2200
rect 1000 2190 1840 2200
rect 3360 2190 4360 2200
rect 6480 2190 6720 2200
rect 7000 2190 7280 2200
rect 7520 2190 7640 2200
rect 8360 2190 8840 2200
rect 9000 2190 9240 2200
rect 0 2180 800 2190
rect 1000 2180 1840 2190
rect 3360 2180 4360 2190
rect 6480 2180 6720 2190
rect 7000 2180 7280 2190
rect 7520 2180 7640 2190
rect 8360 2180 8840 2190
rect 9000 2180 9240 2190
rect 0 2170 800 2180
rect 1000 2170 1840 2180
rect 2680 2170 2720 2180
rect 3360 2170 4360 2180
rect 6520 2170 6720 2180
rect 7080 2170 7280 2180
rect 7320 2170 7360 2180
rect 7520 2170 7680 2180
rect 8400 2170 9240 2180
rect 0 2160 800 2170
rect 1000 2160 1840 2170
rect 2680 2160 2720 2170
rect 3360 2160 4360 2170
rect 6520 2160 6720 2170
rect 7080 2160 7280 2170
rect 7320 2160 7360 2170
rect 7520 2160 7680 2170
rect 8400 2160 9240 2170
rect 0 2150 800 2160
rect 1000 2150 1840 2160
rect 2680 2150 2720 2160
rect 3360 2150 4360 2160
rect 6520 2150 6720 2160
rect 7080 2150 7280 2160
rect 7320 2150 7360 2160
rect 7520 2150 7680 2160
rect 8400 2150 9240 2160
rect 0 2140 800 2150
rect 1000 2140 1840 2150
rect 2680 2140 2720 2150
rect 3360 2140 4360 2150
rect 6520 2140 6720 2150
rect 7080 2140 7280 2150
rect 7320 2140 7360 2150
rect 7520 2140 7680 2150
rect 8400 2140 9240 2150
rect 0 2130 760 2140
rect 960 2130 1840 2140
rect 3360 2130 4360 2140
rect 6520 2130 6720 2140
rect 7320 2130 7400 2140
rect 7480 2130 7720 2140
rect 8400 2130 9200 2140
rect 0 2120 760 2130
rect 960 2120 1840 2130
rect 3360 2120 4360 2130
rect 6520 2120 6720 2130
rect 7320 2120 7400 2130
rect 7480 2120 7720 2130
rect 8400 2120 9200 2130
rect 0 2110 760 2120
rect 960 2110 1840 2120
rect 3360 2110 4360 2120
rect 6520 2110 6720 2120
rect 7320 2110 7400 2120
rect 7480 2110 7720 2120
rect 8400 2110 9200 2120
rect 0 2100 760 2110
rect 960 2100 1840 2110
rect 3360 2100 4360 2110
rect 6520 2100 6720 2110
rect 7320 2100 7400 2110
rect 7480 2100 7720 2110
rect 8400 2100 9200 2110
rect 0 2090 760 2100
rect 960 2090 1840 2100
rect 3360 2090 4320 2100
rect 6560 2090 6760 2100
rect 7320 2090 7840 2100
rect 8480 2090 9200 2100
rect 9600 2090 9640 2100
rect 0 2080 760 2090
rect 960 2080 1840 2090
rect 3360 2080 4320 2090
rect 6560 2080 6760 2090
rect 7320 2080 7840 2090
rect 8480 2080 9200 2090
rect 9600 2080 9640 2090
rect 0 2070 760 2080
rect 960 2070 1840 2080
rect 3360 2070 4320 2080
rect 6560 2070 6760 2080
rect 7320 2070 7840 2080
rect 8480 2070 9200 2080
rect 9600 2070 9640 2080
rect 0 2060 760 2070
rect 960 2060 1840 2070
rect 3360 2060 4320 2070
rect 6560 2060 6760 2070
rect 7320 2060 7840 2070
rect 8480 2060 9200 2070
rect 9600 2060 9640 2070
rect 0 2050 720 2060
rect 960 2050 1840 2060
rect 3360 2050 4360 2060
rect 6560 2050 6760 2060
rect 7360 2050 7720 2060
rect 7800 2050 7840 2060
rect 8560 2050 9080 2060
rect 9280 2050 9320 2060
rect 9400 2050 9440 2060
rect 0 2040 720 2050
rect 960 2040 1840 2050
rect 3360 2040 4360 2050
rect 6560 2040 6760 2050
rect 7360 2040 7720 2050
rect 7800 2040 7840 2050
rect 8560 2040 9080 2050
rect 9280 2040 9320 2050
rect 9400 2040 9440 2050
rect 0 2030 720 2040
rect 960 2030 1840 2040
rect 3360 2030 4360 2040
rect 6560 2030 6760 2040
rect 7360 2030 7720 2040
rect 7800 2030 7840 2040
rect 8560 2030 9080 2040
rect 9280 2030 9320 2040
rect 9400 2030 9440 2040
rect 0 2020 720 2030
rect 960 2020 1840 2030
rect 3360 2020 4360 2030
rect 6560 2020 6760 2030
rect 7360 2020 7720 2030
rect 7800 2020 7840 2030
rect 8560 2020 9080 2030
rect 9280 2020 9320 2030
rect 9400 2020 9440 2030
rect 0 2010 720 2020
rect 960 2010 1840 2020
rect 3360 2010 4320 2020
rect 6560 2010 6760 2020
rect 7360 2010 7720 2020
rect 8680 2010 9040 2020
rect 0 2000 720 2010
rect 960 2000 1840 2010
rect 3360 2000 4320 2010
rect 6560 2000 6760 2010
rect 7360 2000 7720 2010
rect 8680 2000 9040 2010
rect 0 1990 720 2000
rect 960 1990 1840 2000
rect 3360 1990 4320 2000
rect 6560 1990 6760 2000
rect 7360 1990 7720 2000
rect 8680 1990 9040 2000
rect 0 1980 720 1990
rect 960 1980 1840 1990
rect 3360 1980 4320 1990
rect 6560 1980 6760 1990
rect 7360 1980 7720 1990
rect 8680 1980 9040 1990
rect 0 1970 680 1980
rect 960 1970 1840 1980
rect 3360 1970 4360 1980
rect 6560 1970 6760 1980
rect 7360 1970 7720 1980
rect 0 1960 680 1970
rect 960 1960 1840 1970
rect 3360 1960 4360 1970
rect 6560 1960 6760 1970
rect 7360 1960 7720 1970
rect 0 1950 680 1960
rect 960 1950 1840 1960
rect 3360 1950 4360 1960
rect 6560 1950 6760 1960
rect 7360 1950 7720 1960
rect 0 1940 680 1950
rect 960 1940 1840 1950
rect 3360 1940 4360 1950
rect 6560 1940 6760 1950
rect 7360 1940 7720 1950
rect 0 1930 680 1940
rect 920 1930 1840 1940
rect 3360 1930 4360 1940
rect 6560 1930 6760 1940
rect 7360 1930 7720 1940
rect 0 1920 680 1930
rect 920 1920 1840 1930
rect 3360 1920 4360 1930
rect 6560 1920 6760 1930
rect 7360 1920 7720 1930
rect 0 1910 680 1920
rect 920 1910 1840 1920
rect 3360 1910 4360 1920
rect 6560 1910 6760 1920
rect 7360 1910 7720 1920
rect 0 1900 680 1910
rect 920 1900 1840 1910
rect 3360 1900 4360 1910
rect 6560 1900 6760 1910
rect 7360 1900 7720 1910
rect 0 1890 640 1900
rect 920 1890 1840 1900
rect 3360 1890 4280 1900
rect 6600 1890 6760 1900
rect 7360 1890 7720 1900
rect 0 1880 640 1890
rect 920 1880 1840 1890
rect 3360 1880 4280 1890
rect 6600 1880 6760 1890
rect 7360 1880 7720 1890
rect 0 1870 640 1880
rect 920 1870 1840 1880
rect 3360 1870 4280 1880
rect 6600 1870 6760 1880
rect 7360 1870 7720 1880
rect 0 1860 640 1870
rect 920 1860 1840 1870
rect 3360 1860 4280 1870
rect 6600 1860 6760 1870
rect 7360 1860 7720 1870
rect 0 1850 640 1860
rect 920 1850 1840 1860
rect 2760 1850 2800 1860
rect 3360 1850 4280 1860
rect 6600 1850 6800 1860
rect 7360 1850 7720 1860
rect 0 1840 640 1850
rect 920 1840 1840 1850
rect 2760 1840 2800 1850
rect 3360 1840 4280 1850
rect 6600 1840 6800 1850
rect 7360 1840 7720 1850
rect 0 1830 640 1840
rect 920 1830 1840 1840
rect 2760 1830 2800 1840
rect 3360 1830 4280 1840
rect 6600 1830 6800 1840
rect 7360 1830 7720 1840
rect 0 1820 640 1830
rect 920 1820 1840 1830
rect 2760 1820 2800 1830
rect 3360 1820 4280 1830
rect 6600 1820 6800 1830
rect 7360 1820 7720 1830
rect 0 1810 600 1820
rect 920 1810 1840 1820
rect 3320 1810 4080 1820
rect 4200 1810 4280 1820
rect 6600 1810 6800 1820
rect 7360 1810 7760 1820
rect 0 1800 600 1810
rect 920 1800 1840 1810
rect 3320 1800 4080 1810
rect 4200 1800 4280 1810
rect 6600 1800 6800 1810
rect 7360 1800 7760 1810
rect 0 1790 600 1800
rect 920 1790 1840 1800
rect 3320 1790 4080 1800
rect 4200 1790 4280 1800
rect 6600 1790 6800 1800
rect 7360 1790 7760 1800
rect 0 1780 600 1790
rect 920 1780 1840 1790
rect 3320 1780 4080 1790
rect 4200 1780 4280 1790
rect 6600 1780 6800 1790
rect 7360 1780 7760 1790
rect 0 1770 600 1780
rect 920 1770 1840 1780
rect 3320 1770 4040 1780
rect 4240 1770 4280 1780
rect 6640 1770 6800 1780
rect 7360 1770 7760 1780
rect 0 1760 600 1770
rect 920 1760 1840 1770
rect 3320 1760 4040 1770
rect 4240 1760 4280 1770
rect 6640 1760 6800 1770
rect 7360 1760 7760 1770
rect 0 1750 600 1760
rect 920 1750 1840 1760
rect 3320 1750 4040 1760
rect 4240 1750 4280 1760
rect 6640 1750 6800 1760
rect 7360 1750 7760 1760
rect 0 1740 600 1750
rect 920 1740 1840 1750
rect 3320 1740 4040 1750
rect 4240 1740 4280 1750
rect 6640 1740 6800 1750
rect 7360 1740 7760 1750
rect 0 1730 560 1740
rect 880 1730 1880 1740
rect 3320 1730 4040 1740
rect 4240 1730 4280 1740
rect 4320 1730 4360 1740
rect 6680 1730 6800 1740
rect 7360 1730 7760 1740
rect 0 1720 560 1730
rect 880 1720 1880 1730
rect 3320 1720 4040 1730
rect 4240 1720 4280 1730
rect 4320 1720 4360 1730
rect 6680 1720 6800 1730
rect 7360 1720 7760 1730
rect 0 1710 560 1720
rect 880 1710 1880 1720
rect 3320 1710 4040 1720
rect 4240 1710 4280 1720
rect 4320 1710 4360 1720
rect 6680 1710 6800 1720
rect 7360 1710 7760 1720
rect 0 1700 560 1710
rect 880 1700 1880 1710
rect 3320 1700 4040 1710
rect 4240 1700 4280 1710
rect 4320 1700 4360 1710
rect 6680 1700 6800 1710
rect 7360 1700 7760 1710
rect 0 1690 560 1700
rect 880 1690 1880 1700
rect 3280 1690 4040 1700
rect 4320 1690 4360 1700
rect 6200 1690 6240 1700
rect 6680 1690 6800 1700
rect 7360 1690 7760 1700
rect 0 1680 560 1690
rect 880 1680 1880 1690
rect 3280 1680 4040 1690
rect 4320 1680 4360 1690
rect 6200 1680 6240 1690
rect 6680 1680 6800 1690
rect 7360 1680 7760 1690
rect 0 1670 560 1680
rect 880 1670 1880 1680
rect 3280 1670 4040 1680
rect 4320 1670 4360 1680
rect 6200 1670 6240 1680
rect 6680 1670 6800 1680
rect 7360 1670 7760 1680
rect 0 1660 560 1670
rect 880 1660 1880 1670
rect 3280 1660 4040 1670
rect 4320 1660 4360 1670
rect 6200 1660 6240 1670
rect 6680 1660 6800 1670
rect 7360 1660 7760 1670
rect 0 1650 560 1660
rect 880 1650 1880 1660
rect 3280 1650 4080 1660
rect 4320 1650 4360 1660
rect 6200 1650 6280 1660
rect 6680 1650 6800 1660
rect 7360 1650 7760 1660
rect 0 1640 560 1650
rect 880 1640 1880 1650
rect 3280 1640 4080 1650
rect 4320 1640 4360 1650
rect 6200 1640 6280 1650
rect 6680 1640 6800 1650
rect 7360 1640 7760 1650
rect 0 1630 560 1640
rect 880 1630 1880 1640
rect 3280 1630 4080 1640
rect 4320 1630 4360 1640
rect 6200 1630 6280 1640
rect 6680 1630 6800 1640
rect 7360 1630 7760 1640
rect 0 1620 560 1630
rect 880 1620 1880 1630
rect 3280 1620 4080 1630
rect 4320 1620 4360 1630
rect 6200 1620 6280 1630
rect 6680 1620 6800 1630
rect 7360 1620 7760 1630
rect 0 1610 520 1620
rect 880 1610 1920 1620
rect 3240 1610 4080 1620
rect 4400 1610 4440 1620
rect 6200 1610 6280 1620
rect 6720 1610 6800 1620
rect 7400 1610 7760 1620
rect 0 1600 520 1610
rect 880 1600 1920 1610
rect 3240 1600 4080 1610
rect 4400 1600 4440 1610
rect 6200 1600 6280 1610
rect 6720 1600 6800 1610
rect 7400 1600 7760 1610
rect 0 1590 520 1600
rect 880 1590 1920 1600
rect 3240 1590 4080 1600
rect 4400 1590 4440 1600
rect 6200 1590 6280 1600
rect 6720 1590 6800 1600
rect 7400 1590 7760 1600
rect 0 1580 520 1590
rect 880 1580 1920 1590
rect 3240 1580 4080 1590
rect 4400 1580 4440 1590
rect 6200 1580 6280 1590
rect 6720 1580 6800 1590
rect 7400 1580 7760 1590
rect 0 1570 520 1580
rect 840 1570 1920 1580
rect 3200 1570 4080 1580
rect 4360 1570 4480 1580
rect 6240 1570 6280 1580
rect 6720 1570 6800 1580
rect 7400 1570 7760 1580
rect 0 1560 520 1570
rect 840 1560 1920 1570
rect 3200 1560 4080 1570
rect 4360 1560 4480 1570
rect 6240 1560 6280 1570
rect 6720 1560 6800 1570
rect 7400 1560 7760 1570
rect 0 1550 520 1560
rect 840 1550 1920 1560
rect 3200 1550 4080 1560
rect 4360 1550 4480 1560
rect 6240 1550 6280 1560
rect 6720 1550 6800 1560
rect 7400 1550 7760 1560
rect 0 1540 520 1550
rect 840 1540 1920 1550
rect 3200 1540 4080 1550
rect 4360 1540 4480 1550
rect 6240 1540 6280 1550
rect 6720 1540 6800 1550
rect 7400 1540 7760 1550
rect 0 1530 520 1540
rect 840 1530 1960 1540
rect 3200 1530 4120 1540
rect 6240 1530 6280 1540
rect 7400 1530 7800 1540
rect 0 1520 520 1530
rect 840 1520 1960 1530
rect 3200 1520 4120 1530
rect 6240 1520 6280 1530
rect 7400 1520 7800 1530
rect 0 1510 520 1520
rect 840 1510 1960 1520
rect 3200 1510 4120 1520
rect 6240 1510 6280 1520
rect 7400 1510 7800 1520
rect 0 1500 520 1510
rect 840 1500 1960 1510
rect 3200 1500 4120 1510
rect 6240 1500 6280 1510
rect 7400 1500 7800 1510
rect 0 1490 480 1500
rect 840 1490 920 1500
rect 1000 1490 2000 1500
rect 3160 1490 4120 1500
rect 4440 1490 4480 1500
rect 6200 1490 6280 1500
rect 7400 1490 7800 1500
rect 0 1480 480 1490
rect 840 1480 920 1490
rect 1000 1480 2000 1490
rect 3160 1480 4120 1490
rect 4440 1480 4480 1490
rect 6200 1480 6280 1490
rect 7400 1480 7800 1490
rect 0 1470 480 1480
rect 840 1470 920 1480
rect 1000 1470 2000 1480
rect 3160 1470 4120 1480
rect 4440 1470 4480 1480
rect 6200 1470 6280 1480
rect 7400 1470 7800 1480
rect 0 1460 480 1470
rect 840 1460 920 1470
rect 1000 1460 2000 1470
rect 3160 1460 4120 1470
rect 4440 1460 4480 1470
rect 6200 1460 6280 1470
rect 7400 1460 7800 1470
rect 0 1450 480 1460
rect 1040 1450 2000 1460
rect 3120 1450 4120 1460
rect 4400 1450 4440 1460
rect 6200 1450 6320 1460
rect 7400 1450 7800 1460
rect 0 1440 480 1450
rect 1040 1440 2000 1450
rect 3120 1440 4120 1450
rect 4400 1440 4440 1450
rect 6200 1440 6320 1450
rect 7400 1440 7800 1450
rect 0 1430 480 1440
rect 1040 1430 2000 1440
rect 3120 1430 4120 1440
rect 4400 1430 4440 1440
rect 6200 1430 6320 1440
rect 7400 1430 7800 1440
rect 0 1420 480 1430
rect 1040 1420 2000 1430
rect 3120 1420 4120 1430
rect 4400 1420 4440 1430
rect 6200 1420 6320 1430
rect 7400 1420 7800 1430
rect 0 1410 480 1420
rect 1040 1410 2040 1420
rect 3080 1410 4160 1420
rect 4400 1410 4440 1420
rect 6200 1410 6320 1420
rect 7400 1410 7800 1420
rect 0 1400 480 1410
rect 1040 1400 2040 1410
rect 3080 1400 4160 1410
rect 4400 1400 4440 1410
rect 6200 1400 6320 1410
rect 7400 1400 7800 1410
rect 0 1390 480 1400
rect 1040 1390 2040 1400
rect 3080 1390 4160 1400
rect 4400 1390 4440 1400
rect 6200 1390 6320 1400
rect 7400 1390 7800 1400
rect 0 1380 480 1390
rect 1040 1380 2040 1390
rect 3080 1380 4160 1390
rect 4400 1380 4440 1390
rect 6200 1380 6320 1390
rect 7400 1380 7800 1390
rect 0 1370 440 1380
rect 1040 1370 2080 1380
rect 3000 1370 3520 1380
rect 3640 1370 4160 1380
rect 6200 1370 6320 1380
rect 7400 1370 7840 1380
rect 0 1360 440 1370
rect 1040 1360 2080 1370
rect 3000 1360 3520 1370
rect 3640 1360 4160 1370
rect 6200 1360 6320 1370
rect 7400 1360 7840 1370
rect 0 1350 440 1360
rect 1040 1350 2080 1360
rect 3000 1350 3520 1360
rect 3640 1350 4160 1360
rect 6200 1350 6320 1360
rect 7400 1350 7840 1360
rect 0 1340 440 1350
rect 1040 1340 2080 1350
rect 3000 1340 3520 1350
rect 3640 1340 4160 1350
rect 6200 1340 6320 1350
rect 7400 1340 7840 1350
rect 0 1330 440 1340
rect 1040 1330 2080 1340
rect 2960 1330 3480 1340
rect 3680 1330 4160 1340
rect 6200 1330 6320 1340
rect 7400 1330 7840 1340
rect 0 1320 440 1330
rect 1040 1320 2080 1330
rect 2960 1320 3480 1330
rect 3680 1320 4160 1330
rect 6200 1320 6320 1330
rect 7400 1320 7840 1330
rect 0 1310 440 1320
rect 1040 1310 2080 1320
rect 2960 1310 3480 1320
rect 3680 1310 4160 1320
rect 6200 1310 6320 1320
rect 7400 1310 7840 1320
rect 0 1300 440 1310
rect 1040 1300 2080 1310
rect 2960 1300 3480 1310
rect 3680 1300 4160 1310
rect 6200 1300 6320 1310
rect 7400 1300 7840 1310
rect 0 1290 440 1300
rect 1000 1290 2040 1300
rect 2880 1290 3480 1300
rect 3760 1290 4200 1300
rect 6200 1290 6320 1300
rect 7440 1290 7840 1300
rect 0 1280 440 1290
rect 1000 1280 2040 1290
rect 2880 1280 3480 1290
rect 3760 1280 4200 1290
rect 6200 1280 6320 1290
rect 7440 1280 7840 1290
rect 0 1270 440 1280
rect 1000 1270 2040 1280
rect 2880 1270 3480 1280
rect 3760 1270 4200 1280
rect 6200 1270 6320 1280
rect 7440 1270 7840 1280
rect 0 1260 440 1270
rect 1000 1260 2040 1270
rect 2880 1260 3480 1270
rect 3760 1260 4200 1270
rect 6200 1260 6320 1270
rect 7440 1260 7840 1270
rect 0 1250 400 1260
rect 1000 1250 2040 1260
rect 2840 1250 3480 1260
rect 3800 1250 4200 1260
rect 6240 1250 6320 1260
rect 7440 1250 7840 1260
rect 0 1240 400 1250
rect 1000 1240 2040 1250
rect 2840 1240 3480 1250
rect 3800 1240 4200 1250
rect 6240 1240 6320 1250
rect 7440 1240 7840 1250
rect 0 1230 400 1240
rect 1000 1230 2040 1240
rect 2840 1230 3480 1240
rect 3800 1230 4200 1240
rect 6240 1230 6320 1240
rect 7440 1230 7840 1240
rect 0 1220 400 1230
rect 1000 1220 2040 1230
rect 2840 1220 3480 1230
rect 3800 1220 4200 1230
rect 6240 1220 6320 1230
rect 7440 1220 7840 1230
rect 0 1210 400 1220
rect 1000 1210 2000 1220
rect 2760 1210 3520 1220
rect 3840 1210 4200 1220
rect 6240 1210 6360 1220
rect 7440 1210 7840 1220
rect 0 1200 400 1210
rect 1000 1200 2000 1210
rect 2760 1200 3520 1210
rect 3840 1200 4200 1210
rect 6240 1200 6360 1210
rect 7440 1200 7840 1210
rect 0 1190 400 1200
rect 1000 1190 2000 1200
rect 2760 1190 3520 1200
rect 3840 1190 4200 1200
rect 6240 1190 6360 1200
rect 7440 1190 7840 1200
rect 0 1180 400 1190
rect 1000 1180 2000 1190
rect 2760 1180 3520 1190
rect 3840 1180 4200 1190
rect 6240 1180 6360 1190
rect 7440 1180 7840 1190
rect 0 1170 400 1180
rect 1000 1170 2000 1180
rect 2880 1170 3560 1180
rect 3920 1170 4200 1180
rect 6280 1170 6360 1180
rect 7440 1170 7880 1180
rect 0 1160 400 1170
rect 1000 1160 2000 1170
rect 2880 1160 3560 1170
rect 3920 1160 4200 1170
rect 6280 1160 6360 1170
rect 7440 1160 7880 1170
rect 0 1150 400 1160
rect 1000 1150 2000 1160
rect 2880 1150 3560 1160
rect 3920 1150 4200 1160
rect 6280 1150 6360 1160
rect 7440 1150 7880 1160
rect 0 1140 400 1150
rect 1000 1140 2000 1150
rect 2880 1140 3560 1150
rect 3920 1140 4200 1150
rect 6280 1140 6360 1150
rect 7440 1140 7880 1150
rect 0 1130 360 1140
rect 640 1130 760 1140
rect 1000 1130 1560 1140
rect 1600 1130 2000 1140
rect 2880 1130 3600 1140
rect 3960 1130 4200 1140
rect 6280 1130 6400 1140
rect 7440 1130 7880 1140
rect 0 1120 360 1130
rect 640 1120 760 1130
rect 1000 1120 1560 1130
rect 1600 1120 2000 1130
rect 2880 1120 3600 1130
rect 3960 1120 4200 1130
rect 6280 1120 6400 1130
rect 7440 1120 7880 1130
rect 0 1110 360 1120
rect 640 1110 760 1120
rect 1000 1110 1560 1120
rect 1600 1110 2000 1120
rect 2880 1110 3600 1120
rect 3960 1110 4200 1120
rect 6280 1110 6400 1120
rect 7440 1110 7880 1120
rect 0 1100 360 1110
rect 640 1100 760 1110
rect 1000 1100 1560 1110
rect 1600 1100 2000 1110
rect 2880 1100 3600 1110
rect 3960 1100 4200 1110
rect 6280 1100 6400 1110
rect 7440 1100 7880 1110
rect 0 1090 360 1100
rect 640 1090 720 1100
rect 1000 1090 1480 1100
rect 1640 1090 1960 1100
rect 2920 1090 3640 1100
rect 4040 1090 4080 1100
rect 4120 1090 4200 1100
rect 6280 1090 6440 1100
rect 7440 1090 7880 1100
rect 0 1080 360 1090
rect 640 1080 720 1090
rect 1000 1080 1480 1090
rect 1640 1080 1960 1090
rect 2920 1080 3640 1090
rect 4040 1080 4080 1090
rect 4120 1080 4200 1090
rect 6280 1080 6440 1090
rect 7440 1080 7880 1090
rect 0 1070 360 1080
rect 640 1070 720 1080
rect 1000 1070 1480 1080
rect 1640 1070 1960 1080
rect 2920 1070 3640 1080
rect 4040 1070 4080 1080
rect 4120 1070 4200 1080
rect 6280 1070 6440 1080
rect 7440 1070 7880 1080
rect 0 1060 360 1070
rect 640 1060 720 1070
rect 1000 1060 1480 1070
rect 1640 1060 1960 1070
rect 2920 1060 3640 1070
rect 4040 1060 4080 1070
rect 4120 1060 4200 1070
rect 6280 1060 6440 1070
rect 7440 1060 7880 1070
rect 0 1050 320 1060
rect 640 1050 720 1060
rect 960 1050 1440 1060
rect 1680 1050 1960 1060
rect 2920 1050 3680 1060
rect 4120 1050 4200 1060
rect 6280 1050 6400 1060
rect 7440 1050 7880 1060
rect 0 1040 320 1050
rect 640 1040 720 1050
rect 960 1040 1440 1050
rect 1680 1040 1960 1050
rect 2920 1040 3680 1050
rect 4120 1040 4200 1050
rect 6280 1040 6400 1050
rect 7440 1040 7880 1050
rect 0 1030 320 1040
rect 640 1030 720 1040
rect 960 1030 1440 1040
rect 1680 1030 1960 1040
rect 2920 1030 3680 1040
rect 4120 1030 4200 1040
rect 6280 1030 6400 1040
rect 7440 1030 7880 1040
rect 0 1020 320 1030
rect 640 1020 720 1030
rect 960 1020 1440 1030
rect 1680 1020 1960 1030
rect 2920 1020 3680 1030
rect 4120 1020 4200 1030
rect 6280 1020 6400 1030
rect 7440 1020 7880 1030
rect 0 1010 320 1020
rect 680 1010 720 1020
rect 960 1010 1400 1020
rect 1640 1010 1960 1020
rect 2920 1010 3680 1020
rect 6320 1010 6360 1020
rect 7440 1010 7880 1020
rect 0 1000 320 1010
rect 680 1000 720 1010
rect 960 1000 1400 1010
rect 1640 1000 1960 1010
rect 2920 1000 3680 1010
rect 6320 1000 6360 1010
rect 7440 1000 7880 1010
rect 0 990 320 1000
rect 680 990 720 1000
rect 960 990 1400 1000
rect 1640 990 1960 1000
rect 2920 990 3680 1000
rect 6320 990 6360 1000
rect 7440 990 7880 1000
rect 0 980 320 990
rect 680 980 720 990
rect 960 980 1400 990
rect 1640 980 1960 990
rect 2920 980 3680 990
rect 6320 980 6360 990
rect 7440 980 7880 990
rect 0 970 280 980
rect 960 970 1360 980
rect 1600 970 1960 980
rect 2880 970 3760 980
rect 6320 970 6360 980
rect 7440 970 7920 980
rect 0 960 280 970
rect 960 960 1360 970
rect 1600 960 1960 970
rect 2880 960 3760 970
rect 6320 960 6360 970
rect 7440 960 7920 970
rect 0 950 280 960
rect 960 950 1360 960
rect 1600 950 1960 960
rect 2880 950 3760 960
rect 6320 950 6360 960
rect 7440 950 7920 960
rect 0 940 280 950
rect 960 940 1360 950
rect 1600 940 1960 950
rect 2880 940 3760 950
rect 6320 940 6360 950
rect 7440 940 7920 950
rect 0 930 280 940
rect 960 930 1320 940
rect 1560 930 1960 940
rect 2840 930 3800 940
rect 4840 930 4880 940
rect 5160 930 5200 940
rect 6320 930 6360 940
rect 7440 930 7920 940
rect 0 920 280 930
rect 960 920 1320 930
rect 1560 920 1960 930
rect 2840 920 3800 930
rect 4840 920 4880 930
rect 5160 920 5200 930
rect 6320 920 6360 930
rect 7440 920 7920 930
rect 0 910 280 920
rect 960 910 1320 920
rect 1560 910 1960 920
rect 2840 910 3800 920
rect 4840 910 4880 920
rect 5160 910 5200 920
rect 6320 910 6360 920
rect 7440 910 7920 920
rect 0 900 280 910
rect 960 900 1320 910
rect 1560 900 1960 910
rect 2840 900 3800 910
rect 4840 900 4880 910
rect 5160 900 5200 910
rect 6320 900 6360 910
rect 7440 900 7920 910
rect 0 890 240 900
rect 960 890 1240 900
rect 1520 890 2000 900
rect 2760 890 3800 900
rect 4880 890 5080 900
rect 5200 890 5280 900
rect 6320 890 6360 900
rect 7440 890 7920 900
rect 0 880 240 890
rect 960 880 1240 890
rect 1520 880 2000 890
rect 2760 880 3800 890
rect 4880 880 5080 890
rect 5200 880 5280 890
rect 6320 880 6360 890
rect 7440 880 7920 890
rect 0 870 240 880
rect 960 870 1240 880
rect 1520 870 2000 880
rect 2760 870 3800 880
rect 4880 870 5080 880
rect 5200 870 5280 880
rect 6320 870 6360 880
rect 7440 870 7920 880
rect 0 860 240 870
rect 960 860 1240 870
rect 1520 860 2000 870
rect 2760 860 3800 870
rect 4880 860 5080 870
rect 5200 860 5280 870
rect 6320 860 6360 870
rect 7440 860 7920 870
rect 0 850 200 860
rect 920 850 1200 860
rect 1480 850 2000 860
rect 2680 850 3840 860
rect 4920 850 5200 860
rect 5320 850 5360 860
rect 6320 850 6400 860
rect 7440 850 7920 860
rect 0 840 200 850
rect 920 840 1200 850
rect 1480 840 2000 850
rect 2680 840 3840 850
rect 4920 840 5200 850
rect 5320 840 5360 850
rect 6320 840 6400 850
rect 7440 840 7920 850
rect 0 830 200 840
rect 920 830 1200 840
rect 1480 830 2000 840
rect 2680 830 3840 840
rect 4920 830 5200 840
rect 5320 830 5360 840
rect 6320 830 6400 840
rect 7440 830 7920 840
rect 0 820 200 830
rect 920 820 1200 830
rect 1480 820 2000 830
rect 2680 820 3840 830
rect 4920 820 5200 830
rect 5320 820 5360 830
rect 6320 820 6400 830
rect 7440 820 7920 830
rect 0 810 160 820
rect 920 810 1160 820
rect 1480 810 2000 820
rect 2600 810 3880 820
rect 4920 810 5160 820
rect 6320 810 6400 820
rect 7440 810 7920 820
rect 0 800 160 810
rect 920 800 1160 810
rect 1480 800 2000 810
rect 2600 800 3880 810
rect 4920 800 5160 810
rect 6320 800 6400 810
rect 7440 800 7920 810
rect 0 790 160 800
rect 920 790 1160 800
rect 1480 790 2000 800
rect 2600 790 3880 800
rect 4920 790 5160 800
rect 6320 790 6400 800
rect 7440 790 7920 800
rect 0 780 160 790
rect 920 780 1160 790
rect 1480 780 2000 790
rect 2600 780 3880 790
rect 4920 780 5160 790
rect 6320 780 6400 790
rect 7440 780 7920 790
rect 0 770 120 780
rect 920 770 1080 780
rect 1440 770 2040 780
rect 2560 770 3520 780
rect 3920 770 3960 780
rect 4920 770 5320 780
rect 5360 770 5400 780
rect 6320 770 6400 780
rect 7440 770 7960 780
rect 0 760 120 770
rect 920 760 1080 770
rect 1440 760 2040 770
rect 2560 760 3520 770
rect 3920 760 3960 770
rect 4920 760 5320 770
rect 5360 760 5400 770
rect 6320 760 6400 770
rect 7440 760 7960 770
rect 0 750 120 760
rect 920 750 1080 760
rect 1440 750 2040 760
rect 2560 750 3520 760
rect 3920 750 3960 760
rect 4920 750 5320 760
rect 5360 750 5400 760
rect 6320 750 6400 760
rect 7440 750 7960 760
rect 0 740 120 750
rect 920 740 1080 750
rect 1440 740 2040 750
rect 2560 740 3520 750
rect 3920 740 3960 750
rect 4920 740 5320 750
rect 5360 740 5400 750
rect 6320 740 6400 750
rect 7440 740 7960 750
rect 0 730 80 740
rect 920 730 1040 740
rect 1400 730 2040 740
rect 2480 730 3360 740
rect 3960 730 4000 740
rect 4920 730 5120 740
rect 5200 730 5360 740
rect 5400 730 5440 740
rect 6320 730 6440 740
rect 7440 730 7960 740
rect 0 720 80 730
rect 920 720 1040 730
rect 1400 720 2040 730
rect 2480 720 3360 730
rect 3960 720 4000 730
rect 4920 720 5120 730
rect 5200 720 5360 730
rect 5400 720 5440 730
rect 6320 720 6440 730
rect 7440 720 7960 730
rect 0 710 80 720
rect 920 710 1040 720
rect 1400 710 2040 720
rect 2480 710 3360 720
rect 3960 710 4000 720
rect 4920 710 5120 720
rect 5200 710 5360 720
rect 5400 710 5440 720
rect 6320 710 6440 720
rect 7440 710 7960 720
rect 0 700 80 710
rect 920 700 1040 710
rect 1400 700 2040 710
rect 2480 700 3360 710
rect 3960 700 4000 710
rect 4920 700 5120 710
rect 5200 700 5360 710
rect 5400 700 5440 710
rect 6320 700 6440 710
rect 7440 700 7960 710
rect 0 690 40 700
rect 1360 690 2080 700
rect 2400 690 3280 700
rect 4960 690 5120 700
rect 5200 690 5400 700
rect 5440 690 5480 700
rect 6360 690 6440 700
rect 7440 690 7960 700
rect 0 680 40 690
rect 1360 680 2080 690
rect 2400 680 3280 690
rect 4960 680 5120 690
rect 5200 680 5400 690
rect 5440 680 5480 690
rect 6360 680 6440 690
rect 7440 680 7960 690
rect 0 670 40 680
rect 1360 670 2080 680
rect 2400 670 3280 680
rect 4960 670 5120 680
rect 5200 670 5400 680
rect 5440 670 5480 680
rect 6360 670 6440 680
rect 7440 670 7960 680
rect 0 660 40 670
rect 1360 660 2080 670
rect 2400 660 3280 670
rect 4960 660 5120 670
rect 5200 660 5400 670
rect 5440 660 5480 670
rect 6360 660 6440 670
rect 7440 660 7960 670
rect 1360 650 2080 660
rect 2320 650 3200 660
rect 4960 650 5160 660
rect 5200 650 5280 660
rect 5320 650 5400 660
rect 5440 650 5480 660
rect 6360 650 6480 660
rect 7440 650 8000 660
rect 1360 640 2080 650
rect 2320 640 3200 650
rect 4960 640 5160 650
rect 5200 640 5280 650
rect 5320 640 5400 650
rect 5440 640 5480 650
rect 6360 640 6480 650
rect 7440 640 8000 650
rect 1360 630 2080 640
rect 2320 630 3200 640
rect 4960 630 5160 640
rect 5200 630 5280 640
rect 5320 630 5400 640
rect 5440 630 5480 640
rect 6360 630 6480 640
rect 7440 630 8000 640
rect 1360 620 2080 630
rect 2320 620 3200 630
rect 4960 620 5160 630
rect 5200 620 5280 630
rect 5320 620 5400 630
rect 5440 620 5480 630
rect 6360 620 6480 630
rect 7440 620 8000 630
rect 1440 610 2120 620
rect 2280 610 3120 620
rect 4960 610 5560 620
rect 6360 610 6520 620
rect 7440 610 8000 620
rect 1440 600 2120 610
rect 2280 600 3120 610
rect 4960 600 5560 610
rect 6360 600 6520 610
rect 7440 600 8000 610
rect 1440 590 2120 600
rect 2280 590 3120 600
rect 4960 590 5560 600
rect 6360 590 6520 600
rect 7440 590 8000 600
rect 1440 580 2120 590
rect 2280 580 3120 590
rect 4960 580 5560 590
rect 6360 580 6520 590
rect 7440 580 8000 590
rect 1480 570 2120 580
rect 2200 570 3000 580
rect 4960 570 5560 580
rect 6360 570 6520 580
rect 7440 570 8040 580
rect 1480 560 2120 570
rect 2200 560 3000 570
rect 4960 560 5560 570
rect 6360 560 6520 570
rect 7440 560 8040 570
rect 1480 550 2120 560
rect 2200 550 3000 560
rect 4960 550 5560 560
rect 6360 550 6520 560
rect 7440 550 8040 560
rect 1480 540 2120 550
rect 2200 540 3000 550
rect 4960 540 5560 550
rect 6360 540 6520 550
rect 7440 540 8040 550
rect 1520 530 2880 540
rect 4960 530 5360 540
rect 5480 530 5600 540
rect 6360 530 6560 540
rect 7440 530 8080 540
rect 1520 520 2880 530
rect 4960 520 5360 530
rect 5480 520 5600 530
rect 6360 520 6560 530
rect 7440 520 8080 530
rect 1520 510 2880 520
rect 4960 510 5360 520
rect 5480 510 5600 520
rect 6360 510 6560 520
rect 7440 510 8080 520
rect 1520 500 2880 510
rect 4960 500 5360 510
rect 5480 500 5600 510
rect 6360 500 6560 510
rect 7440 500 8080 510
rect 1560 490 2120 500
rect 2160 490 2760 500
rect 4480 490 4520 500
rect 4960 490 5360 500
rect 5480 490 5680 500
rect 6320 490 6560 500
rect 7440 490 8120 500
rect 1560 480 2120 490
rect 2160 480 2760 490
rect 4480 480 4520 490
rect 4960 480 5360 490
rect 5480 480 5680 490
rect 6320 480 6560 490
rect 7440 480 8120 490
rect 1560 470 2120 480
rect 2160 470 2760 480
rect 4480 470 4520 480
rect 4960 470 5360 480
rect 5480 470 5680 480
rect 6320 470 6560 480
rect 7440 470 8120 480
rect 1560 460 2120 470
rect 2160 460 2760 470
rect 4480 460 4520 470
rect 4960 460 5360 470
rect 5480 460 5680 470
rect 6320 460 6560 470
rect 7440 460 8120 470
rect 680 450 800 460
rect 1720 450 1800 460
rect 2320 450 2560 460
rect 4320 450 4440 460
rect 5000 450 5680 460
rect 6360 450 6600 460
rect 7440 450 8200 460
rect 680 440 800 450
rect 1720 440 1800 450
rect 2320 440 2560 450
rect 4320 440 4440 450
rect 5000 440 5680 450
rect 6360 440 6600 450
rect 7440 440 8200 450
rect 680 430 800 440
rect 1720 430 1800 440
rect 2320 430 2560 440
rect 4320 430 4440 440
rect 5000 430 5680 440
rect 6360 430 6600 440
rect 7440 430 8200 440
rect 680 420 800 430
rect 1720 420 1800 430
rect 2320 420 2560 430
rect 4320 420 4440 430
rect 5000 420 5680 430
rect 6360 420 6600 430
rect 7440 420 8200 430
rect 680 410 760 420
rect 5000 410 5200 420
rect 5280 410 5320 420
rect 5360 410 5720 420
rect 6360 410 6600 420
rect 7440 410 8280 420
rect 680 400 760 410
rect 5000 400 5200 410
rect 5280 400 5320 410
rect 5360 400 5720 410
rect 6360 400 6600 410
rect 7440 400 8280 410
rect 680 390 760 400
rect 5000 390 5200 400
rect 5280 390 5320 400
rect 5360 390 5720 400
rect 6360 390 6600 400
rect 7440 390 8280 400
rect 680 380 760 390
rect 5000 380 5200 390
rect 5280 380 5320 390
rect 5360 380 5720 390
rect 6360 380 6600 390
rect 7440 380 8280 390
rect 680 370 800 380
rect 840 370 920 380
rect 5000 370 5200 380
rect 5280 370 5320 380
rect 5400 370 5760 380
rect 6360 370 6640 380
rect 7440 370 8280 380
rect 680 360 800 370
rect 840 360 920 370
rect 5000 360 5200 370
rect 5280 360 5320 370
rect 5400 360 5760 370
rect 6360 360 6640 370
rect 7440 360 8280 370
rect 680 350 800 360
rect 840 350 920 360
rect 5000 350 5200 360
rect 5280 350 5320 360
rect 5400 350 5760 360
rect 6360 350 6640 360
rect 7440 350 8280 360
rect 680 340 800 350
rect 840 340 920 350
rect 5000 340 5200 350
rect 5280 340 5320 350
rect 5400 340 5760 350
rect 6360 340 6640 350
rect 7440 340 8280 350
rect 840 330 880 340
rect 5000 330 5720 340
rect 6360 330 6680 340
rect 7440 330 8320 340
rect 840 320 880 330
rect 5000 320 5720 330
rect 6360 320 6680 330
rect 7440 320 8320 330
rect 840 310 880 320
rect 5000 310 5720 320
rect 6360 310 6680 320
rect 7440 310 8320 320
rect 840 300 880 310
rect 5000 300 5720 310
rect 6360 300 6680 310
rect 7440 300 8320 310
rect 5000 290 5720 300
rect 5840 290 5880 300
rect 6360 290 6720 300
rect 7440 290 8360 300
rect 5000 280 5720 290
rect 5840 280 5880 290
rect 6360 280 6720 290
rect 7440 280 8360 290
rect 5000 270 5720 280
rect 5840 270 5880 280
rect 6360 270 6720 280
rect 7440 270 8360 280
rect 5000 260 5720 270
rect 5840 260 5880 270
rect 6360 260 6720 270
rect 7440 260 8360 270
rect 5000 250 5720 260
rect 5800 250 5960 260
rect 6360 250 6720 260
rect 7400 250 8400 260
rect 5000 240 5720 250
rect 5800 240 5960 250
rect 6360 240 6720 250
rect 7400 240 8400 250
rect 5000 230 5720 240
rect 5800 230 5960 240
rect 6360 230 6720 240
rect 7400 230 8400 240
rect 5000 220 5720 230
rect 5800 220 5960 230
rect 6360 220 6720 230
rect 7400 220 8400 230
rect 5000 210 6000 220
rect 6360 210 6760 220
rect 7400 210 8440 220
rect 5000 200 6000 210
rect 6360 200 6760 210
rect 7400 200 8440 210
rect 5000 190 6000 200
rect 6360 190 6760 200
rect 7400 190 8440 200
rect 5000 180 6000 190
rect 6360 180 6760 190
rect 7400 180 8440 190
rect 5040 170 5360 180
rect 5720 170 5960 180
rect 6400 170 6800 180
rect 7400 170 8480 180
rect 8920 170 9000 180
rect 5040 160 5360 170
rect 5720 160 5960 170
rect 6400 160 6800 170
rect 7400 160 8480 170
rect 8920 160 9000 170
rect 5040 150 5360 160
rect 5720 150 5960 160
rect 6400 150 6800 160
rect 7400 150 8480 160
rect 8920 150 9000 160
rect 5040 140 5360 150
rect 5720 140 5960 150
rect 6400 140 6800 150
rect 7400 140 8480 150
rect 8920 140 9000 150
rect 400 130 480 140
rect 5040 130 5320 140
rect 6400 130 6800 140
rect 7400 130 8520 140
rect 8960 130 9040 140
rect 400 120 480 130
rect 5040 120 5320 130
rect 6400 120 6800 130
rect 7400 120 8520 130
rect 8960 120 9040 130
rect 400 110 480 120
rect 5040 110 5320 120
rect 6400 110 6800 120
rect 7400 110 8520 120
rect 8960 110 9040 120
rect 400 100 480 110
rect 5040 100 5320 110
rect 6400 100 6800 110
rect 7400 100 8520 110
rect 8960 100 9040 110
rect 360 90 520 100
rect 5040 90 5360 100
rect 6440 90 6840 100
rect 7400 90 8560 100
rect 9280 90 9320 100
rect 360 80 520 90
rect 5040 80 5360 90
rect 6440 80 6840 90
rect 7400 80 8560 90
rect 9280 80 9320 90
rect 360 70 520 80
rect 5040 70 5360 80
rect 6440 70 6840 80
rect 7400 70 8560 80
rect 9280 70 9320 80
rect 360 60 520 70
rect 5040 60 5360 70
rect 6440 60 6840 70
rect 7400 60 8560 70
rect 9280 60 9320 70
rect 360 50 600 60
rect 5080 50 5360 60
rect 5680 50 5800 60
rect 6480 50 6840 60
rect 7360 50 8600 60
rect 8960 50 9000 60
rect 9240 50 9360 60
rect 360 40 600 50
rect 5080 40 5360 50
rect 5680 40 5800 50
rect 6480 40 6840 50
rect 7360 40 8600 50
rect 8960 40 9000 50
rect 9240 40 9360 50
rect 360 30 600 40
rect 5080 30 5360 40
rect 5680 30 5800 40
rect 6480 30 6840 40
rect 7360 30 8600 40
rect 8960 30 9000 40
rect 9240 30 9360 40
rect 360 20 600 30
rect 5080 20 5360 30
rect 5680 20 5800 30
rect 6480 20 6840 30
rect 7360 20 8600 30
rect 8960 20 9000 30
rect 9240 20 9360 30
rect 240 10 280 20
rect 360 10 600 20
rect 5080 10 5400 20
rect 5640 10 5840 20
rect 6480 10 6880 20
rect 7360 10 8560 20
rect 8920 10 9000 20
rect 9240 10 9400 20
rect 240 0 280 10
rect 360 0 600 10
rect 5080 0 5400 10
rect 5640 0 5840 10
rect 6480 0 6880 10
rect 7360 0 8560 10
rect 8920 0 9000 10
rect 9240 0 9400 10
<< metal1 >>
rect 2200 7490 2280 7500
rect 3640 7490 3680 7500
rect 9800 7490 9990 7500
rect 2200 7480 2280 7490
rect 3640 7480 3680 7490
rect 9800 7480 9990 7490
rect 2200 7470 2280 7480
rect 3640 7470 3680 7480
rect 9800 7470 9990 7480
rect 2200 7460 2280 7470
rect 3640 7460 3680 7470
rect 9800 7460 9990 7470
rect 2160 7450 2200 7460
rect 9760 7450 9800 7460
rect 9920 7450 9960 7460
rect 2160 7440 2200 7450
rect 9760 7440 9800 7450
rect 9920 7440 9960 7450
rect 2160 7430 2200 7440
rect 9760 7430 9800 7440
rect 9920 7430 9960 7440
rect 2160 7420 2200 7430
rect 9760 7420 9800 7430
rect 9920 7420 9960 7430
rect 2120 7410 2160 7420
rect 9680 7410 9760 7420
rect 9840 7410 9920 7420
rect 2120 7400 2160 7410
rect 9680 7400 9760 7410
rect 9840 7400 9920 7410
rect 2120 7390 2160 7400
rect 9680 7390 9760 7400
rect 9840 7390 9920 7400
rect 2120 7380 2160 7390
rect 9680 7380 9760 7390
rect 9840 7380 9920 7390
rect 2080 7370 2120 7380
rect 9640 7370 9990 7380
rect 2080 7360 2120 7370
rect 9640 7360 9990 7370
rect 2080 7350 2120 7360
rect 9640 7350 9990 7360
rect 2080 7340 2120 7350
rect 9640 7340 9990 7350
rect 2040 7330 2080 7340
rect 3320 7330 3360 7340
rect 9640 7330 9840 7340
rect 9880 7330 9960 7340
rect 2040 7320 2080 7330
rect 3320 7320 3360 7330
rect 9640 7320 9840 7330
rect 9880 7320 9960 7330
rect 2040 7310 2080 7320
rect 3320 7310 3360 7320
rect 9640 7310 9840 7320
rect 9880 7310 9960 7320
rect 2040 7300 2080 7310
rect 3320 7300 3360 7310
rect 9640 7300 9840 7310
rect 9880 7300 9960 7310
rect 2040 7290 2080 7300
rect 2520 7290 2560 7300
rect 3320 7290 3360 7300
rect 9880 7290 9960 7300
rect 2040 7280 2080 7290
rect 2520 7280 2560 7290
rect 3320 7280 3360 7290
rect 9880 7280 9960 7290
rect 2040 7270 2080 7280
rect 2520 7270 2560 7280
rect 3320 7270 3360 7280
rect 9880 7270 9960 7280
rect 2040 7260 2080 7270
rect 2520 7260 2560 7270
rect 3320 7260 3360 7270
rect 9880 7260 9960 7270
rect 2000 7250 2040 7260
rect 2440 7250 2560 7260
rect 3320 7250 3360 7260
rect 9880 7250 9960 7260
rect 2000 7240 2040 7250
rect 2440 7240 2560 7250
rect 3320 7240 3360 7250
rect 9880 7240 9960 7250
rect 2000 7230 2040 7240
rect 2440 7230 2560 7240
rect 3320 7230 3360 7240
rect 9880 7230 9960 7240
rect 2000 7220 2040 7230
rect 2440 7220 2560 7230
rect 3320 7220 3360 7230
rect 9880 7220 9960 7230
rect 2000 7210 2040 7220
rect 2120 7210 2280 7220
rect 2400 7210 2440 7220
rect 3320 7210 3400 7220
rect 3840 7210 3880 7220
rect 9840 7210 9960 7220
rect 2000 7200 2040 7210
rect 2120 7200 2280 7210
rect 2400 7200 2440 7210
rect 3320 7200 3400 7210
rect 3840 7200 3880 7210
rect 9840 7200 9960 7210
rect 2000 7190 2040 7200
rect 2120 7190 2280 7200
rect 2400 7190 2440 7200
rect 3320 7190 3400 7200
rect 3840 7190 3880 7200
rect 9840 7190 9960 7200
rect 2000 7180 2040 7190
rect 2120 7180 2280 7190
rect 2400 7180 2440 7190
rect 3320 7180 3400 7190
rect 3840 7180 3880 7190
rect 9840 7180 9960 7190
rect 1960 7170 2000 7180
rect 2080 7170 2320 7180
rect 3320 7170 3360 7180
rect 3840 7170 3880 7180
rect 9840 7170 9990 7180
rect 1960 7160 2000 7170
rect 2080 7160 2320 7170
rect 3320 7160 3360 7170
rect 3840 7160 3880 7170
rect 9840 7160 9990 7170
rect 1960 7150 2000 7160
rect 2080 7150 2320 7160
rect 3320 7150 3360 7160
rect 3840 7150 3880 7160
rect 9840 7150 9990 7160
rect 1960 7140 2000 7150
rect 2080 7140 2320 7150
rect 3320 7140 3360 7150
rect 3840 7140 3880 7150
rect 9840 7140 9990 7150
rect 1960 7130 2000 7140
rect 2040 7130 2200 7140
rect 3840 7130 3880 7140
rect 9680 7130 9720 7140
rect 9840 7130 9880 7140
rect 9920 7130 9990 7140
rect 1960 7120 2000 7130
rect 2040 7120 2200 7130
rect 3840 7120 3880 7130
rect 9680 7120 9720 7130
rect 9840 7120 9880 7130
rect 9920 7120 9990 7130
rect 1960 7110 2000 7120
rect 2040 7110 2200 7120
rect 3840 7110 3880 7120
rect 9680 7110 9720 7120
rect 9840 7110 9880 7120
rect 9920 7110 9990 7120
rect 1960 7100 2000 7110
rect 2040 7100 2200 7110
rect 3840 7100 3880 7110
rect 9680 7100 9720 7110
rect 9840 7100 9880 7110
rect 9920 7100 9990 7110
rect 1920 7090 2040 7100
rect 2120 7090 2160 7100
rect 3400 7090 3480 7100
rect 3640 7090 3680 7100
rect 9680 7090 9720 7100
rect 9800 7090 9840 7100
rect 9960 7090 9990 7100
rect 1920 7080 2040 7090
rect 2120 7080 2160 7090
rect 3400 7080 3480 7090
rect 3640 7080 3680 7090
rect 9680 7080 9720 7090
rect 9800 7080 9840 7090
rect 9960 7080 9990 7090
rect 1920 7070 2040 7080
rect 2120 7070 2160 7080
rect 3400 7070 3480 7080
rect 3640 7070 3680 7080
rect 9680 7070 9720 7080
rect 9800 7070 9840 7080
rect 9960 7070 9990 7080
rect 1920 7060 2040 7070
rect 2120 7060 2160 7070
rect 3400 7060 3480 7070
rect 3640 7060 3680 7070
rect 9680 7060 9720 7070
rect 9800 7060 9840 7070
rect 9960 7060 9990 7070
rect 1960 7050 2000 7060
rect 2080 7050 2120 7060
rect 2200 7050 3080 7060
rect 3440 7050 3520 7060
rect 3640 7050 3680 7060
rect 9680 7050 9800 7060
rect 9920 7050 9990 7060
rect 1960 7040 2000 7050
rect 2080 7040 2120 7050
rect 2200 7040 3080 7050
rect 3440 7040 3520 7050
rect 3640 7040 3680 7050
rect 9680 7040 9800 7050
rect 9920 7040 9990 7050
rect 1960 7030 2000 7040
rect 2080 7030 2120 7040
rect 2200 7030 3080 7040
rect 3440 7030 3520 7040
rect 3640 7030 3680 7040
rect 9680 7030 9800 7040
rect 9920 7030 9990 7040
rect 1960 7020 2000 7030
rect 2080 7020 2120 7030
rect 2200 7020 3080 7030
rect 3440 7020 3520 7030
rect 3640 7020 3680 7030
rect 9680 7020 9800 7030
rect 9920 7020 9990 7030
rect 2000 7010 2040 7020
rect 2160 7010 2240 7020
rect 2440 7010 2720 7020
rect 3200 7010 3240 7020
rect 3480 7010 3560 7020
rect 9680 7010 9720 7020
rect 9760 7010 9990 7020
rect 2000 7000 2040 7010
rect 2160 7000 2240 7010
rect 2440 7000 2720 7010
rect 3200 7000 3240 7010
rect 3480 7000 3560 7010
rect 9680 7000 9720 7010
rect 9760 7000 9990 7010
rect 2000 6990 2040 7000
rect 2160 6990 2240 7000
rect 2440 6990 2720 7000
rect 3200 6990 3240 7000
rect 3480 6990 3560 7000
rect 9680 6990 9720 7000
rect 9760 6990 9990 7000
rect 2000 6980 2040 6990
rect 2160 6980 2240 6990
rect 2440 6980 2720 6990
rect 3200 6980 3240 6990
rect 3480 6980 3560 6990
rect 9680 6980 9720 6990
rect 9760 6980 9990 6990
rect 2160 6970 2280 6980
rect 3320 6970 3360 6980
rect 3520 6970 3640 6980
rect 9640 6970 9680 6980
rect 9720 6970 9880 6980
rect 2160 6960 2280 6970
rect 3320 6960 3360 6970
rect 3520 6960 3640 6970
rect 9640 6960 9680 6970
rect 9720 6960 9880 6970
rect 2160 6950 2280 6960
rect 3320 6950 3360 6960
rect 3520 6950 3640 6960
rect 9640 6950 9680 6960
rect 9720 6950 9880 6960
rect 2160 6940 2280 6950
rect 3320 6940 3360 6950
rect 3520 6940 3640 6950
rect 9640 6940 9680 6950
rect 9720 6940 9880 6950
rect 1920 6930 1960 6940
rect 2200 6930 2320 6940
rect 3440 6930 3480 6940
rect 3560 6930 3720 6940
rect 9680 6930 9840 6940
rect 1920 6920 1960 6930
rect 2200 6920 2320 6930
rect 3440 6920 3480 6930
rect 3560 6920 3720 6930
rect 9680 6920 9840 6930
rect 1920 6910 1960 6920
rect 2200 6910 2320 6920
rect 3440 6910 3480 6920
rect 3560 6910 3720 6920
rect 9680 6910 9840 6920
rect 1920 6900 1960 6910
rect 2200 6900 2320 6910
rect 3440 6900 3480 6910
rect 3560 6900 3720 6910
rect 9680 6900 9840 6910
rect 2240 6890 2400 6900
rect 3520 6890 3560 6900
rect 3640 6890 3760 6900
rect 9680 6890 9880 6900
rect 2240 6880 2400 6890
rect 3520 6880 3560 6890
rect 3640 6880 3760 6890
rect 9680 6880 9880 6890
rect 2240 6870 2400 6880
rect 3520 6870 3560 6880
rect 3640 6870 3760 6880
rect 9680 6870 9880 6880
rect 2240 6860 2400 6870
rect 3520 6860 3560 6870
rect 3640 6860 3760 6870
rect 9680 6860 9880 6870
rect 2280 6850 2480 6860
rect 3680 6850 3800 6860
rect 9680 6850 9880 6860
rect 9920 6850 9990 6860
rect 2280 6840 2480 6850
rect 3680 6840 3800 6850
rect 9680 6840 9880 6850
rect 9920 6840 9990 6850
rect 2280 6830 2480 6840
rect 3680 6830 3800 6840
rect 9680 6830 9880 6840
rect 9920 6830 9990 6840
rect 2280 6820 2480 6830
rect 3680 6820 3800 6830
rect 9680 6820 9880 6830
rect 9920 6820 9990 6830
rect 1880 6810 1920 6820
rect 1960 6810 2040 6820
rect 2280 6810 2560 6820
rect 3720 6810 3840 6820
rect 9680 6810 9880 6820
rect 9920 6810 9990 6820
rect 1880 6800 1920 6810
rect 1960 6800 2040 6810
rect 2280 6800 2560 6810
rect 3720 6800 3840 6810
rect 9680 6800 9880 6810
rect 9920 6800 9990 6810
rect 1880 6790 1920 6800
rect 1960 6790 2040 6800
rect 2280 6790 2560 6800
rect 3720 6790 3840 6800
rect 9680 6790 9880 6800
rect 9920 6790 9990 6800
rect 1880 6780 1920 6790
rect 1960 6780 2040 6790
rect 2280 6780 2560 6790
rect 3720 6780 3840 6790
rect 9680 6780 9880 6790
rect 9920 6780 9990 6790
rect 1880 6770 1960 6780
rect 2000 6770 2040 6780
rect 2240 6770 2280 6780
rect 2520 6770 2600 6780
rect 2640 6770 2840 6780
rect 3720 6770 3760 6780
rect 3800 6770 3840 6780
rect 9600 6770 9640 6780
rect 9680 6770 9840 6780
rect 9960 6770 9990 6780
rect 1880 6760 1960 6770
rect 2000 6760 2040 6770
rect 2240 6760 2280 6770
rect 2520 6760 2600 6770
rect 2640 6760 2840 6770
rect 3720 6760 3760 6770
rect 3800 6760 3840 6770
rect 9600 6760 9640 6770
rect 9680 6760 9840 6770
rect 9960 6760 9990 6770
rect 1880 6750 1960 6760
rect 2000 6750 2040 6760
rect 2240 6750 2280 6760
rect 2520 6750 2600 6760
rect 2640 6750 2840 6760
rect 3720 6750 3760 6760
rect 3800 6750 3840 6760
rect 9600 6750 9640 6760
rect 9680 6750 9840 6760
rect 9960 6750 9990 6760
rect 1880 6740 1960 6750
rect 2000 6740 2040 6750
rect 2240 6740 2280 6750
rect 2520 6740 2600 6750
rect 2640 6740 2840 6750
rect 3720 6740 3760 6750
rect 3800 6740 3840 6750
rect 9600 6740 9640 6750
rect 9680 6740 9840 6750
rect 9960 6740 9990 6750
rect 1880 6730 2000 6740
rect 2200 6730 2240 6740
rect 2520 6730 2560 6740
rect 3000 6730 3160 6740
rect 3840 6730 3880 6740
rect 9600 6730 9640 6740
rect 9680 6730 9840 6740
rect 1880 6720 2000 6730
rect 2200 6720 2240 6730
rect 2520 6720 2560 6730
rect 3000 6720 3160 6730
rect 3840 6720 3880 6730
rect 9600 6720 9640 6730
rect 9680 6720 9840 6730
rect 1880 6710 2000 6720
rect 2200 6710 2240 6720
rect 2520 6710 2560 6720
rect 3000 6710 3160 6720
rect 3840 6710 3880 6720
rect 9600 6710 9640 6720
rect 9680 6710 9840 6720
rect 1880 6700 2000 6710
rect 2200 6700 2240 6710
rect 2520 6700 2560 6710
rect 3000 6700 3160 6710
rect 3840 6700 3880 6710
rect 9600 6700 9640 6710
rect 9680 6700 9840 6710
rect 1880 6690 1960 6700
rect 2200 6690 2240 6700
rect 2560 6690 2640 6700
rect 3280 6690 3400 6700
rect 3880 6690 3920 6700
rect 9600 6690 9640 6700
rect 9680 6690 9840 6700
rect 9880 6690 9920 6700
rect 1880 6680 1960 6690
rect 2200 6680 2240 6690
rect 2560 6680 2640 6690
rect 3280 6680 3400 6690
rect 3880 6680 3920 6690
rect 9600 6680 9640 6690
rect 9680 6680 9840 6690
rect 9880 6680 9920 6690
rect 1880 6670 1960 6680
rect 2200 6670 2240 6680
rect 2560 6670 2640 6680
rect 3280 6670 3400 6680
rect 3880 6670 3920 6680
rect 9600 6670 9640 6680
rect 9680 6670 9840 6680
rect 9880 6670 9920 6680
rect 1880 6660 1960 6670
rect 2200 6660 2240 6670
rect 2560 6660 2640 6670
rect 3280 6660 3400 6670
rect 3880 6660 3920 6670
rect 9600 6660 9640 6670
rect 9680 6660 9840 6670
rect 9880 6660 9920 6670
rect 1840 6650 1920 6660
rect 2600 6650 2680 6660
rect 3480 6650 3520 6660
rect 9680 6650 9800 6660
rect 1840 6640 1920 6650
rect 2600 6640 2680 6650
rect 3480 6640 3520 6650
rect 9680 6640 9800 6650
rect 1840 6630 1920 6640
rect 2600 6630 2680 6640
rect 3480 6630 3520 6640
rect 9680 6630 9800 6640
rect 1840 6620 1920 6630
rect 2600 6620 2680 6630
rect 3480 6620 3520 6630
rect 9680 6620 9800 6630
rect 1760 6610 1800 6620
rect 2120 6610 2160 6620
rect 2640 6610 2680 6620
rect 3600 6610 3640 6620
rect 3920 6610 3960 6620
rect 1760 6600 1800 6610
rect 2120 6600 2160 6610
rect 2640 6600 2680 6610
rect 3600 6600 3640 6610
rect 3920 6600 3960 6610
rect 1760 6590 1800 6600
rect 2120 6590 2160 6600
rect 2640 6590 2680 6600
rect 3600 6590 3640 6600
rect 3920 6590 3960 6600
rect 1760 6580 1800 6590
rect 2120 6580 2160 6590
rect 2640 6580 2680 6590
rect 3600 6580 3640 6590
rect 3920 6580 3960 6590
rect 1560 6570 1600 6580
rect 1800 6570 1840 6580
rect 2000 6570 2040 6580
rect 2640 6570 2680 6580
rect 1560 6560 1600 6570
rect 1800 6560 1840 6570
rect 2000 6560 2040 6570
rect 2640 6560 2680 6570
rect 1560 6550 1600 6560
rect 1800 6550 1840 6560
rect 2000 6550 2040 6560
rect 2640 6550 2680 6560
rect 1560 6540 1600 6550
rect 1800 6540 1840 6550
rect 2000 6540 2040 6550
rect 2640 6540 2680 6550
rect 1440 6530 1520 6540
rect 1560 6530 1640 6540
rect 1720 6530 1760 6540
rect 1840 6530 1880 6540
rect 2600 6530 2640 6540
rect 3960 6530 4000 6540
rect 1440 6520 1520 6530
rect 1560 6520 1640 6530
rect 1720 6520 1760 6530
rect 1840 6520 1880 6530
rect 2600 6520 2640 6530
rect 3960 6520 4000 6530
rect 1440 6510 1520 6520
rect 1560 6510 1640 6520
rect 1720 6510 1760 6520
rect 1840 6510 1880 6520
rect 2600 6510 2640 6520
rect 3960 6510 4000 6520
rect 1440 6500 1520 6510
rect 1560 6500 1640 6510
rect 1720 6500 1760 6510
rect 1840 6500 1880 6510
rect 2600 6500 2640 6510
rect 3960 6500 4000 6510
rect 1280 6490 1320 6500
rect 1360 6490 1400 6500
rect 1520 6490 1600 6500
rect 1640 6490 1680 6500
rect 1760 6490 1800 6500
rect 1840 6490 1960 6500
rect 2080 6490 2120 6500
rect 2400 6490 2520 6500
rect 2560 6490 2600 6500
rect 6400 6490 6520 6500
rect 9880 6490 9990 6500
rect 1280 6480 1320 6490
rect 1360 6480 1400 6490
rect 1520 6480 1600 6490
rect 1640 6480 1680 6490
rect 1760 6480 1800 6490
rect 1840 6480 1960 6490
rect 2080 6480 2120 6490
rect 2400 6480 2520 6490
rect 2560 6480 2600 6490
rect 6400 6480 6520 6490
rect 9880 6480 9990 6490
rect 1280 6470 1320 6480
rect 1360 6470 1400 6480
rect 1520 6470 1600 6480
rect 1640 6470 1680 6480
rect 1760 6470 1800 6480
rect 1840 6470 1960 6480
rect 2080 6470 2120 6480
rect 2400 6470 2520 6480
rect 2560 6470 2600 6480
rect 6400 6470 6520 6480
rect 9880 6470 9990 6480
rect 1280 6460 1320 6470
rect 1360 6460 1400 6470
rect 1520 6460 1600 6470
rect 1640 6460 1680 6470
rect 1760 6460 1800 6470
rect 1840 6460 1960 6470
rect 2080 6460 2120 6470
rect 2400 6460 2520 6470
rect 2560 6460 2600 6470
rect 6400 6460 6520 6470
rect 9880 6460 9990 6470
rect 1240 6450 1280 6460
rect 1360 6450 1400 6460
rect 1440 6450 1480 6460
rect 1560 6450 1640 6460
rect 1960 6450 2080 6460
rect 2480 6450 2520 6460
rect 3920 6450 3960 6460
rect 6120 6450 6200 6460
rect 6400 6450 6560 6460
rect 9760 6450 9840 6460
rect 9920 6450 9990 6460
rect 1240 6440 1280 6450
rect 1360 6440 1400 6450
rect 1440 6440 1480 6450
rect 1560 6440 1640 6450
rect 1960 6440 2080 6450
rect 2480 6440 2520 6450
rect 3920 6440 3960 6450
rect 6120 6440 6200 6450
rect 6400 6440 6560 6450
rect 9760 6440 9840 6450
rect 9920 6440 9990 6450
rect 1240 6430 1280 6440
rect 1360 6430 1400 6440
rect 1440 6430 1480 6440
rect 1560 6430 1640 6440
rect 1960 6430 2080 6440
rect 2480 6430 2520 6440
rect 3920 6430 3960 6440
rect 6120 6430 6200 6440
rect 6400 6430 6560 6440
rect 9760 6430 9840 6440
rect 9920 6430 9990 6440
rect 1240 6420 1280 6430
rect 1360 6420 1400 6430
rect 1440 6420 1480 6430
rect 1560 6420 1640 6430
rect 1960 6420 2080 6430
rect 2480 6420 2520 6430
rect 3920 6420 3960 6430
rect 6120 6420 6200 6430
rect 6400 6420 6560 6430
rect 9760 6420 9840 6430
rect 9920 6420 9990 6430
rect 1560 6410 1600 6420
rect 6400 6410 6600 6420
rect 9640 6410 9800 6420
rect 1560 6400 1600 6410
rect 6400 6400 6600 6410
rect 9640 6400 9800 6410
rect 1560 6390 1600 6400
rect 6400 6390 6600 6400
rect 9640 6390 9800 6400
rect 1560 6380 1600 6390
rect 6400 6380 6600 6390
rect 9640 6380 9800 6390
rect 1440 6370 1480 6380
rect 1560 6370 1600 6380
rect 1720 6370 1760 6380
rect 1800 6370 1840 6380
rect 2400 6370 2480 6380
rect 4040 6370 4080 6380
rect 6440 6370 6600 6380
rect 9640 6370 9880 6380
rect 9920 6370 9990 6380
rect 1440 6360 1480 6370
rect 1560 6360 1600 6370
rect 1720 6360 1760 6370
rect 1800 6360 1840 6370
rect 2400 6360 2480 6370
rect 4040 6360 4080 6370
rect 6440 6360 6600 6370
rect 9640 6360 9880 6370
rect 9920 6360 9990 6370
rect 1440 6350 1480 6360
rect 1560 6350 1600 6360
rect 1720 6350 1760 6360
rect 1800 6350 1840 6360
rect 2400 6350 2480 6360
rect 4040 6350 4080 6360
rect 6440 6350 6600 6360
rect 9640 6350 9880 6360
rect 9920 6350 9990 6360
rect 1440 6340 1480 6350
rect 1560 6340 1600 6350
rect 1720 6340 1760 6350
rect 1800 6340 1840 6350
rect 2400 6340 2480 6350
rect 4040 6340 4080 6350
rect 6440 6340 6600 6350
rect 9640 6340 9880 6350
rect 9920 6340 9990 6350
rect 1680 6330 1720 6340
rect 1800 6330 1840 6340
rect 6520 6330 6720 6340
rect 9640 6330 9720 6340
rect 9760 6330 9840 6340
rect 9920 6330 9990 6340
rect 1680 6320 1720 6330
rect 1800 6320 1840 6330
rect 6520 6320 6720 6330
rect 9640 6320 9720 6330
rect 9760 6320 9840 6330
rect 9920 6320 9990 6330
rect 1680 6310 1720 6320
rect 1800 6310 1840 6320
rect 6520 6310 6720 6320
rect 9640 6310 9720 6320
rect 9760 6310 9840 6320
rect 9920 6310 9990 6320
rect 1680 6300 1720 6310
rect 1800 6300 1840 6310
rect 6520 6300 6720 6310
rect 9640 6300 9720 6310
rect 9760 6300 9840 6310
rect 9920 6300 9990 6310
rect 1520 6290 1560 6300
rect 1640 6290 1720 6300
rect 1760 6290 1800 6300
rect 5400 6290 5440 6300
rect 5480 6290 5520 6300
rect 6600 6290 6760 6300
rect 9640 6290 9680 6300
rect 9800 6290 9840 6300
rect 1520 6280 1560 6290
rect 1640 6280 1720 6290
rect 1760 6280 1800 6290
rect 5400 6280 5440 6290
rect 5480 6280 5520 6290
rect 6600 6280 6760 6290
rect 9640 6280 9680 6290
rect 9800 6280 9840 6290
rect 1520 6270 1560 6280
rect 1640 6270 1720 6280
rect 1760 6270 1800 6280
rect 5400 6270 5440 6280
rect 5480 6270 5520 6280
rect 6600 6270 6760 6280
rect 9640 6270 9680 6280
rect 9800 6270 9840 6280
rect 1520 6260 1560 6270
rect 1640 6260 1720 6270
rect 1760 6260 1800 6270
rect 5400 6260 5440 6270
rect 5480 6260 5520 6270
rect 6600 6260 6760 6270
rect 9640 6260 9680 6270
rect 9800 6260 9840 6270
rect 1600 6250 1680 6260
rect 1720 6250 1800 6260
rect 2440 6250 2480 6260
rect 5360 6250 5400 6260
rect 5480 6250 5520 6260
rect 6640 6250 6760 6260
rect 9520 6250 9600 6260
rect 1600 6240 1680 6250
rect 1720 6240 1800 6250
rect 2440 6240 2480 6250
rect 5360 6240 5400 6250
rect 5480 6240 5520 6250
rect 6640 6240 6760 6250
rect 9520 6240 9600 6250
rect 1600 6230 1680 6240
rect 1720 6230 1800 6240
rect 2440 6230 2480 6240
rect 5360 6230 5400 6240
rect 5480 6230 5520 6240
rect 6640 6230 6760 6240
rect 9520 6230 9600 6240
rect 1600 6220 1680 6230
rect 1720 6220 1800 6230
rect 2440 6220 2480 6230
rect 5360 6220 5400 6230
rect 5480 6220 5520 6230
rect 6640 6220 6760 6230
rect 9520 6220 9600 6230
rect 1560 6210 1600 6220
rect 1640 6210 1720 6220
rect 5320 6210 5360 6220
rect 5440 6210 5480 6220
rect 6680 6210 6760 6220
rect 9400 6210 9440 6220
rect 9680 6210 9720 6220
rect 9760 6210 9800 6220
rect 1560 6200 1600 6210
rect 1640 6200 1720 6210
rect 5320 6200 5360 6210
rect 5440 6200 5480 6210
rect 6680 6200 6760 6210
rect 9400 6200 9440 6210
rect 9680 6200 9720 6210
rect 9760 6200 9800 6210
rect 1560 6190 1600 6200
rect 1640 6190 1720 6200
rect 5320 6190 5360 6200
rect 5440 6190 5480 6200
rect 6680 6190 6760 6200
rect 9400 6190 9440 6200
rect 9680 6190 9720 6200
rect 9760 6190 9800 6200
rect 1560 6180 1600 6190
rect 1640 6180 1720 6190
rect 5320 6180 5360 6190
rect 5440 6180 5480 6190
rect 6680 6180 6760 6190
rect 9400 6180 9440 6190
rect 9680 6180 9720 6190
rect 9760 6180 9800 6190
rect 1680 6170 1720 6180
rect 4240 6170 4280 6180
rect 5400 6170 5440 6180
rect 6680 6170 6760 6180
rect 9280 6170 9480 6180
rect 9680 6170 9720 6180
rect 1680 6160 1720 6170
rect 4240 6160 4280 6170
rect 5400 6160 5440 6170
rect 6680 6160 6760 6170
rect 9280 6160 9480 6170
rect 9680 6160 9720 6170
rect 1680 6150 1720 6160
rect 4240 6150 4280 6160
rect 5400 6150 5440 6160
rect 6680 6150 6760 6160
rect 9280 6150 9480 6160
rect 9680 6150 9720 6160
rect 1680 6140 1720 6150
rect 4240 6140 4280 6150
rect 5400 6140 5440 6150
rect 6680 6140 6760 6150
rect 9280 6140 9480 6150
rect 9680 6140 9720 6150
rect 1360 6130 1400 6140
rect 1600 6130 1640 6140
rect 5280 6130 5320 6140
rect 5360 6130 5400 6140
rect 6720 6130 6840 6140
rect 9200 6130 9280 6140
rect 9320 6130 9400 6140
rect 9440 6130 9480 6140
rect 9640 6130 9720 6140
rect 9800 6130 9840 6140
rect 1360 6120 1400 6130
rect 1600 6120 1640 6130
rect 5280 6120 5320 6130
rect 5360 6120 5400 6130
rect 6720 6120 6840 6130
rect 9200 6120 9280 6130
rect 9320 6120 9400 6130
rect 9440 6120 9480 6130
rect 9640 6120 9720 6130
rect 9800 6120 9840 6130
rect 1360 6110 1400 6120
rect 1600 6110 1640 6120
rect 5280 6110 5320 6120
rect 5360 6110 5400 6120
rect 6720 6110 6840 6120
rect 9200 6110 9280 6120
rect 9320 6110 9400 6120
rect 9440 6110 9480 6120
rect 9640 6110 9720 6120
rect 9800 6110 9840 6120
rect 1360 6100 1400 6110
rect 1600 6100 1640 6110
rect 5280 6100 5320 6110
rect 5360 6100 5400 6110
rect 6720 6100 6840 6110
rect 9200 6100 9280 6110
rect 9320 6100 9400 6110
rect 9440 6100 9480 6110
rect 9640 6100 9720 6110
rect 9800 6100 9840 6110
rect 1320 6090 1440 6100
rect 1600 6090 1640 6100
rect 3760 6090 3840 6100
rect 4280 6090 4320 6100
rect 6760 6090 6840 6100
rect 9120 6090 9280 6100
rect 9640 6090 9720 6100
rect 1320 6080 1440 6090
rect 1600 6080 1640 6090
rect 3760 6080 3840 6090
rect 4280 6080 4320 6090
rect 6760 6080 6840 6090
rect 9120 6080 9280 6090
rect 9640 6080 9720 6090
rect 1320 6070 1440 6080
rect 1600 6070 1640 6080
rect 3760 6070 3840 6080
rect 4280 6070 4320 6080
rect 6760 6070 6840 6080
rect 9120 6070 9280 6080
rect 9640 6070 9720 6080
rect 1320 6060 1440 6070
rect 1600 6060 1640 6070
rect 3760 6060 3840 6070
rect 4280 6060 4320 6070
rect 6760 6060 6840 6070
rect 9120 6060 9280 6070
rect 9640 6060 9720 6070
rect 1320 6050 1360 6060
rect 3200 6050 3280 6060
rect 6760 6050 6800 6060
rect 9040 6050 9160 6060
rect 9640 6050 9720 6060
rect 1320 6040 1360 6050
rect 3200 6040 3280 6050
rect 6760 6040 6800 6050
rect 9040 6040 9160 6050
rect 9640 6040 9720 6050
rect 1320 6030 1360 6040
rect 3200 6030 3280 6040
rect 6760 6030 6800 6040
rect 9040 6030 9160 6040
rect 9640 6030 9720 6040
rect 1320 6020 1360 6030
rect 3200 6020 3280 6030
rect 6760 6020 6800 6030
rect 9040 6020 9160 6030
rect 9640 6020 9720 6030
rect 1200 6010 1360 6020
rect 1600 6010 1680 6020
rect 3160 6010 3200 6020
rect 3240 6010 3280 6020
rect 5200 6010 5240 6020
rect 5320 6010 5360 6020
rect 6800 6010 6840 6020
rect 8840 6010 9040 6020
rect 9240 6010 9360 6020
rect 9640 6010 9720 6020
rect 9840 6010 9880 6020
rect 1200 6000 1360 6010
rect 1600 6000 1680 6010
rect 3160 6000 3200 6010
rect 3240 6000 3280 6010
rect 5200 6000 5240 6010
rect 5320 6000 5360 6010
rect 6800 6000 6840 6010
rect 8840 6000 9040 6010
rect 9240 6000 9360 6010
rect 9640 6000 9720 6010
rect 9840 6000 9880 6010
rect 1200 5990 1360 6000
rect 1600 5990 1680 6000
rect 3160 5990 3200 6000
rect 3240 5990 3280 6000
rect 5200 5990 5240 6000
rect 5320 5990 5360 6000
rect 6800 5990 6840 6000
rect 8840 5990 9040 6000
rect 9240 5990 9360 6000
rect 9640 5990 9720 6000
rect 9840 5990 9880 6000
rect 1200 5980 1360 5990
rect 1600 5980 1680 5990
rect 3160 5980 3200 5990
rect 3240 5980 3280 5990
rect 5200 5980 5240 5990
rect 5320 5980 5360 5990
rect 6800 5980 6840 5990
rect 8840 5980 9040 5990
rect 9240 5980 9360 5990
rect 9640 5980 9720 5990
rect 9840 5980 9880 5990
rect 1120 5970 1160 5980
rect 1240 5970 1280 5980
rect 1640 5970 1680 5980
rect 3120 5970 3160 5980
rect 3240 5970 3280 5980
rect 6840 5970 6960 5980
rect 8680 5970 8960 5980
rect 9320 5970 9360 5980
rect 9680 5970 9760 5980
rect 1120 5960 1160 5970
rect 1240 5960 1280 5970
rect 1640 5960 1680 5970
rect 3120 5960 3160 5970
rect 3240 5960 3280 5970
rect 6840 5960 6960 5970
rect 8680 5960 8960 5970
rect 9320 5960 9360 5970
rect 9680 5960 9760 5970
rect 1120 5950 1160 5960
rect 1240 5950 1280 5960
rect 1640 5950 1680 5960
rect 3120 5950 3160 5960
rect 3240 5950 3280 5960
rect 6840 5950 6960 5960
rect 8680 5950 8960 5960
rect 9320 5950 9360 5960
rect 9680 5950 9760 5960
rect 1120 5940 1160 5950
rect 1240 5940 1280 5950
rect 1640 5940 1680 5950
rect 3120 5940 3160 5950
rect 3240 5940 3280 5950
rect 6840 5940 6960 5950
rect 8680 5940 8960 5950
rect 9320 5940 9360 5950
rect 9680 5940 9760 5950
rect 960 5930 1080 5940
rect 1160 5930 1200 5940
rect 2560 5930 2600 5940
rect 3080 5930 3120 5940
rect 4200 5930 4240 5940
rect 4280 5930 4320 5940
rect 6840 5930 6960 5940
rect 8560 5930 8800 5940
rect 9280 5930 9360 5940
rect 9440 5930 9480 5940
rect 9680 5930 9760 5940
rect 960 5920 1080 5930
rect 1160 5920 1200 5930
rect 2560 5920 2600 5930
rect 3080 5920 3120 5930
rect 4200 5920 4240 5930
rect 4280 5920 4320 5930
rect 6840 5920 6960 5930
rect 8560 5920 8800 5930
rect 9280 5920 9360 5930
rect 9440 5920 9480 5930
rect 9680 5920 9760 5930
rect 960 5910 1080 5920
rect 1160 5910 1200 5920
rect 2560 5910 2600 5920
rect 3080 5910 3120 5920
rect 4200 5910 4240 5920
rect 4280 5910 4320 5920
rect 6840 5910 6960 5920
rect 8560 5910 8800 5920
rect 9280 5910 9360 5920
rect 9440 5910 9480 5920
rect 9680 5910 9760 5920
rect 960 5900 1080 5910
rect 1160 5900 1200 5910
rect 2560 5900 2600 5910
rect 3080 5900 3120 5910
rect 4200 5900 4240 5910
rect 4280 5900 4320 5910
rect 6840 5900 6960 5910
rect 8560 5900 8800 5910
rect 9280 5900 9360 5910
rect 9440 5900 9480 5910
rect 9680 5900 9760 5910
rect 1000 5890 1120 5900
rect 1720 5890 1760 5900
rect 2600 5890 2680 5900
rect 3000 5890 3080 5900
rect 3240 5890 3280 5900
rect 3720 5890 3760 5900
rect 6920 5890 6960 5900
rect 8440 5890 8600 5900
rect 8760 5890 8800 5900
rect 9360 5890 9440 5900
rect 9720 5890 9760 5900
rect 9880 5890 9920 5900
rect 1000 5880 1120 5890
rect 1720 5880 1760 5890
rect 2600 5880 2680 5890
rect 3000 5880 3080 5890
rect 3240 5880 3280 5890
rect 3720 5880 3760 5890
rect 6920 5880 6960 5890
rect 8440 5880 8600 5890
rect 8760 5880 8800 5890
rect 9360 5880 9440 5890
rect 9720 5880 9760 5890
rect 9880 5880 9920 5890
rect 1000 5870 1120 5880
rect 1720 5870 1760 5880
rect 2600 5870 2680 5880
rect 3000 5870 3080 5880
rect 3240 5870 3280 5880
rect 3720 5870 3760 5880
rect 6920 5870 6960 5880
rect 8440 5870 8600 5880
rect 8760 5870 8800 5880
rect 9360 5870 9440 5880
rect 9720 5870 9760 5880
rect 9880 5870 9920 5880
rect 1000 5860 1120 5870
rect 1720 5860 1760 5870
rect 2600 5860 2680 5870
rect 3000 5860 3080 5870
rect 3240 5860 3280 5870
rect 3720 5860 3760 5870
rect 6920 5860 6960 5870
rect 8440 5860 8600 5870
rect 8760 5860 8800 5870
rect 9360 5860 9440 5870
rect 9720 5860 9760 5870
rect 9880 5860 9920 5870
rect 680 5850 720 5860
rect 800 5850 880 5860
rect 960 5850 1000 5860
rect 2680 5850 2720 5860
rect 2840 5850 2960 5860
rect 5280 5850 5320 5860
rect 6920 5850 6960 5860
rect 8280 5850 8600 5860
rect 8720 5850 8800 5860
rect 9280 5850 9360 5860
rect 9880 5850 9920 5860
rect 680 5840 720 5850
rect 800 5840 880 5850
rect 960 5840 1000 5850
rect 2680 5840 2720 5850
rect 2840 5840 2960 5850
rect 5280 5840 5320 5850
rect 6920 5840 6960 5850
rect 8280 5840 8600 5850
rect 8720 5840 8800 5850
rect 9280 5840 9360 5850
rect 9880 5840 9920 5850
rect 680 5830 720 5840
rect 800 5830 880 5840
rect 960 5830 1000 5840
rect 2680 5830 2720 5840
rect 2840 5830 2960 5840
rect 5280 5830 5320 5840
rect 6920 5830 6960 5840
rect 8280 5830 8600 5840
rect 8720 5830 8800 5840
rect 9280 5830 9360 5840
rect 9880 5830 9920 5840
rect 680 5820 720 5830
rect 800 5820 880 5830
rect 960 5820 1000 5830
rect 2680 5820 2720 5830
rect 2840 5820 2960 5830
rect 5280 5820 5320 5830
rect 6920 5820 6960 5830
rect 8280 5820 8600 5830
rect 8720 5820 8800 5830
rect 9280 5820 9360 5830
rect 9880 5820 9920 5830
rect 880 5810 920 5820
rect 2680 5810 2840 5820
rect 3280 5810 3320 5820
rect 3720 5810 3760 5820
rect 5280 5810 5320 5820
rect 6840 5810 6880 5820
rect 6920 5810 6960 5820
rect 8160 5810 8400 5820
rect 8440 5810 8680 5820
rect 8760 5810 8800 5820
rect 8960 5810 9000 5820
rect 9080 5810 9280 5820
rect 880 5800 920 5810
rect 2680 5800 2840 5810
rect 3280 5800 3320 5810
rect 3720 5800 3760 5810
rect 5280 5800 5320 5810
rect 6840 5800 6880 5810
rect 6920 5800 6960 5810
rect 8160 5800 8400 5810
rect 8440 5800 8680 5810
rect 8760 5800 8800 5810
rect 8960 5800 9000 5810
rect 9080 5800 9280 5810
rect 880 5790 920 5800
rect 2680 5790 2840 5800
rect 3280 5790 3320 5800
rect 3720 5790 3760 5800
rect 5280 5790 5320 5800
rect 6840 5790 6880 5800
rect 6920 5790 6960 5800
rect 8160 5790 8400 5800
rect 8440 5790 8680 5800
rect 8760 5790 8800 5800
rect 8960 5790 9000 5800
rect 9080 5790 9280 5800
rect 880 5780 920 5790
rect 2680 5780 2840 5790
rect 3280 5780 3320 5790
rect 3720 5780 3760 5790
rect 5280 5780 5320 5790
rect 6840 5780 6880 5790
rect 6920 5780 6960 5790
rect 8160 5780 8400 5790
rect 8440 5780 8680 5790
rect 8760 5780 8800 5790
rect 8960 5780 9000 5790
rect 9080 5780 9280 5790
rect 880 5770 920 5780
rect 1840 5770 1880 5780
rect 2640 5770 2800 5780
rect 3280 5770 3320 5780
rect 3720 5770 3880 5780
rect 6840 5770 6960 5780
rect 8040 5770 8240 5780
rect 8280 5770 8360 5780
rect 8440 5770 8680 5780
rect 8760 5770 8800 5780
rect 8960 5770 9080 5780
rect 9160 5770 9200 5780
rect 880 5760 920 5770
rect 1840 5760 1880 5770
rect 2640 5760 2800 5770
rect 3280 5760 3320 5770
rect 3720 5760 3880 5770
rect 6840 5760 6960 5770
rect 8040 5760 8240 5770
rect 8280 5760 8360 5770
rect 8440 5760 8680 5770
rect 8760 5760 8800 5770
rect 8960 5760 9080 5770
rect 9160 5760 9200 5770
rect 880 5750 920 5760
rect 1840 5750 1880 5760
rect 2640 5750 2800 5760
rect 3280 5750 3320 5760
rect 3720 5750 3880 5760
rect 6840 5750 6960 5760
rect 8040 5750 8240 5760
rect 8280 5750 8360 5760
rect 8440 5750 8680 5760
rect 8760 5750 8800 5760
rect 8960 5750 9080 5760
rect 9160 5750 9200 5760
rect 880 5740 920 5750
rect 1840 5740 1880 5750
rect 2640 5740 2800 5750
rect 3280 5740 3320 5750
rect 3720 5740 3880 5750
rect 6840 5740 6960 5750
rect 8040 5740 8240 5750
rect 8280 5740 8360 5750
rect 8440 5740 8680 5750
rect 8760 5740 8800 5750
rect 8960 5740 9080 5750
rect 9160 5740 9200 5750
rect 800 5730 880 5740
rect 1160 5730 1240 5740
rect 1840 5730 1880 5740
rect 2240 5730 2280 5740
rect 2600 5730 2760 5740
rect 3280 5730 3320 5740
rect 3720 5730 3760 5740
rect 3840 5730 3880 5740
rect 3920 5730 4000 5740
rect 5080 5730 5120 5740
rect 6840 5730 6920 5740
rect 7920 5730 8120 5740
rect 8320 5730 8360 5740
rect 8440 5730 8680 5740
rect 8800 5730 9040 5740
rect 9920 5730 9960 5740
rect 800 5720 880 5730
rect 1160 5720 1240 5730
rect 1840 5720 1880 5730
rect 2240 5720 2280 5730
rect 2600 5720 2760 5730
rect 3280 5720 3320 5730
rect 3720 5720 3760 5730
rect 3840 5720 3880 5730
rect 3920 5720 4000 5730
rect 5080 5720 5120 5730
rect 6840 5720 6920 5730
rect 7920 5720 8120 5730
rect 8320 5720 8360 5730
rect 8440 5720 8680 5730
rect 8800 5720 9040 5730
rect 9920 5720 9960 5730
rect 800 5710 880 5720
rect 1160 5710 1240 5720
rect 1840 5710 1880 5720
rect 2240 5710 2280 5720
rect 2600 5710 2760 5720
rect 3280 5710 3320 5720
rect 3720 5710 3760 5720
rect 3840 5710 3880 5720
rect 3920 5710 4000 5720
rect 5080 5710 5120 5720
rect 6840 5710 6920 5720
rect 7920 5710 8120 5720
rect 8320 5710 8360 5720
rect 8440 5710 8680 5720
rect 8800 5710 9040 5720
rect 9920 5710 9960 5720
rect 800 5700 880 5710
rect 1160 5700 1240 5710
rect 1840 5700 1880 5710
rect 2240 5700 2280 5710
rect 2600 5700 2760 5710
rect 3280 5700 3320 5710
rect 3720 5700 3760 5710
rect 3840 5700 3880 5710
rect 3920 5700 4000 5710
rect 5080 5700 5120 5710
rect 6840 5700 6920 5710
rect 7920 5700 8120 5710
rect 8320 5700 8360 5710
rect 8440 5700 8680 5710
rect 8800 5700 9040 5710
rect 9920 5700 9960 5710
rect 1160 5690 1200 5700
rect 1840 5690 1880 5700
rect 2560 5690 2680 5700
rect 3280 5690 3320 5700
rect 3680 5690 3720 5700
rect 3760 5690 3880 5700
rect 3920 5690 4000 5700
rect 5120 5690 5160 5700
rect 6880 5690 6920 5700
rect 7760 5690 7800 5700
rect 7920 5690 8000 5700
rect 8320 5690 8400 5700
rect 8480 5690 8760 5700
rect 8920 5690 9000 5700
rect 9960 5690 9990 5700
rect 1160 5680 1200 5690
rect 1840 5680 1880 5690
rect 2560 5680 2680 5690
rect 3280 5680 3320 5690
rect 3680 5680 3720 5690
rect 3760 5680 3880 5690
rect 3920 5680 4000 5690
rect 5120 5680 5160 5690
rect 6880 5680 6920 5690
rect 7760 5680 7800 5690
rect 7920 5680 8000 5690
rect 8320 5680 8400 5690
rect 8480 5680 8760 5690
rect 8920 5680 9000 5690
rect 9960 5680 9990 5690
rect 1160 5670 1200 5680
rect 1840 5670 1880 5680
rect 2560 5670 2680 5680
rect 3280 5670 3320 5680
rect 3680 5670 3720 5680
rect 3760 5670 3880 5680
rect 3920 5670 4000 5680
rect 5120 5670 5160 5680
rect 6880 5670 6920 5680
rect 7760 5670 7800 5680
rect 7920 5670 8000 5680
rect 8320 5670 8400 5680
rect 8480 5670 8760 5680
rect 8920 5670 9000 5680
rect 9960 5670 9990 5680
rect 1160 5660 1200 5670
rect 1840 5660 1880 5670
rect 2560 5660 2680 5670
rect 3280 5660 3320 5670
rect 3680 5660 3720 5670
rect 3760 5660 3880 5670
rect 3920 5660 4000 5670
rect 5120 5660 5160 5670
rect 6880 5660 6920 5670
rect 7760 5660 7800 5670
rect 7920 5660 8000 5670
rect 8320 5660 8400 5670
rect 8480 5660 8760 5670
rect 8920 5660 9000 5670
rect 9960 5660 9990 5670
rect 800 5650 840 5660
rect 1840 5650 1880 5660
rect 2200 5650 2240 5660
rect 2520 5650 2640 5660
rect 3280 5650 3320 5660
rect 3680 5650 3720 5660
rect 3760 5650 3800 5660
rect 5120 5650 5160 5660
rect 5240 5650 5280 5660
rect 6920 5650 6960 5660
rect 7720 5650 7800 5660
rect 7920 5650 8000 5660
rect 8320 5650 8400 5660
rect 800 5640 840 5650
rect 1840 5640 1880 5650
rect 2200 5640 2240 5650
rect 2520 5640 2640 5650
rect 3280 5640 3320 5650
rect 3680 5640 3720 5650
rect 3760 5640 3800 5650
rect 5120 5640 5160 5650
rect 5240 5640 5280 5650
rect 6920 5640 6960 5650
rect 7720 5640 7800 5650
rect 7920 5640 8000 5650
rect 8320 5640 8400 5650
rect 800 5630 840 5640
rect 1840 5630 1880 5640
rect 2200 5630 2240 5640
rect 2520 5630 2640 5640
rect 3280 5630 3320 5640
rect 3680 5630 3720 5640
rect 3760 5630 3800 5640
rect 5120 5630 5160 5640
rect 5240 5630 5280 5640
rect 6920 5630 6960 5640
rect 7720 5630 7800 5640
rect 7920 5630 8000 5640
rect 8320 5630 8400 5640
rect 800 5620 840 5630
rect 1840 5620 1880 5630
rect 2200 5620 2240 5630
rect 2520 5620 2640 5630
rect 3280 5620 3320 5630
rect 3680 5620 3720 5630
rect 3760 5620 3800 5630
rect 5120 5620 5160 5630
rect 5240 5620 5280 5630
rect 6920 5620 6960 5630
rect 7720 5620 7800 5630
rect 7920 5620 8000 5630
rect 8320 5620 8400 5630
rect 720 5610 760 5620
rect 1840 5610 1920 5620
rect 2200 5610 2240 5620
rect 2480 5610 2640 5620
rect 3280 5610 3320 5620
rect 3400 5610 3480 5620
rect 3640 5610 3680 5620
rect 5240 5610 5280 5620
rect 5600 5610 5800 5620
rect 6880 5610 6960 5620
rect 7680 5610 7720 5620
rect 7960 5610 8000 5620
rect 8920 5610 8960 5620
rect 720 5600 760 5610
rect 1840 5600 1920 5610
rect 2200 5600 2240 5610
rect 2480 5600 2640 5610
rect 3280 5600 3320 5610
rect 3400 5600 3480 5610
rect 3640 5600 3680 5610
rect 5240 5600 5280 5610
rect 5600 5600 5800 5610
rect 6880 5600 6960 5610
rect 7680 5600 7720 5610
rect 7960 5600 8000 5610
rect 8920 5600 8960 5610
rect 720 5590 760 5600
rect 1840 5590 1920 5600
rect 2200 5590 2240 5600
rect 2480 5590 2640 5600
rect 3280 5590 3320 5600
rect 3400 5590 3480 5600
rect 3640 5590 3680 5600
rect 5240 5590 5280 5600
rect 5600 5590 5800 5600
rect 6880 5590 6960 5600
rect 7680 5590 7720 5600
rect 7960 5590 8000 5600
rect 8920 5590 8960 5600
rect 720 5580 760 5590
rect 1840 5580 1920 5590
rect 2200 5580 2240 5590
rect 2480 5580 2640 5590
rect 3280 5580 3320 5590
rect 3400 5580 3480 5590
rect 3640 5580 3680 5590
rect 5240 5580 5280 5590
rect 5600 5580 5800 5590
rect 6880 5580 6960 5590
rect 7680 5580 7720 5590
rect 7960 5580 8000 5590
rect 8920 5580 8960 5590
rect 1880 5570 1920 5580
rect 2200 5570 2240 5580
rect 2440 5570 2600 5580
rect 3280 5570 3320 5580
rect 3480 5570 3520 5580
rect 5640 5570 5720 5580
rect 5840 5570 5880 5580
rect 6280 5570 6440 5580
rect 6920 5570 6960 5580
rect 7400 5570 7600 5580
rect 7960 5570 8000 5580
rect 8360 5570 8400 5580
rect 1880 5560 1920 5570
rect 2200 5560 2240 5570
rect 2440 5560 2600 5570
rect 3280 5560 3320 5570
rect 3480 5560 3520 5570
rect 5640 5560 5720 5570
rect 5840 5560 5880 5570
rect 6280 5560 6440 5570
rect 6920 5560 6960 5570
rect 7400 5560 7600 5570
rect 7960 5560 8000 5570
rect 8360 5560 8400 5570
rect 1880 5550 1920 5560
rect 2200 5550 2240 5560
rect 2440 5550 2600 5560
rect 3280 5550 3320 5560
rect 3480 5550 3520 5560
rect 5640 5550 5720 5560
rect 5840 5550 5880 5560
rect 6280 5550 6440 5560
rect 6920 5550 6960 5560
rect 7400 5550 7600 5560
rect 7960 5550 8000 5560
rect 8360 5550 8400 5560
rect 1880 5540 1920 5550
rect 2200 5540 2240 5550
rect 2440 5540 2600 5550
rect 3280 5540 3320 5550
rect 3480 5540 3520 5550
rect 5640 5540 5720 5550
rect 5840 5540 5880 5550
rect 6280 5540 6440 5550
rect 6920 5540 6960 5550
rect 7400 5540 7600 5550
rect 7960 5540 8000 5550
rect 8360 5540 8400 5550
rect 640 5530 680 5540
rect 1880 5530 1960 5540
rect 2200 5530 2240 5540
rect 2400 5530 2600 5540
rect 3240 5530 3320 5540
rect 3480 5530 3520 5540
rect 5120 5530 5160 5540
rect 5720 5530 5920 5540
rect 6240 5530 6280 5540
rect 6440 5530 6520 5540
rect 7400 5530 7480 5540
rect 7760 5530 7800 5540
rect 7960 5530 8040 5540
rect 8120 5530 8200 5540
rect 8720 5530 8760 5540
rect 9000 5530 9040 5540
rect 640 5520 680 5530
rect 1880 5520 1960 5530
rect 2200 5520 2240 5530
rect 2400 5520 2600 5530
rect 3240 5520 3320 5530
rect 3480 5520 3520 5530
rect 5120 5520 5160 5530
rect 5720 5520 5920 5530
rect 6240 5520 6280 5530
rect 6440 5520 6520 5530
rect 7400 5520 7480 5530
rect 7760 5520 7800 5530
rect 7960 5520 8040 5530
rect 8120 5520 8200 5530
rect 8720 5520 8760 5530
rect 9000 5520 9040 5530
rect 640 5510 680 5520
rect 1880 5510 1960 5520
rect 2200 5510 2240 5520
rect 2400 5510 2600 5520
rect 3240 5510 3320 5520
rect 3480 5510 3520 5520
rect 5120 5510 5160 5520
rect 5720 5510 5920 5520
rect 6240 5510 6280 5520
rect 6440 5510 6520 5520
rect 7400 5510 7480 5520
rect 7760 5510 7800 5520
rect 7960 5510 8040 5520
rect 8120 5510 8200 5520
rect 8720 5510 8760 5520
rect 9000 5510 9040 5520
rect 640 5500 680 5510
rect 1880 5500 1960 5510
rect 2200 5500 2240 5510
rect 2400 5500 2600 5510
rect 3240 5500 3320 5510
rect 3480 5500 3520 5510
rect 5120 5500 5160 5510
rect 5720 5500 5920 5510
rect 6240 5500 6280 5510
rect 6440 5500 6520 5510
rect 7400 5500 7480 5510
rect 7760 5500 7800 5510
rect 7960 5500 8040 5510
rect 8120 5500 8200 5510
rect 8720 5500 8760 5510
rect 9000 5500 9040 5510
rect 440 5490 640 5500
rect 920 5490 1000 5500
rect 1880 5490 1960 5500
rect 2200 5490 2240 5500
rect 2400 5490 2560 5500
rect 3240 5490 3320 5500
rect 3560 5490 3600 5500
rect 5120 5490 5160 5500
rect 5720 5490 5920 5500
rect 6200 5490 6240 5500
rect 6360 5490 6440 5500
rect 7400 5490 7480 5500
rect 7760 5490 7800 5500
rect 7960 5490 8160 5500
rect 8520 5490 8600 5500
rect 9120 5490 9160 5500
rect 440 5480 640 5490
rect 920 5480 1000 5490
rect 1880 5480 1960 5490
rect 2200 5480 2240 5490
rect 2400 5480 2560 5490
rect 3240 5480 3320 5490
rect 3560 5480 3600 5490
rect 5120 5480 5160 5490
rect 5720 5480 5920 5490
rect 6200 5480 6240 5490
rect 6360 5480 6440 5490
rect 7400 5480 7480 5490
rect 7760 5480 7800 5490
rect 7960 5480 8160 5490
rect 8520 5480 8600 5490
rect 9120 5480 9160 5490
rect 440 5470 640 5480
rect 920 5470 1000 5480
rect 1880 5470 1960 5480
rect 2200 5470 2240 5480
rect 2400 5470 2560 5480
rect 3240 5470 3320 5480
rect 3560 5470 3600 5480
rect 5120 5470 5160 5480
rect 5720 5470 5920 5480
rect 6200 5470 6240 5480
rect 6360 5470 6440 5480
rect 7400 5470 7480 5480
rect 7760 5470 7800 5480
rect 7960 5470 8160 5480
rect 8520 5470 8600 5480
rect 9120 5470 9160 5480
rect 440 5460 640 5470
rect 920 5460 1000 5470
rect 1880 5460 1960 5470
rect 2200 5460 2240 5470
rect 2400 5460 2560 5470
rect 3240 5460 3320 5470
rect 3560 5460 3600 5470
rect 5120 5460 5160 5470
rect 5720 5460 5920 5470
rect 6200 5460 6240 5470
rect 6360 5460 6440 5470
rect 7400 5460 7480 5470
rect 7760 5460 7800 5470
rect 7960 5460 8160 5470
rect 8520 5460 8600 5470
rect 9120 5460 9160 5470
rect 480 5450 520 5460
rect 1920 5450 1960 5460
rect 2400 5450 2440 5460
rect 2560 5450 2600 5460
rect 2880 5450 2920 5460
rect 3240 5450 3320 5460
rect 5120 5450 5160 5460
rect 5480 5450 5600 5460
rect 5640 5450 5720 5460
rect 5800 5450 5920 5460
rect 6200 5450 6240 5460
rect 6360 5450 6480 5460
rect 7400 5450 7520 5460
rect 7960 5450 8160 5460
rect 8480 5450 8520 5460
rect 9520 5450 9560 5460
rect 480 5440 520 5450
rect 1920 5440 1960 5450
rect 2400 5440 2440 5450
rect 2560 5440 2600 5450
rect 2880 5440 2920 5450
rect 3240 5440 3320 5450
rect 5120 5440 5160 5450
rect 5480 5440 5600 5450
rect 5640 5440 5720 5450
rect 5800 5440 5920 5450
rect 6200 5440 6240 5450
rect 6360 5440 6480 5450
rect 7400 5440 7520 5450
rect 7960 5440 8160 5450
rect 8480 5440 8520 5450
rect 9520 5440 9560 5450
rect 480 5430 520 5440
rect 1920 5430 1960 5440
rect 2400 5430 2440 5440
rect 2560 5430 2600 5440
rect 2880 5430 2920 5440
rect 3240 5430 3320 5440
rect 5120 5430 5160 5440
rect 5480 5430 5600 5440
rect 5640 5430 5720 5440
rect 5800 5430 5920 5440
rect 6200 5430 6240 5440
rect 6360 5430 6480 5440
rect 7400 5430 7520 5440
rect 7960 5430 8160 5440
rect 8480 5430 8520 5440
rect 9520 5430 9560 5440
rect 480 5420 520 5430
rect 1920 5420 1960 5430
rect 2400 5420 2440 5430
rect 2560 5420 2600 5430
rect 2880 5420 2920 5430
rect 3240 5420 3320 5430
rect 5120 5420 5160 5430
rect 5480 5420 5600 5430
rect 5640 5420 5720 5430
rect 5800 5420 5920 5430
rect 6200 5420 6240 5430
rect 6360 5420 6480 5430
rect 7400 5420 7520 5430
rect 7960 5420 8160 5430
rect 8480 5420 8520 5430
rect 9520 5420 9560 5430
rect 440 5410 480 5420
rect 560 5410 600 5420
rect 1920 5410 1960 5420
rect 2400 5410 2440 5420
rect 2560 5410 2680 5420
rect 2880 5410 3080 5420
rect 3160 5410 3240 5420
rect 5200 5410 5240 5420
rect 5440 5410 5560 5420
rect 5840 5410 5920 5420
rect 6200 5410 6240 5420
rect 6560 5410 6600 5420
rect 7400 5410 7520 5420
rect 7800 5410 7880 5420
rect 7960 5410 8160 5420
rect 8280 5410 8320 5420
rect 8960 5410 9000 5420
rect 9080 5410 9120 5420
rect 440 5400 480 5410
rect 560 5400 600 5410
rect 1920 5400 1960 5410
rect 2400 5400 2440 5410
rect 2560 5400 2680 5410
rect 2880 5400 3080 5410
rect 3160 5400 3240 5410
rect 5200 5400 5240 5410
rect 5440 5400 5560 5410
rect 5840 5400 5920 5410
rect 6200 5400 6240 5410
rect 6560 5400 6600 5410
rect 7400 5400 7520 5410
rect 7800 5400 7880 5410
rect 7960 5400 8160 5410
rect 8280 5400 8320 5410
rect 8960 5400 9000 5410
rect 9080 5400 9120 5410
rect 440 5390 480 5400
rect 560 5390 600 5400
rect 1920 5390 1960 5400
rect 2400 5390 2440 5400
rect 2560 5390 2680 5400
rect 2880 5390 3080 5400
rect 3160 5390 3240 5400
rect 5200 5390 5240 5400
rect 5440 5390 5560 5400
rect 5840 5390 5920 5400
rect 6200 5390 6240 5400
rect 6560 5390 6600 5400
rect 7400 5390 7520 5400
rect 7800 5390 7880 5400
rect 7960 5390 8160 5400
rect 8280 5390 8320 5400
rect 8960 5390 9000 5400
rect 9080 5390 9120 5400
rect 440 5380 480 5390
rect 560 5380 600 5390
rect 1920 5380 1960 5390
rect 2400 5380 2440 5390
rect 2560 5380 2680 5390
rect 2880 5380 3080 5390
rect 3160 5380 3240 5390
rect 5200 5380 5240 5390
rect 5440 5380 5560 5390
rect 5840 5380 5920 5390
rect 6200 5380 6240 5390
rect 6560 5380 6600 5390
rect 7400 5380 7520 5390
rect 7800 5380 7880 5390
rect 7960 5380 8160 5390
rect 8280 5380 8320 5390
rect 8960 5380 9000 5390
rect 9080 5380 9120 5390
rect 360 5370 400 5380
rect 1920 5370 2000 5380
rect 2400 5370 2440 5380
rect 2480 5370 2520 5380
rect 2560 5370 2600 5380
rect 2720 5370 3040 5380
rect 3480 5370 3520 5380
rect 5600 5370 5760 5380
rect 5840 5370 5880 5380
rect 6360 5370 6400 5380
rect 6640 5370 6680 5380
rect 7400 5370 7520 5380
rect 7640 5370 7800 5380
rect 7840 5370 7880 5380
rect 7960 5370 8120 5380
rect 8160 5370 8200 5380
rect 8840 5370 8880 5380
rect 9240 5370 9280 5380
rect 9360 5370 9400 5380
rect 360 5360 400 5370
rect 1920 5360 2000 5370
rect 2400 5360 2440 5370
rect 2480 5360 2520 5370
rect 2560 5360 2600 5370
rect 2720 5360 3040 5370
rect 3480 5360 3520 5370
rect 5600 5360 5760 5370
rect 5840 5360 5880 5370
rect 6360 5360 6400 5370
rect 6640 5360 6680 5370
rect 7400 5360 7520 5370
rect 7640 5360 7800 5370
rect 7840 5360 7880 5370
rect 7960 5360 8120 5370
rect 8160 5360 8200 5370
rect 8840 5360 8880 5370
rect 9240 5360 9280 5370
rect 9360 5360 9400 5370
rect 360 5350 400 5360
rect 1920 5350 2000 5360
rect 2400 5350 2440 5360
rect 2480 5350 2520 5360
rect 2560 5350 2600 5360
rect 2720 5350 3040 5360
rect 3480 5350 3520 5360
rect 5600 5350 5760 5360
rect 5840 5350 5880 5360
rect 6360 5350 6400 5360
rect 6640 5350 6680 5360
rect 7400 5350 7520 5360
rect 7640 5350 7800 5360
rect 7840 5350 7880 5360
rect 7960 5350 8120 5360
rect 8160 5350 8200 5360
rect 8840 5350 8880 5360
rect 9240 5350 9280 5360
rect 9360 5350 9400 5360
rect 360 5340 400 5350
rect 1920 5340 2000 5350
rect 2400 5340 2440 5350
rect 2480 5340 2520 5350
rect 2560 5340 2600 5350
rect 2720 5340 3040 5350
rect 3480 5340 3520 5350
rect 5600 5340 5760 5350
rect 5840 5340 5880 5350
rect 6360 5340 6400 5350
rect 6640 5340 6680 5350
rect 7400 5340 7520 5350
rect 7640 5340 7800 5350
rect 7840 5340 7880 5350
rect 7960 5340 8120 5350
rect 8160 5340 8200 5350
rect 8840 5340 8880 5350
rect 9240 5340 9280 5350
rect 9360 5340 9400 5350
rect 560 5330 600 5340
rect 1920 5330 2000 5340
rect 2400 5330 2480 5340
rect 2520 5330 2600 5340
rect 2720 5330 3040 5340
rect 5160 5330 5200 5340
rect 5760 5330 5800 5340
rect 6200 5330 6560 5340
rect 6640 5330 6720 5340
rect 7360 5330 7720 5340
rect 7840 5330 7880 5340
rect 8320 5330 8360 5340
rect 8480 5330 8520 5340
rect 8760 5330 8800 5340
rect 9360 5330 9400 5340
rect 9600 5330 9640 5340
rect 560 5320 600 5330
rect 1920 5320 2000 5330
rect 2400 5320 2480 5330
rect 2520 5320 2600 5330
rect 2720 5320 3040 5330
rect 5160 5320 5200 5330
rect 5760 5320 5800 5330
rect 6200 5320 6560 5330
rect 6640 5320 6720 5330
rect 7360 5320 7720 5330
rect 7840 5320 7880 5330
rect 8320 5320 8360 5330
rect 8480 5320 8520 5330
rect 8760 5320 8800 5330
rect 9360 5320 9400 5330
rect 9600 5320 9640 5330
rect 560 5310 600 5320
rect 1920 5310 2000 5320
rect 2400 5310 2480 5320
rect 2520 5310 2600 5320
rect 2720 5310 3040 5320
rect 5160 5310 5200 5320
rect 5760 5310 5800 5320
rect 6200 5310 6560 5320
rect 6640 5310 6720 5320
rect 7360 5310 7720 5320
rect 7840 5310 7880 5320
rect 8320 5310 8360 5320
rect 8480 5310 8520 5320
rect 8760 5310 8800 5320
rect 9360 5310 9400 5320
rect 9600 5310 9640 5320
rect 560 5300 600 5310
rect 1920 5300 2000 5310
rect 2400 5300 2480 5310
rect 2520 5300 2600 5310
rect 2720 5300 3040 5310
rect 5160 5300 5200 5310
rect 5760 5300 5800 5310
rect 6200 5300 6560 5310
rect 6640 5300 6720 5310
rect 7360 5300 7720 5310
rect 7840 5300 7880 5310
rect 8320 5300 8360 5310
rect 8480 5300 8520 5310
rect 8760 5300 8800 5310
rect 9360 5300 9400 5310
rect 9600 5300 9640 5310
rect 600 5290 640 5300
rect 1920 5290 2000 5300
rect 2400 5290 2440 5300
rect 2600 5290 2640 5300
rect 2800 5290 3000 5300
rect 6320 5290 6360 5300
rect 7320 5290 7640 5300
rect 7840 5290 7920 5300
rect 8600 5290 8680 5300
rect 8920 5290 8960 5300
rect 9080 5290 9120 5300
rect 9400 5290 9440 5300
rect 9880 5290 9920 5300
rect 600 5280 640 5290
rect 1920 5280 2000 5290
rect 2400 5280 2440 5290
rect 2600 5280 2640 5290
rect 2800 5280 3000 5290
rect 6320 5280 6360 5290
rect 7320 5280 7640 5290
rect 7840 5280 7920 5290
rect 8600 5280 8680 5290
rect 8920 5280 8960 5290
rect 9080 5280 9120 5290
rect 9400 5280 9440 5290
rect 9880 5280 9920 5290
rect 600 5270 640 5280
rect 1920 5270 2000 5280
rect 2400 5270 2440 5280
rect 2600 5270 2640 5280
rect 2800 5270 3000 5280
rect 6320 5270 6360 5280
rect 7320 5270 7640 5280
rect 7840 5270 7920 5280
rect 8600 5270 8680 5280
rect 8920 5270 8960 5280
rect 9080 5270 9120 5280
rect 9400 5270 9440 5280
rect 9880 5270 9920 5280
rect 600 5260 640 5270
rect 1920 5260 2000 5270
rect 2400 5260 2440 5270
rect 2600 5260 2640 5270
rect 2800 5260 3000 5270
rect 6320 5260 6360 5270
rect 7320 5260 7640 5270
rect 7840 5260 7920 5270
rect 8600 5260 8680 5270
rect 8920 5260 8960 5270
rect 9080 5260 9120 5270
rect 9400 5260 9440 5270
rect 9880 5260 9920 5270
rect 1960 5250 2040 5260
rect 2880 5250 2960 5260
rect 7360 5250 7480 5260
rect 7560 5250 7680 5260
rect 7840 5250 7920 5260
rect 8440 5250 8480 5260
rect 8800 5250 8840 5260
rect 8880 5250 8920 5260
rect 1960 5240 2040 5250
rect 2880 5240 2960 5250
rect 7360 5240 7480 5250
rect 7560 5240 7680 5250
rect 7840 5240 7920 5250
rect 8440 5240 8480 5250
rect 8800 5240 8840 5250
rect 8880 5240 8920 5250
rect 1960 5230 2040 5240
rect 2880 5230 2960 5240
rect 7360 5230 7480 5240
rect 7560 5230 7680 5240
rect 7840 5230 7920 5240
rect 8440 5230 8480 5240
rect 8800 5230 8840 5240
rect 8880 5230 8920 5240
rect 1960 5220 2040 5230
rect 2880 5220 2960 5230
rect 7360 5220 7480 5230
rect 7560 5220 7680 5230
rect 7840 5220 7920 5230
rect 8440 5220 8480 5230
rect 8800 5220 8840 5230
rect 8880 5220 8920 5230
rect 680 5210 720 5220
rect 1960 5210 2040 5220
rect 2680 5210 2720 5220
rect 2920 5210 3000 5220
rect 5080 5210 5160 5220
rect 7360 5210 7440 5220
rect 7520 5210 7680 5220
rect 7840 5210 7960 5220
rect 8280 5210 8320 5220
rect 8640 5210 8680 5220
rect 8800 5210 8840 5220
rect 8880 5210 8920 5220
rect 9360 5210 9400 5220
rect 9760 5210 9800 5220
rect 680 5200 720 5210
rect 1960 5200 2040 5210
rect 2680 5200 2720 5210
rect 2920 5200 3000 5210
rect 5080 5200 5160 5210
rect 7360 5200 7440 5210
rect 7520 5200 7680 5210
rect 7840 5200 7960 5210
rect 8280 5200 8320 5210
rect 8640 5200 8680 5210
rect 8800 5200 8840 5210
rect 8880 5200 8920 5210
rect 9360 5200 9400 5210
rect 9760 5200 9800 5210
rect 680 5190 720 5200
rect 1960 5190 2040 5200
rect 2680 5190 2720 5200
rect 2920 5190 3000 5200
rect 5080 5190 5160 5200
rect 7360 5190 7440 5200
rect 7520 5190 7680 5200
rect 7840 5190 7960 5200
rect 8280 5190 8320 5200
rect 8640 5190 8680 5200
rect 8800 5190 8840 5200
rect 8880 5190 8920 5200
rect 9360 5190 9400 5200
rect 9760 5190 9800 5200
rect 680 5180 720 5190
rect 1960 5180 2040 5190
rect 2680 5180 2720 5190
rect 2920 5180 3000 5190
rect 5080 5180 5160 5190
rect 7360 5180 7440 5190
rect 7520 5180 7680 5190
rect 7840 5180 7960 5190
rect 8280 5180 8320 5190
rect 8640 5180 8680 5190
rect 8800 5180 8840 5190
rect 8880 5180 8920 5190
rect 9360 5180 9400 5190
rect 9760 5180 9800 5190
rect 680 5170 720 5180
rect 1800 5170 1880 5180
rect 1960 5170 2040 5180
rect 2720 5170 2800 5180
rect 3000 5170 3040 5180
rect 5120 5170 5160 5180
rect 7360 5170 7440 5180
rect 7560 5170 7600 5180
rect 7880 5170 7960 5180
rect 8000 5170 8040 5180
rect 8200 5170 8280 5180
rect 8720 5170 8760 5180
rect 8880 5170 8920 5180
rect 9360 5170 9400 5180
rect 9680 5170 9720 5180
rect 9840 5170 9880 5180
rect 680 5160 720 5170
rect 1800 5160 1880 5170
rect 1960 5160 2040 5170
rect 2720 5160 2800 5170
rect 3000 5160 3040 5170
rect 5120 5160 5160 5170
rect 7360 5160 7440 5170
rect 7560 5160 7600 5170
rect 7880 5160 7960 5170
rect 8000 5160 8040 5170
rect 8200 5160 8280 5170
rect 8720 5160 8760 5170
rect 8880 5160 8920 5170
rect 9360 5160 9400 5170
rect 9680 5160 9720 5170
rect 9840 5160 9880 5170
rect 680 5150 720 5160
rect 1800 5150 1880 5160
rect 1960 5150 2040 5160
rect 2720 5150 2800 5160
rect 3000 5150 3040 5160
rect 5120 5150 5160 5160
rect 7360 5150 7440 5160
rect 7560 5150 7600 5160
rect 7880 5150 7960 5160
rect 8000 5150 8040 5160
rect 8200 5150 8280 5160
rect 8720 5150 8760 5160
rect 8880 5150 8920 5160
rect 9360 5150 9400 5160
rect 9680 5150 9720 5160
rect 9840 5150 9880 5160
rect 680 5140 720 5150
rect 1800 5140 1880 5150
rect 1960 5140 2040 5150
rect 2720 5140 2800 5150
rect 3000 5140 3040 5150
rect 5120 5140 5160 5150
rect 7360 5140 7440 5150
rect 7560 5140 7600 5150
rect 7880 5140 7960 5150
rect 8000 5140 8040 5150
rect 8200 5140 8280 5150
rect 8720 5140 8760 5150
rect 8880 5140 8920 5150
rect 9360 5140 9400 5150
rect 9680 5140 9720 5150
rect 9840 5140 9880 5150
rect 600 5130 760 5140
rect 1800 5130 1880 5140
rect 1960 5130 2080 5140
rect 2800 5130 2920 5140
rect 2960 5130 3040 5140
rect 3400 5130 3440 5140
rect 7320 5130 7440 5140
rect 7880 5130 7960 5140
rect 8000 5130 8040 5140
rect 8080 5130 8240 5140
rect 8800 5130 8840 5140
rect 9440 5130 9520 5140
rect 9560 5130 9600 5140
rect 600 5120 760 5130
rect 1800 5120 1880 5130
rect 1960 5120 2080 5130
rect 2800 5120 2920 5130
rect 2960 5120 3040 5130
rect 3400 5120 3440 5130
rect 7320 5120 7440 5130
rect 7880 5120 7960 5130
rect 8000 5120 8040 5130
rect 8080 5120 8240 5130
rect 8800 5120 8840 5130
rect 9440 5120 9520 5130
rect 9560 5120 9600 5130
rect 600 5110 760 5120
rect 1800 5110 1880 5120
rect 1960 5110 2080 5120
rect 2800 5110 2920 5120
rect 2960 5110 3040 5120
rect 3400 5110 3440 5120
rect 7320 5110 7440 5120
rect 7880 5110 7960 5120
rect 8000 5110 8040 5120
rect 8080 5110 8240 5120
rect 8800 5110 8840 5120
rect 9440 5110 9520 5120
rect 9560 5110 9600 5120
rect 600 5100 760 5110
rect 1800 5100 1880 5110
rect 1960 5100 2080 5110
rect 2800 5100 2920 5110
rect 2960 5100 3040 5110
rect 3400 5100 3440 5110
rect 7320 5100 7440 5110
rect 7880 5100 7960 5110
rect 8000 5100 8040 5110
rect 8080 5100 8240 5110
rect 8800 5100 8840 5110
rect 9440 5100 9520 5110
rect 9560 5100 9600 5110
rect 600 5090 640 5100
rect 680 5090 760 5100
rect 1760 5090 1880 5100
rect 1960 5090 2080 5100
rect 2840 5090 2960 5100
rect 5160 5090 5200 5100
rect 7320 5090 7440 5100
rect 7880 5090 8000 5100
rect 8120 5090 8280 5100
rect 8640 5090 8680 5100
rect 8840 5090 8920 5100
rect 9200 5090 9240 5100
rect 9560 5090 9600 5100
rect 9720 5090 9760 5100
rect 600 5080 640 5090
rect 680 5080 760 5090
rect 1760 5080 1880 5090
rect 1960 5080 2080 5090
rect 2840 5080 2960 5090
rect 5160 5080 5200 5090
rect 7320 5080 7440 5090
rect 7880 5080 8000 5090
rect 8120 5080 8280 5090
rect 8640 5080 8680 5090
rect 8840 5080 8920 5090
rect 9200 5080 9240 5090
rect 9560 5080 9600 5090
rect 9720 5080 9760 5090
rect 600 5070 640 5080
rect 680 5070 760 5080
rect 1760 5070 1880 5080
rect 1960 5070 2080 5080
rect 2840 5070 2960 5080
rect 5160 5070 5200 5080
rect 7320 5070 7440 5080
rect 7880 5070 8000 5080
rect 8120 5070 8280 5080
rect 8640 5070 8680 5080
rect 8840 5070 8920 5080
rect 9200 5070 9240 5080
rect 9560 5070 9600 5080
rect 9720 5070 9760 5080
rect 600 5060 640 5070
rect 680 5060 760 5070
rect 1760 5060 1880 5070
rect 1960 5060 2080 5070
rect 2840 5060 2960 5070
rect 5160 5060 5200 5070
rect 7320 5060 7440 5070
rect 7880 5060 8000 5070
rect 8120 5060 8280 5070
rect 8640 5060 8680 5070
rect 8840 5060 8920 5070
rect 9200 5060 9240 5070
rect 9560 5060 9600 5070
rect 9720 5060 9760 5070
rect 400 5050 640 5060
rect 1760 5050 1880 5060
rect 2000 5050 2080 5060
rect 2880 5050 3040 5060
rect 3360 5050 3400 5060
rect 7320 5050 7480 5060
rect 7880 5050 8000 5060
rect 8040 5050 8160 5060
rect 8400 5050 8440 5060
rect 9000 5050 9040 5060
rect 9360 5050 9400 5060
rect 400 5040 640 5050
rect 1760 5040 1880 5050
rect 2000 5040 2080 5050
rect 2880 5040 3040 5050
rect 3360 5040 3400 5050
rect 7320 5040 7480 5050
rect 7880 5040 8000 5050
rect 8040 5040 8160 5050
rect 8400 5040 8440 5050
rect 9000 5040 9040 5050
rect 9360 5040 9400 5050
rect 400 5030 640 5040
rect 1760 5030 1880 5040
rect 2000 5030 2080 5040
rect 2880 5030 3040 5040
rect 3360 5030 3400 5040
rect 7320 5030 7480 5040
rect 7880 5030 8000 5040
rect 8040 5030 8160 5040
rect 8400 5030 8440 5040
rect 9000 5030 9040 5040
rect 9360 5030 9400 5040
rect 400 5020 640 5030
rect 1760 5020 1880 5030
rect 2000 5020 2080 5030
rect 2880 5020 3040 5030
rect 3360 5020 3400 5030
rect 7320 5020 7480 5030
rect 7880 5020 8000 5030
rect 8040 5020 8160 5030
rect 8400 5020 8440 5030
rect 9000 5020 9040 5030
rect 9360 5020 9400 5030
rect 400 5010 480 5020
rect 1760 5010 1840 5020
rect 2000 5010 2120 5020
rect 2760 5010 3040 5020
rect 3320 5010 3360 5020
rect 7320 5010 7360 5020
rect 7880 5010 8000 5020
rect 8400 5010 8440 5020
rect 400 5000 480 5010
rect 1760 5000 1840 5010
rect 2000 5000 2120 5010
rect 2760 5000 3040 5010
rect 3320 5000 3360 5010
rect 7320 5000 7360 5010
rect 7880 5000 8000 5010
rect 8400 5000 8440 5010
rect 400 4990 480 5000
rect 1760 4990 1840 5000
rect 2000 4990 2120 5000
rect 2760 4990 3040 5000
rect 3320 4990 3360 5000
rect 7320 4990 7360 5000
rect 7880 4990 8000 5000
rect 8400 4990 8440 5000
rect 400 4980 480 4990
rect 1760 4980 1840 4990
rect 2000 4980 2120 4990
rect 2760 4980 3040 4990
rect 3320 4980 3360 4990
rect 7320 4980 7360 4990
rect 7880 4980 8000 4990
rect 8400 4980 8440 4990
rect 400 4970 560 4980
rect 2080 4970 2160 4980
rect 2680 4970 2720 4980
rect 2760 4970 2960 4980
rect 3320 4970 3360 4980
rect 4000 4970 4040 4980
rect 4200 4970 4280 4980
rect 4320 4970 4360 4980
rect 7320 4970 7360 4980
rect 7800 4970 7840 4980
rect 7960 4970 8000 4980
rect 8440 4970 8480 4980
rect 8600 4970 8640 4980
rect 9120 4970 9160 4980
rect 9240 4970 9360 4980
rect 9520 4970 9600 4980
rect 400 4960 560 4970
rect 2080 4960 2160 4970
rect 2680 4960 2720 4970
rect 2760 4960 2960 4970
rect 3320 4960 3360 4970
rect 4000 4960 4040 4970
rect 4200 4960 4280 4970
rect 4320 4960 4360 4970
rect 7320 4960 7360 4970
rect 7800 4960 7840 4970
rect 7960 4960 8000 4970
rect 8440 4960 8480 4970
rect 8600 4960 8640 4970
rect 9120 4960 9160 4970
rect 9240 4960 9360 4970
rect 9520 4960 9600 4970
rect 400 4950 560 4960
rect 2080 4950 2160 4960
rect 2680 4950 2720 4960
rect 2760 4950 2960 4960
rect 3320 4950 3360 4960
rect 4000 4950 4040 4960
rect 4200 4950 4280 4960
rect 4320 4950 4360 4960
rect 7320 4950 7360 4960
rect 7800 4950 7840 4960
rect 7960 4950 8000 4960
rect 8440 4950 8480 4960
rect 8600 4950 8640 4960
rect 9120 4950 9160 4960
rect 9240 4950 9360 4960
rect 9520 4950 9600 4960
rect 400 4940 560 4950
rect 2080 4940 2160 4950
rect 2680 4940 2720 4950
rect 2760 4940 2960 4950
rect 3320 4940 3360 4950
rect 4000 4940 4040 4950
rect 4200 4940 4280 4950
rect 4320 4940 4360 4950
rect 7320 4940 7360 4950
rect 7800 4940 7840 4950
rect 7960 4940 8000 4950
rect 8440 4940 8480 4950
rect 8600 4940 8640 4950
rect 9120 4940 9160 4950
rect 9240 4940 9360 4950
rect 9520 4940 9600 4950
rect 240 4930 320 4940
rect 400 4930 720 4940
rect 1040 4930 1080 4940
rect 2160 4930 2200 4940
rect 2240 4930 2320 4940
rect 2640 4930 2880 4940
rect 3280 4930 3320 4940
rect 4000 4930 4040 4940
rect 4360 4930 4400 4940
rect 5640 4930 5720 4940
rect 5840 4930 5920 4940
rect 6320 4930 6400 4940
rect 7720 4930 7760 4940
rect 7960 4930 8000 4940
rect 8560 4930 8600 4940
rect 9480 4930 9520 4940
rect 240 4920 320 4930
rect 400 4920 720 4930
rect 1040 4920 1080 4930
rect 2160 4920 2200 4930
rect 2240 4920 2320 4930
rect 2640 4920 2880 4930
rect 3280 4920 3320 4930
rect 4000 4920 4040 4930
rect 4360 4920 4400 4930
rect 5640 4920 5720 4930
rect 5840 4920 5920 4930
rect 6320 4920 6400 4930
rect 7720 4920 7760 4930
rect 7960 4920 8000 4930
rect 8560 4920 8600 4930
rect 9480 4920 9520 4930
rect 240 4910 320 4920
rect 400 4910 720 4920
rect 1040 4910 1080 4920
rect 2160 4910 2200 4920
rect 2240 4910 2320 4920
rect 2640 4910 2880 4920
rect 3280 4910 3320 4920
rect 4000 4910 4040 4920
rect 4360 4910 4400 4920
rect 5640 4910 5720 4920
rect 5840 4910 5920 4920
rect 6320 4910 6400 4920
rect 7720 4910 7760 4920
rect 7960 4910 8000 4920
rect 8560 4910 8600 4920
rect 9480 4910 9520 4920
rect 240 4900 320 4910
rect 400 4900 720 4910
rect 1040 4900 1080 4910
rect 2160 4900 2200 4910
rect 2240 4900 2320 4910
rect 2640 4900 2880 4910
rect 3280 4900 3320 4910
rect 4000 4900 4040 4910
rect 4360 4900 4400 4910
rect 5640 4900 5720 4910
rect 5840 4900 5920 4910
rect 6320 4900 6400 4910
rect 7720 4900 7760 4910
rect 7960 4900 8000 4910
rect 8560 4900 8600 4910
rect 9480 4900 9520 4910
rect 80 4890 760 4900
rect 1040 4890 1080 4900
rect 2200 4890 2360 4900
rect 2680 4890 2800 4900
rect 3160 4890 3200 4900
rect 3280 4890 3320 4900
rect 4160 4890 4200 4900
rect 4480 4890 4680 4900
rect 4720 4890 4760 4900
rect 5600 4890 5680 4900
rect 5840 4890 5960 4900
rect 6040 4890 6080 4900
rect 6120 4890 6200 4900
rect 6280 4890 6440 4900
rect 7360 4890 7400 4900
rect 7960 4890 8000 4900
rect 8320 4890 8360 4900
rect 8720 4890 8760 4900
rect 8880 4890 8920 4900
rect 80 4880 760 4890
rect 1040 4880 1080 4890
rect 2200 4880 2360 4890
rect 2680 4880 2800 4890
rect 3160 4880 3200 4890
rect 3280 4880 3320 4890
rect 4160 4880 4200 4890
rect 4480 4880 4680 4890
rect 4720 4880 4760 4890
rect 5600 4880 5680 4890
rect 5840 4880 5960 4890
rect 6040 4880 6080 4890
rect 6120 4880 6200 4890
rect 6280 4880 6440 4890
rect 7360 4880 7400 4890
rect 7960 4880 8000 4890
rect 8320 4880 8360 4890
rect 8720 4880 8760 4890
rect 8880 4880 8920 4890
rect 80 4870 760 4880
rect 1040 4870 1080 4880
rect 2200 4870 2360 4880
rect 2680 4870 2800 4880
rect 3160 4870 3200 4880
rect 3280 4870 3320 4880
rect 4160 4870 4200 4880
rect 4480 4870 4680 4880
rect 4720 4870 4760 4880
rect 5600 4870 5680 4880
rect 5840 4870 5960 4880
rect 6040 4870 6080 4880
rect 6120 4870 6200 4880
rect 6280 4870 6440 4880
rect 7360 4870 7400 4880
rect 7960 4870 8000 4880
rect 8320 4870 8360 4880
rect 8720 4870 8760 4880
rect 8880 4870 8920 4880
rect 80 4860 760 4870
rect 1040 4860 1080 4870
rect 2200 4860 2360 4870
rect 2680 4860 2800 4870
rect 3160 4860 3200 4870
rect 3280 4860 3320 4870
rect 4160 4860 4200 4870
rect 4480 4860 4680 4870
rect 4720 4860 4760 4870
rect 5600 4860 5680 4870
rect 5840 4860 5960 4870
rect 6040 4860 6080 4870
rect 6120 4860 6200 4870
rect 6280 4860 6440 4870
rect 7360 4860 7400 4870
rect 7960 4860 8000 4870
rect 8320 4860 8360 4870
rect 8720 4860 8760 4870
rect 8880 4860 8920 4870
rect 160 4850 800 4860
rect 1040 4850 1120 4860
rect 2320 4850 2360 4860
rect 2680 4850 2800 4860
rect 3080 4850 3160 4860
rect 3240 4850 3280 4860
rect 3320 4850 3360 4860
rect 3680 4850 3720 4860
rect 3840 4850 3880 4860
rect 3920 4850 3960 4860
rect 4880 4850 4920 4860
rect 5560 4850 5680 4860
rect 6000 4850 6480 4860
rect 7360 4850 7400 4860
rect 7960 4850 8080 4860
rect 8440 4850 8480 4860
rect 9360 4850 9400 4860
rect 9600 4850 9640 4860
rect 160 4840 800 4850
rect 1040 4840 1120 4850
rect 2320 4840 2360 4850
rect 2680 4840 2800 4850
rect 3080 4840 3160 4850
rect 3240 4840 3280 4850
rect 3320 4840 3360 4850
rect 3680 4840 3720 4850
rect 3840 4840 3880 4850
rect 3920 4840 3960 4850
rect 4880 4840 4920 4850
rect 5560 4840 5680 4850
rect 6000 4840 6480 4850
rect 7360 4840 7400 4850
rect 7960 4840 8080 4850
rect 8440 4840 8480 4850
rect 9360 4840 9400 4850
rect 9600 4840 9640 4850
rect 160 4830 800 4840
rect 1040 4830 1120 4840
rect 2320 4830 2360 4840
rect 2680 4830 2800 4840
rect 3080 4830 3160 4840
rect 3240 4830 3280 4840
rect 3320 4830 3360 4840
rect 3680 4830 3720 4840
rect 3840 4830 3880 4840
rect 3920 4830 3960 4840
rect 4880 4830 4920 4840
rect 5560 4830 5680 4840
rect 6000 4830 6480 4840
rect 7360 4830 7400 4840
rect 7960 4830 8080 4840
rect 8440 4830 8480 4840
rect 9360 4830 9400 4840
rect 9600 4830 9640 4840
rect 160 4820 800 4830
rect 1040 4820 1120 4830
rect 2320 4820 2360 4830
rect 2680 4820 2800 4830
rect 3080 4820 3160 4830
rect 3240 4820 3280 4830
rect 3320 4820 3360 4830
rect 3680 4820 3720 4830
rect 3840 4820 3880 4830
rect 3920 4820 3960 4830
rect 4880 4820 4920 4830
rect 5560 4820 5680 4830
rect 6000 4820 6480 4830
rect 7360 4820 7400 4830
rect 7960 4820 8080 4830
rect 8440 4820 8480 4830
rect 9360 4820 9400 4830
rect 9600 4820 9640 4830
rect 200 4810 480 4820
rect 560 4810 880 4820
rect 1040 4810 1120 4820
rect 2760 4810 2920 4820
rect 3040 4810 3160 4820
rect 3200 4810 3280 4820
rect 3320 4810 3360 4820
rect 3720 4810 3800 4820
rect 3880 4810 3960 4820
rect 4920 4810 5000 4820
rect 5200 4810 5240 4820
rect 5520 4810 5560 4820
rect 5600 4810 5640 4820
rect 6000 4810 6240 4820
rect 6360 4810 6520 4820
rect 7840 4810 7920 4820
rect 7960 4810 8000 4820
rect 8080 4810 8120 4820
rect 8720 4810 8760 4820
rect 8920 4810 8960 4820
rect 9440 4810 9480 4820
rect 9680 4810 9720 4820
rect 200 4800 480 4810
rect 560 4800 880 4810
rect 1040 4800 1120 4810
rect 2760 4800 2920 4810
rect 3040 4800 3160 4810
rect 3200 4800 3280 4810
rect 3320 4800 3360 4810
rect 3720 4800 3800 4810
rect 3880 4800 3960 4810
rect 4920 4800 5000 4810
rect 5200 4800 5240 4810
rect 5520 4800 5560 4810
rect 5600 4800 5640 4810
rect 6000 4800 6240 4810
rect 6360 4800 6520 4810
rect 7840 4800 7920 4810
rect 7960 4800 8000 4810
rect 8080 4800 8120 4810
rect 8720 4800 8760 4810
rect 8920 4800 8960 4810
rect 9440 4800 9480 4810
rect 9680 4800 9720 4810
rect 200 4790 480 4800
rect 560 4790 880 4800
rect 1040 4790 1120 4800
rect 2760 4790 2920 4800
rect 3040 4790 3160 4800
rect 3200 4790 3280 4800
rect 3320 4790 3360 4800
rect 3720 4790 3800 4800
rect 3880 4790 3960 4800
rect 4920 4790 5000 4800
rect 5200 4790 5240 4800
rect 5520 4790 5560 4800
rect 5600 4790 5640 4800
rect 6000 4790 6240 4800
rect 6360 4790 6520 4800
rect 7840 4790 7920 4800
rect 7960 4790 8000 4800
rect 8080 4790 8120 4800
rect 8720 4790 8760 4800
rect 8920 4790 8960 4800
rect 9440 4790 9480 4800
rect 9680 4790 9720 4800
rect 200 4780 480 4790
rect 560 4780 880 4790
rect 1040 4780 1120 4790
rect 2760 4780 2920 4790
rect 3040 4780 3160 4790
rect 3200 4780 3280 4790
rect 3320 4780 3360 4790
rect 3720 4780 3800 4790
rect 3880 4780 3960 4790
rect 4920 4780 5000 4790
rect 5200 4780 5240 4790
rect 5520 4780 5560 4790
rect 5600 4780 5640 4790
rect 6000 4780 6240 4790
rect 6360 4780 6520 4790
rect 7840 4780 7920 4790
rect 7960 4780 8000 4790
rect 8080 4780 8120 4790
rect 8720 4780 8760 4790
rect 8920 4780 8960 4790
rect 9440 4780 9480 4790
rect 9680 4780 9720 4790
rect 160 4770 360 4780
rect 480 4770 1000 4780
rect 1040 4770 1160 4780
rect 2360 4770 2440 4780
rect 2840 4770 3120 4780
rect 3280 4770 3320 4780
rect 3840 4770 3880 4780
rect 5480 4770 5520 4780
rect 5560 4770 5600 4780
rect 6400 4770 6560 4780
rect 7360 4770 7400 4780
rect 8880 4770 8920 4780
rect 160 4760 360 4770
rect 480 4760 1000 4770
rect 1040 4760 1160 4770
rect 2360 4760 2440 4770
rect 2840 4760 3120 4770
rect 3280 4760 3320 4770
rect 3840 4760 3880 4770
rect 5480 4760 5520 4770
rect 5560 4760 5600 4770
rect 6400 4760 6560 4770
rect 7360 4760 7400 4770
rect 8880 4760 8920 4770
rect 160 4750 360 4760
rect 480 4750 1000 4760
rect 1040 4750 1160 4760
rect 2360 4750 2440 4760
rect 2840 4750 3120 4760
rect 3280 4750 3320 4760
rect 3840 4750 3880 4760
rect 5480 4750 5520 4760
rect 5560 4750 5600 4760
rect 6400 4750 6560 4760
rect 7360 4750 7400 4760
rect 8880 4750 8920 4760
rect 160 4740 360 4750
rect 480 4740 1000 4750
rect 1040 4740 1160 4750
rect 2360 4740 2440 4750
rect 2840 4740 3120 4750
rect 3280 4740 3320 4750
rect 3840 4740 3880 4750
rect 5480 4740 5520 4750
rect 5560 4740 5600 4750
rect 6400 4740 6560 4750
rect 7360 4740 7400 4750
rect 8880 4740 8920 4750
rect 160 4730 440 4740
rect 600 4730 1040 4740
rect 1080 4730 1160 4740
rect 2400 4730 2520 4740
rect 2840 4730 2960 4740
rect 3000 4730 3120 4740
rect 3320 4730 3360 4740
rect 3560 4730 3600 4740
rect 3760 4730 3800 4740
rect 5080 4730 5120 4740
rect 5480 4730 5520 4740
rect 5560 4730 5600 4740
rect 6440 4730 6560 4740
rect 7360 4730 7440 4740
rect 9800 4730 9840 4740
rect 160 4720 440 4730
rect 600 4720 1040 4730
rect 1080 4720 1160 4730
rect 2400 4720 2520 4730
rect 2840 4720 2960 4730
rect 3000 4720 3120 4730
rect 3320 4720 3360 4730
rect 3560 4720 3600 4730
rect 3760 4720 3800 4730
rect 5080 4720 5120 4730
rect 5480 4720 5520 4730
rect 5560 4720 5600 4730
rect 6440 4720 6560 4730
rect 7360 4720 7440 4730
rect 9800 4720 9840 4730
rect 160 4710 440 4720
rect 600 4710 1040 4720
rect 1080 4710 1160 4720
rect 2400 4710 2520 4720
rect 2840 4710 2960 4720
rect 3000 4710 3120 4720
rect 3320 4710 3360 4720
rect 3560 4710 3600 4720
rect 3760 4710 3800 4720
rect 5080 4710 5120 4720
rect 5480 4710 5520 4720
rect 5560 4710 5600 4720
rect 6440 4710 6560 4720
rect 7360 4710 7440 4720
rect 9800 4710 9840 4720
rect 160 4700 440 4710
rect 600 4700 1040 4710
rect 1080 4700 1160 4710
rect 2400 4700 2520 4710
rect 2840 4700 2960 4710
rect 3000 4700 3120 4710
rect 3320 4700 3360 4710
rect 3560 4700 3600 4710
rect 3760 4700 3800 4710
rect 5080 4700 5120 4710
rect 5480 4700 5520 4710
rect 5560 4700 5600 4710
rect 6440 4700 6560 4710
rect 7360 4700 7440 4710
rect 9800 4700 9840 4710
rect 120 4690 520 4700
rect 760 4690 1040 4700
rect 1120 4690 1200 4700
rect 2440 4690 2560 4700
rect 2600 4690 2960 4700
rect 3000 4690 3120 4700
rect 3160 4690 3200 4700
rect 3320 4690 3360 4700
rect 3520 4690 3560 4700
rect 5080 4690 5120 4700
rect 5480 4690 5520 4700
rect 5560 4690 5640 4700
rect 6440 4690 6560 4700
rect 8200 4690 8240 4700
rect 120 4680 520 4690
rect 760 4680 1040 4690
rect 1120 4680 1200 4690
rect 2440 4680 2560 4690
rect 2600 4680 2960 4690
rect 3000 4680 3120 4690
rect 3160 4680 3200 4690
rect 3320 4680 3360 4690
rect 3520 4680 3560 4690
rect 5080 4680 5120 4690
rect 5480 4680 5520 4690
rect 5560 4680 5640 4690
rect 6440 4680 6560 4690
rect 8200 4680 8240 4690
rect 120 4670 520 4680
rect 760 4670 1040 4680
rect 1120 4670 1200 4680
rect 2440 4670 2560 4680
rect 2600 4670 2960 4680
rect 3000 4670 3120 4680
rect 3160 4670 3200 4680
rect 3320 4670 3360 4680
rect 3520 4670 3560 4680
rect 5080 4670 5120 4680
rect 5480 4670 5520 4680
rect 5560 4670 5640 4680
rect 6440 4670 6560 4680
rect 8200 4670 8240 4680
rect 120 4660 520 4670
rect 760 4660 1040 4670
rect 1120 4660 1200 4670
rect 2440 4660 2560 4670
rect 2600 4660 2960 4670
rect 3000 4660 3120 4670
rect 3160 4660 3200 4670
rect 3320 4660 3360 4670
rect 3520 4660 3560 4670
rect 5080 4660 5120 4670
rect 5480 4660 5520 4670
rect 5560 4660 5640 4670
rect 6440 4660 6560 4670
rect 8200 4660 8240 4670
rect 0 4650 600 4660
rect 840 4650 1200 4660
rect 2560 4650 3200 4660
rect 3280 4650 3320 4660
rect 5120 4650 5200 4660
rect 5520 4650 5560 4660
rect 5720 4650 5800 4660
rect 6080 4650 6200 4660
rect 6400 4650 6520 4660
rect 8360 4650 8400 4660
rect 8760 4650 8800 4660
rect 0 4640 600 4650
rect 840 4640 1200 4650
rect 2560 4640 3200 4650
rect 3280 4640 3320 4650
rect 5120 4640 5200 4650
rect 5520 4640 5560 4650
rect 5720 4640 5800 4650
rect 6080 4640 6200 4650
rect 6400 4640 6520 4650
rect 8360 4640 8400 4650
rect 8760 4640 8800 4650
rect 0 4630 600 4640
rect 840 4630 1200 4640
rect 2560 4630 3200 4640
rect 3280 4630 3320 4640
rect 5120 4630 5200 4640
rect 5520 4630 5560 4640
rect 5720 4630 5800 4640
rect 6080 4630 6200 4640
rect 6400 4630 6520 4640
rect 8360 4630 8400 4640
rect 8760 4630 8800 4640
rect 0 4620 600 4630
rect 840 4620 1200 4630
rect 2560 4620 3200 4630
rect 3280 4620 3320 4630
rect 5120 4620 5200 4630
rect 5520 4620 5560 4630
rect 5720 4620 5800 4630
rect 6080 4620 6200 4630
rect 6400 4620 6520 4630
rect 8360 4620 8400 4630
rect 8760 4620 8800 4630
rect 0 4610 680 4620
rect 880 4610 1240 4620
rect 2840 4610 3040 4620
rect 3120 4610 3280 4620
rect 5520 4610 5600 4620
rect 5640 4610 5680 4620
rect 6120 4610 6280 4620
rect 6520 4610 6560 4620
rect 7840 4610 7880 4620
rect 8080 4610 8160 4620
rect 8880 4610 8920 4620
rect 9240 4610 9280 4620
rect 0 4600 680 4610
rect 880 4600 1240 4610
rect 2840 4600 3040 4610
rect 3120 4600 3280 4610
rect 5520 4600 5600 4610
rect 5640 4600 5680 4610
rect 6120 4600 6280 4610
rect 6520 4600 6560 4610
rect 7840 4600 7880 4610
rect 8080 4600 8160 4610
rect 8880 4600 8920 4610
rect 9240 4600 9280 4610
rect 0 4590 680 4600
rect 880 4590 1240 4600
rect 2840 4590 3040 4600
rect 3120 4590 3280 4600
rect 5520 4590 5600 4600
rect 5640 4590 5680 4600
rect 6120 4590 6280 4600
rect 6520 4590 6560 4600
rect 7840 4590 7880 4600
rect 8080 4590 8160 4600
rect 8880 4590 8920 4600
rect 9240 4590 9280 4600
rect 0 4580 680 4590
rect 880 4580 1240 4590
rect 2840 4580 3040 4590
rect 3120 4580 3280 4590
rect 5520 4580 5600 4590
rect 5640 4580 5680 4590
rect 6120 4580 6280 4590
rect 6520 4580 6560 4590
rect 7840 4580 7880 4590
rect 8080 4580 8160 4590
rect 8880 4580 8920 4590
rect 9240 4580 9280 4590
rect 0 4570 720 4580
rect 920 4570 1240 4580
rect 3040 4570 3080 4580
rect 3120 4570 3240 4580
rect 3440 4570 3480 4580
rect 5200 4570 5240 4580
rect 5560 4570 5600 4580
rect 5760 4570 5800 4580
rect 6280 4570 6320 4580
rect 6480 4570 6520 4580
rect 7560 4570 7600 4580
rect 7720 4570 7760 4580
rect 8040 4570 8080 4580
rect 8240 4570 8280 4580
rect 8600 4570 8640 4580
rect 8920 4570 8960 4580
rect 0 4560 720 4570
rect 920 4560 1240 4570
rect 3040 4560 3080 4570
rect 3120 4560 3240 4570
rect 3440 4560 3480 4570
rect 5200 4560 5240 4570
rect 5560 4560 5600 4570
rect 5760 4560 5800 4570
rect 6280 4560 6320 4570
rect 6480 4560 6520 4570
rect 7560 4560 7600 4570
rect 7720 4560 7760 4570
rect 8040 4560 8080 4570
rect 8240 4560 8280 4570
rect 8600 4560 8640 4570
rect 8920 4560 8960 4570
rect 0 4550 720 4560
rect 920 4550 1240 4560
rect 3040 4550 3080 4560
rect 3120 4550 3240 4560
rect 3440 4550 3480 4560
rect 5200 4550 5240 4560
rect 5560 4550 5600 4560
rect 5760 4550 5800 4560
rect 6280 4550 6320 4560
rect 6480 4550 6520 4560
rect 7560 4550 7600 4560
rect 7720 4550 7760 4560
rect 8040 4550 8080 4560
rect 8240 4550 8280 4560
rect 8600 4550 8640 4560
rect 8920 4550 8960 4560
rect 0 4540 720 4550
rect 920 4540 1240 4550
rect 3040 4540 3080 4550
rect 3120 4540 3240 4550
rect 3440 4540 3480 4550
rect 5200 4540 5240 4550
rect 5560 4540 5600 4550
rect 5760 4540 5800 4550
rect 6280 4540 6320 4550
rect 6480 4540 6520 4550
rect 7560 4540 7600 4550
rect 7720 4540 7760 4550
rect 8040 4540 8080 4550
rect 8240 4540 8280 4550
rect 8600 4540 8640 4550
rect 8920 4540 8960 4550
rect 0 4530 760 4540
rect 960 4530 1160 4540
rect 2960 4530 3000 4540
rect 3040 4530 3080 4540
rect 3200 4530 3240 4540
rect 3880 4530 3920 4540
rect 5760 4530 5800 4540
rect 6280 4530 6320 4540
rect 6400 4530 6520 4540
rect 7400 4530 7440 4540
rect 7600 4530 7640 4540
rect 7840 4530 7880 4540
rect 0 4520 760 4530
rect 960 4520 1160 4530
rect 2960 4520 3000 4530
rect 3040 4520 3080 4530
rect 3200 4520 3240 4530
rect 3880 4520 3920 4530
rect 5760 4520 5800 4530
rect 6280 4520 6320 4530
rect 6400 4520 6520 4530
rect 7400 4520 7440 4530
rect 7600 4520 7640 4530
rect 7840 4520 7880 4530
rect 0 4510 760 4520
rect 960 4510 1160 4520
rect 2960 4510 3000 4520
rect 3040 4510 3080 4520
rect 3200 4510 3240 4520
rect 3880 4510 3920 4520
rect 5760 4510 5800 4520
rect 6280 4510 6320 4520
rect 6400 4510 6520 4520
rect 7400 4510 7440 4520
rect 7600 4510 7640 4520
rect 7840 4510 7880 4520
rect 0 4500 760 4510
rect 960 4500 1160 4510
rect 2960 4500 3000 4510
rect 3040 4500 3080 4510
rect 3200 4500 3240 4510
rect 3880 4500 3920 4510
rect 5760 4500 5800 4510
rect 6280 4500 6320 4510
rect 6400 4500 6520 4510
rect 7400 4500 7440 4510
rect 7600 4500 7640 4510
rect 7840 4500 7880 4510
rect 0 4490 640 4500
rect 1000 4490 1200 4500
rect 3040 4490 3080 4500
rect 3840 4490 3960 4500
rect 5760 4490 5800 4500
rect 6240 4490 6280 4500
rect 6360 4490 6520 4500
rect 9960 4490 9990 4500
rect 0 4480 640 4490
rect 1000 4480 1200 4490
rect 3040 4480 3080 4490
rect 3840 4480 3960 4490
rect 5760 4480 5800 4490
rect 6240 4480 6280 4490
rect 6360 4480 6520 4490
rect 9960 4480 9990 4490
rect 0 4470 640 4480
rect 1000 4470 1200 4480
rect 3040 4470 3080 4480
rect 3840 4470 3960 4480
rect 5760 4470 5800 4480
rect 6240 4470 6280 4480
rect 6360 4470 6520 4480
rect 9960 4470 9990 4480
rect 0 4460 640 4470
rect 1000 4460 1200 4470
rect 3040 4460 3080 4470
rect 3840 4460 3960 4470
rect 5760 4460 5800 4470
rect 6240 4460 6280 4470
rect 6360 4460 6520 4470
rect 9960 4460 9990 4470
rect 0 4450 480 4460
rect 520 4450 600 4460
rect 1040 4450 1160 4460
rect 2800 4450 2880 4460
rect 2960 4450 3000 4460
rect 3120 4450 3240 4460
rect 3840 4450 3960 4460
rect 4600 4450 4680 4460
rect 6200 4450 6240 4460
rect 6320 4450 6360 4460
rect 6440 4450 6480 4460
rect 7760 4450 7800 4460
rect 7840 4450 7880 4460
rect 9920 4450 9960 4460
rect 0 4440 480 4450
rect 520 4440 600 4450
rect 1040 4440 1160 4450
rect 2800 4440 2880 4450
rect 2960 4440 3000 4450
rect 3120 4440 3240 4450
rect 3840 4440 3960 4450
rect 4600 4440 4680 4450
rect 6200 4440 6240 4450
rect 6320 4440 6360 4450
rect 6440 4440 6480 4450
rect 7760 4440 7800 4450
rect 7840 4440 7880 4450
rect 9920 4440 9960 4450
rect 0 4430 480 4440
rect 520 4430 600 4440
rect 1040 4430 1160 4440
rect 2800 4430 2880 4440
rect 2960 4430 3000 4440
rect 3120 4430 3240 4440
rect 3840 4430 3960 4440
rect 4600 4430 4680 4440
rect 6200 4430 6240 4440
rect 6320 4430 6360 4440
rect 6440 4430 6480 4440
rect 7760 4430 7800 4440
rect 7840 4430 7880 4440
rect 9920 4430 9960 4440
rect 0 4420 480 4430
rect 520 4420 600 4430
rect 1040 4420 1160 4430
rect 2800 4420 2880 4430
rect 2960 4420 3000 4430
rect 3120 4420 3240 4430
rect 3840 4420 3960 4430
rect 4600 4420 4680 4430
rect 6200 4420 6240 4430
rect 6320 4420 6360 4430
rect 6440 4420 6480 4430
rect 7760 4420 7800 4430
rect 7840 4420 7880 4430
rect 9920 4420 9960 4430
rect 0 4410 280 4420
rect 320 4410 400 4420
rect 2640 4410 2680 4420
rect 2800 4410 2880 4420
rect 3080 4410 3240 4420
rect 3360 4410 3400 4420
rect 3800 4410 3960 4420
rect 4240 4410 4320 4420
rect 4720 4410 4760 4420
rect 4800 4410 4880 4420
rect 5280 4410 5320 4420
rect 6200 4410 6320 4420
rect 8000 4410 8040 4420
rect 8120 4410 8160 4420
rect 8640 4410 8680 4420
rect 9880 4410 9920 4420
rect 0 4400 280 4410
rect 320 4400 400 4410
rect 2640 4400 2680 4410
rect 2800 4400 2880 4410
rect 3080 4400 3240 4410
rect 3360 4400 3400 4410
rect 3800 4400 3960 4410
rect 4240 4400 4320 4410
rect 4720 4400 4760 4410
rect 4800 4400 4880 4410
rect 5280 4400 5320 4410
rect 6200 4400 6320 4410
rect 8000 4400 8040 4410
rect 8120 4400 8160 4410
rect 8640 4400 8680 4410
rect 9880 4400 9920 4410
rect 0 4390 280 4400
rect 320 4390 400 4400
rect 2640 4390 2680 4400
rect 2800 4390 2880 4400
rect 3080 4390 3240 4400
rect 3360 4390 3400 4400
rect 3800 4390 3960 4400
rect 4240 4390 4320 4400
rect 4720 4390 4760 4400
rect 4800 4390 4880 4400
rect 5280 4390 5320 4400
rect 6200 4390 6320 4400
rect 8000 4390 8040 4400
rect 8120 4390 8160 4400
rect 8640 4390 8680 4400
rect 9880 4390 9920 4400
rect 0 4380 280 4390
rect 320 4380 400 4390
rect 2640 4380 2680 4390
rect 2800 4380 2880 4390
rect 3080 4380 3240 4390
rect 3360 4380 3400 4390
rect 3800 4380 3960 4390
rect 4240 4380 4320 4390
rect 4720 4380 4760 4390
rect 4800 4380 4880 4390
rect 5280 4380 5320 4390
rect 6200 4380 6320 4390
rect 8000 4380 8040 4390
rect 8120 4380 8160 4390
rect 8640 4380 8680 4390
rect 9880 4380 9920 4390
rect 0 4370 240 4380
rect 2800 4370 2880 4380
rect 3080 4370 3120 4380
rect 3160 4370 3240 4380
rect 3840 4370 3920 4380
rect 4280 4370 4320 4380
rect 4880 4370 4920 4380
rect 8120 4370 8200 4380
rect 8480 4370 8520 4380
rect 8720 4370 8760 4380
rect 9880 4370 9920 4380
rect 0 4360 240 4370
rect 2800 4360 2880 4370
rect 3080 4360 3120 4370
rect 3160 4360 3240 4370
rect 3840 4360 3920 4370
rect 4280 4360 4320 4370
rect 4880 4360 4920 4370
rect 8120 4360 8200 4370
rect 8480 4360 8520 4370
rect 8720 4360 8760 4370
rect 9880 4360 9920 4370
rect 0 4350 240 4360
rect 2800 4350 2880 4360
rect 3080 4350 3120 4360
rect 3160 4350 3240 4360
rect 3840 4350 3920 4360
rect 4280 4350 4320 4360
rect 4880 4350 4920 4360
rect 8120 4350 8200 4360
rect 8480 4350 8520 4360
rect 8720 4350 8760 4360
rect 9880 4350 9920 4360
rect 0 4340 240 4350
rect 2800 4340 2880 4350
rect 3080 4340 3120 4350
rect 3160 4340 3240 4350
rect 3840 4340 3920 4350
rect 4280 4340 4320 4350
rect 4880 4340 4920 4350
rect 8120 4340 8200 4350
rect 8480 4340 8520 4350
rect 8720 4340 8760 4350
rect 9880 4340 9920 4350
rect 0 4330 240 4340
rect 2800 4330 2880 4340
rect 3080 4330 3160 4340
rect 3240 4330 3280 4340
rect 4160 4330 4280 4340
rect 4520 4330 4560 4340
rect 4920 4330 4960 4340
rect 7360 4330 7400 4340
rect 8160 4330 8200 4340
rect 8520 4330 8560 4340
rect 0 4320 240 4330
rect 2800 4320 2880 4330
rect 3080 4320 3160 4330
rect 3240 4320 3280 4330
rect 4160 4320 4280 4330
rect 4520 4320 4560 4330
rect 4920 4320 4960 4330
rect 7360 4320 7400 4330
rect 8160 4320 8200 4330
rect 8520 4320 8560 4330
rect 0 4310 240 4320
rect 2800 4310 2880 4320
rect 3080 4310 3160 4320
rect 3240 4310 3280 4320
rect 4160 4310 4280 4320
rect 4520 4310 4560 4320
rect 4920 4310 4960 4320
rect 7360 4310 7400 4320
rect 8160 4310 8200 4320
rect 8520 4310 8560 4320
rect 0 4300 240 4310
rect 2800 4300 2880 4310
rect 3080 4300 3160 4310
rect 3240 4300 3280 4310
rect 4160 4300 4280 4310
rect 4520 4300 4560 4310
rect 4920 4300 4960 4310
rect 7360 4300 7400 4310
rect 8160 4300 8200 4310
rect 8520 4300 8560 4310
rect 0 4290 80 4300
rect 2800 4290 2920 4300
rect 3000 4290 3040 4300
rect 3080 4290 3120 4300
rect 3240 4290 3320 4300
rect 4120 4290 4160 4300
rect 4960 4290 5000 4300
rect 5320 4290 5360 4300
rect 7200 4290 7240 4300
rect 8160 4290 8200 4300
rect 8640 4290 8680 4300
rect 8720 4290 8760 4300
rect 0 4280 80 4290
rect 2800 4280 2920 4290
rect 3000 4280 3040 4290
rect 3080 4280 3120 4290
rect 3240 4280 3320 4290
rect 4120 4280 4160 4290
rect 4960 4280 5000 4290
rect 5320 4280 5360 4290
rect 7200 4280 7240 4290
rect 8160 4280 8200 4290
rect 8640 4280 8680 4290
rect 8720 4280 8760 4290
rect 0 4270 80 4280
rect 2800 4270 2920 4280
rect 3000 4270 3040 4280
rect 3080 4270 3120 4280
rect 3240 4270 3320 4280
rect 4120 4270 4160 4280
rect 4960 4270 5000 4280
rect 5320 4270 5360 4280
rect 7200 4270 7240 4280
rect 8160 4270 8200 4280
rect 8640 4270 8680 4280
rect 8720 4270 8760 4280
rect 0 4260 80 4270
rect 2800 4260 2920 4270
rect 3000 4260 3040 4270
rect 3080 4260 3120 4270
rect 3240 4260 3320 4270
rect 4120 4260 4160 4270
rect 4960 4260 5000 4270
rect 5320 4260 5360 4270
rect 7200 4260 7240 4270
rect 8160 4260 8200 4270
rect 8640 4260 8680 4270
rect 8720 4260 8760 4270
rect 0 4250 120 4260
rect 2800 4250 2880 4260
rect 2960 4250 3040 4260
rect 3240 4250 3280 4260
rect 4120 4250 4160 4260
rect 4480 4250 4520 4260
rect 7160 4250 7240 4260
rect 7440 4250 7480 4260
rect 8160 4250 8200 4260
rect 8520 4250 8560 4260
rect 9760 4250 9800 4260
rect 0 4240 120 4250
rect 2800 4240 2880 4250
rect 2960 4240 3040 4250
rect 3240 4240 3280 4250
rect 4120 4240 4160 4250
rect 4480 4240 4520 4250
rect 7160 4240 7240 4250
rect 7440 4240 7480 4250
rect 8160 4240 8200 4250
rect 8520 4240 8560 4250
rect 9760 4240 9800 4250
rect 0 4230 120 4240
rect 2800 4230 2880 4240
rect 2960 4230 3040 4240
rect 3240 4230 3280 4240
rect 4120 4230 4160 4240
rect 4480 4230 4520 4240
rect 7160 4230 7240 4240
rect 7440 4230 7480 4240
rect 8160 4230 8200 4240
rect 8520 4230 8560 4240
rect 9760 4230 9800 4240
rect 0 4220 120 4230
rect 2800 4220 2880 4230
rect 2960 4220 3040 4230
rect 3240 4220 3280 4230
rect 4120 4220 4160 4230
rect 4480 4220 4520 4230
rect 7160 4220 7240 4230
rect 7440 4220 7480 4230
rect 8160 4220 8200 4230
rect 8520 4220 8560 4230
rect 9760 4220 9800 4230
rect 0 4210 120 4220
rect 2560 4210 2600 4220
rect 2760 4210 2800 4220
rect 2840 4210 2960 4220
rect 3000 4210 3040 4220
rect 3240 4210 3280 4220
rect 4080 4210 4120 4220
rect 4400 4210 4440 4220
rect 5000 4210 5040 4220
rect 5360 4210 5400 4220
rect 8160 4210 8200 4220
rect 9280 4210 9320 4220
rect 0 4200 120 4210
rect 2560 4200 2600 4210
rect 2760 4200 2800 4210
rect 2840 4200 2960 4210
rect 3000 4200 3040 4210
rect 3240 4200 3280 4210
rect 4080 4200 4120 4210
rect 4400 4200 4440 4210
rect 5000 4200 5040 4210
rect 5360 4200 5400 4210
rect 8160 4200 8200 4210
rect 9280 4200 9320 4210
rect 0 4190 120 4200
rect 2560 4190 2600 4200
rect 2760 4190 2800 4200
rect 2840 4190 2960 4200
rect 3000 4190 3040 4200
rect 3240 4190 3280 4200
rect 4080 4190 4120 4200
rect 4400 4190 4440 4200
rect 5000 4190 5040 4200
rect 5360 4190 5400 4200
rect 8160 4190 8200 4200
rect 9280 4190 9320 4200
rect 0 4180 120 4190
rect 2560 4180 2600 4190
rect 2760 4180 2800 4190
rect 2840 4180 2960 4190
rect 3000 4180 3040 4190
rect 3240 4180 3280 4190
rect 4080 4180 4120 4190
rect 4400 4180 4440 4190
rect 5000 4180 5040 4190
rect 5360 4180 5400 4190
rect 8160 4180 8200 4190
rect 9280 4180 9320 4190
rect 0 4170 160 4180
rect 2560 4170 2880 4180
rect 2960 4170 3000 4180
rect 3120 4170 3160 4180
rect 3200 4170 3280 4180
rect 5040 4170 5080 4180
rect 0 4160 160 4170
rect 2560 4160 2880 4170
rect 2960 4160 3000 4170
rect 3120 4160 3160 4170
rect 3200 4160 3280 4170
rect 5040 4160 5080 4170
rect 0 4150 160 4160
rect 2560 4150 2880 4160
rect 2960 4150 3000 4160
rect 3120 4150 3160 4160
rect 3200 4150 3280 4160
rect 5040 4150 5080 4160
rect 0 4140 160 4150
rect 2560 4140 2880 4150
rect 2960 4140 3000 4150
rect 3120 4140 3160 4150
rect 3200 4140 3280 4150
rect 5040 4140 5080 4150
rect 80 4130 160 4140
rect 2600 4130 2640 4140
rect 2680 4130 2960 4140
rect 3000 4130 3040 4140
rect 3080 4130 3120 4140
rect 4040 4130 4080 4140
rect 4720 4130 4760 4140
rect 4880 4130 4920 4140
rect 5080 4130 5120 4140
rect 7240 4130 7280 4140
rect 7400 4130 7480 4140
rect 9920 4130 9960 4140
rect 80 4120 160 4130
rect 2600 4120 2640 4130
rect 2680 4120 2960 4130
rect 3000 4120 3040 4130
rect 3080 4120 3120 4130
rect 4040 4120 4080 4130
rect 4720 4120 4760 4130
rect 4880 4120 4920 4130
rect 5080 4120 5120 4130
rect 7240 4120 7280 4130
rect 7400 4120 7480 4130
rect 9920 4120 9960 4130
rect 80 4110 160 4120
rect 2600 4110 2640 4120
rect 2680 4110 2960 4120
rect 3000 4110 3040 4120
rect 3080 4110 3120 4120
rect 4040 4110 4080 4120
rect 4720 4110 4760 4120
rect 4880 4110 4920 4120
rect 5080 4110 5120 4120
rect 7240 4110 7280 4120
rect 7400 4110 7480 4120
rect 9920 4110 9960 4120
rect 80 4100 160 4110
rect 2600 4100 2640 4110
rect 2680 4100 2960 4110
rect 3000 4100 3040 4110
rect 3080 4100 3120 4110
rect 4040 4100 4080 4110
rect 4720 4100 4760 4110
rect 4880 4100 4920 4110
rect 5080 4100 5120 4110
rect 7240 4100 7280 4110
rect 7400 4100 7480 4110
rect 9920 4100 9960 4110
rect 120 4090 160 4100
rect 2600 4090 3080 4100
rect 4640 4090 4680 4100
rect 5120 4090 5160 4100
rect 5400 4090 5440 4100
rect 5640 4090 5680 4100
rect 7480 4090 7600 4100
rect 8760 4090 8800 4100
rect 120 4080 160 4090
rect 2600 4080 3080 4090
rect 4640 4080 4680 4090
rect 5120 4080 5160 4090
rect 5400 4080 5440 4090
rect 5640 4080 5680 4090
rect 7480 4080 7600 4090
rect 8760 4080 8800 4090
rect 120 4070 160 4080
rect 2600 4070 3080 4080
rect 4640 4070 4680 4080
rect 5120 4070 5160 4080
rect 5400 4070 5440 4080
rect 5640 4070 5680 4080
rect 7480 4070 7600 4080
rect 8760 4070 8800 4080
rect 120 4060 160 4070
rect 2600 4060 3080 4070
rect 4640 4060 4680 4070
rect 5120 4060 5160 4070
rect 5400 4060 5440 4070
rect 5640 4060 5680 4070
rect 7480 4060 7600 4070
rect 8760 4060 8800 4070
rect 2600 4050 2960 4060
rect 3000 4050 3040 4060
rect 4000 4050 4040 4060
rect 5120 4050 5160 4060
rect 5680 4050 5720 4060
rect 7200 4050 7240 4060
rect 7600 4050 7760 4060
rect 2600 4040 2960 4050
rect 3000 4040 3040 4050
rect 4000 4040 4040 4050
rect 5120 4040 5160 4050
rect 5680 4040 5720 4050
rect 7200 4040 7240 4050
rect 7600 4040 7760 4050
rect 2600 4030 2960 4040
rect 3000 4030 3040 4040
rect 4000 4030 4040 4040
rect 5120 4030 5160 4040
rect 5680 4030 5720 4040
rect 7200 4030 7240 4040
rect 7600 4030 7760 4040
rect 2600 4020 2960 4030
rect 3000 4020 3040 4030
rect 4000 4020 4040 4030
rect 5120 4020 5160 4030
rect 5680 4020 5720 4030
rect 7200 4020 7240 4030
rect 7600 4020 7760 4030
rect 2600 4010 3080 4020
rect 4640 4010 4680 4020
rect 5720 4010 5760 4020
rect 7720 4010 7840 4020
rect 8400 4010 8440 4020
rect 2600 4000 3080 4010
rect 4640 4000 4680 4010
rect 5720 4000 5760 4010
rect 7720 4000 7840 4010
rect 8400 4000 8440 4010
rect 2600 3990 3080 4000
rect 4640 3990 4680 4000
rect 5720 3990 5760 4000
rect 7720 3990 7840 4000
rect 8400 3990 8440 4000
rect 2600 3980 3080 3990
rect 4640 3980 4680 3990
rect 5720 3980 5760 3990
rect 7720 3980 7840 3990
rect 8400 3980 8440 3990
rect 2600 3970 3120 3980
rect 3920 3970 3960 3980
rect 5160 3970 5200 3980
rect 5480 3970 5520 3980
rect 5800 3970 6000 3980
rect 6240 3970 6320 3980
rect 7160 3970 7200 3980
rect 7880 3970 7960 3980
rect 8120 3970 8160 3980
rect 8520 3970 8560 3980
rect 2600 3960 3120 3970
rect 3920 3960 3960 3970
rect 5160 3960 5200 3970
rect 5480 3960 5520 3970
rect 5800 3960 6000 3970
rect 6240 3960 6320 3970
rect 7160 3960 7200 3970
rect 7880 3960 7960 3970
rect 8120 3960 8160 3970
rect 8520 3960 8560 3970
rect 2600 3950 3120 3960
rect 3920 3950 3960 3960
rect 5160 3950 5200 3960
rect 5480 3950 5520 3960
rect 5800 3950 6000 3960
rect 6240 3950 6320 3960
rect 7160 3950 7200 3960
rect 7880 3950 7960 3960
rect 8120 3950 8160 3960
rect 8520 3950 8560 3960
rect 2600 3940 3120 3950
rect 3920 3940 3960 3950
rect 5160 3940 5200 3950
rect 5480 3940 5520 3950
rect 5800 3940 6000 3950
rect 6240 3940 6320 3950
rect 7160 3940 7200 3950
rect 7880 3940 7960 3950
rect 8120 3940 8160 3950
rect 8520 3940 8560 3950
rect 2600 3930 2920 3940
rect 2960 3930 3040 3940
rect 3880 3930 3920 3940
rect 4200 3930 4280 3940
rect 5200 3930 5240 3940
rect 5400 3930 5480 3940
rect 6040 3930 6320 3940
rect 7920 3930 7960 3940
rect 8080 3930 8120 3940
rect 8520 3930 8560 3940
rect 8640 3930 8680 3940
rect 2600 3920 2920 3930
rect 2960 3920 3040 3930
rect 3880 3920 3920 3930
rect 4200 3920 4280 3930
rect 5200 3920 5240 3930
rect 5400 3920 5480 3930
rect 6040 3920 6320 3930
rect 7920 3920 7960 3930
rect 8080 3920 8120 3930
rect 8520 3920 8560 3930
rect 8640 3920 8680 3930
rect 2600 3910 2920 3920
rect 2960 3910 3040 3920
rect 3880 3910 3920 3920
rect 4200 3910 4280 3920
rect 5200 3910 5240 3920
rect 5400 3910 5480 3920
rect 6040 3910 6320 3920
rect 7920 3910 7960 3920
rect 8080 3910 8120 3920
rect 8520 3910 8560 3920
rect 8640 3910 8680 3920
rect 2600 3900 2920 3910
rect 2960 3900 3040 3910
rect 3880 3900 3920 3910
rect 4200 3900 4280 3910
rect 5200 3900 5240 3910
rect 5400 3900 5480 3910
rect 6040 3900 6320 3910
rect 7920 3900 7960 3910
rect 8080 3900 8120 3910
rect 8520 3900 8560 3910
rect 8640 3900 8680 3910
rect 2520 3890 2880 3900
rect 4120 3890 4280 3900
rect 6000 3890 6320 3900
rect 7960 3890 8000 3900
rect 9600 3890 9680 3900
rect 2520 3880 2880 3890
rect 4120 3880 4280 3890
rect 6000 3880 6320 3890
rect 7960 3880 8000 3890
rect 9600 3880 9680 3890
rect 2520 3870 2880 3880
rect 4120 3870 4280 3880
rect 6000 3870 6320 3880
rect 7960 3870 8000 3880
rect 9600 3870 9680 3880
rect 2520 3860 2880 3870
rect 4120 3860 4280 3870
rect 6000 3860 6320 3870
rect 7960 3860 8000 3870
rect 9600 3860 9680 3870
rect 2240 3850 2280 3860
rect 2400 3850 2480 3860
rect 2560 3850 2880 3860
rect 3840 3850 3880 3860
rect 4120 3850 4160 3860
rect 4240 3850 4280 3860
rect 5240 3850 5280 3860
rect 5960 3850 6320 3860
rect 8000 3850 8120 3860
rect 8160 3850 8240 3860
rect 9600 3850 9640 3860
rect 9680 3850 9720 3860
rect 2240 3840 2280 3850
rect 2400 3840 2480 3850
rect 2560 3840 2880 3850
rect 3840 3840 3880 3850
rect 4120 3840 4160 3850
rect 4240 3840 4280 3850
rect 5240 3840 5280 3850
rect 5960 3840 6320 3850
rect 8000 3840 8120 3850
rect 8160 3840 8240 3850
rect 9600 3840 9640 3850
rect 9680 3840 9720 3850
rect 2240 3830 2280 3840
rect 2400 3830 2480 3840
rect 2560 3830 2880 3840
rect 3840 3830 3880 3840
rect 4120 3830 4160 3840
rect 4240 3830 4280 3840
rect 5240 3830 5280 3840
rect 5960 3830 6320 3840
rect 8000 3830 8120 3840
rect 8160 3830 8240 3840
rect 9600 3830 9640 3840
rect 9680 3830 9720 3840
rect 2240 3820 2280 3830
rect 2400 3820 2480 3830
rect 2560 3820 2880 3830
rect 3840 3820 3880 3830
rect 4120 3820 4160 3830
rect 4240 3820 4280 3830
rect 5240 3820 5280 3830
rect 5960 3820 6320 3830
rect 8000 3820 8120 3830
rect 8160 3820 8240 3830
rect 9600 3820 9640 3830
rect 9680 3820 9720 3830
rect 2600 3810 2920 3820
rect 3840 3810 3880 3820
rect 4240 3810 4280 3820
rect 5960 3810 6280 3820
rect 7080 3810 7120 3820
rect 8080 3810 8120 3820
rect 8160 3810 8200 3820
rect 9680 3810 9720 3820
rect 2600 3800 2920 3810
rect 3840 3800 3880 3810
rect 4240 3800 4280 3810
rect 5960 3800 6280 3810
rect 7080 3800 7120 3810
rect 8080 3800 8120 3810
rect 8160 3800 8200 3810
rect 9680 3800 9720 3810
rect 2600 3790 2920 3800
rect 3840 3790 3880 3800
rect 4240 3790 4280 3800
rect 5960 3790 6280 3800
rect 7080 3790 7120 3800
rect 8080 3790 8120 3800
rect 8160 3790 8200 3800
rect 9680 3790 9720 3800
rect 2600 3780 2920 3790
rect 3840 3780 3880 3790
rect 4240 3780 4280 3790
rect 5960 3780 6280 3790
rect 7080 3780 7120 3790
rect 8080 3780 8120 3790
rect 8160 3780 8200 3790
rect 9680 3780 9720 3790
rect 1640 3770 1720 3780
rect 2560 3770 2600 3780
rect 2640 3770 2920 3780
rect 3280 3770 3320 3780
rect 4000 3770 4040 3780
rect 4080 3770 4120 3780
rect 5280 3770 5320 3780
rect 6000 3770 6320 3780
rect 8120 3770 8160 3780
rect 8320 3770 8360 3780
rect 9680 3770 9720 3780
rect 1640 3760 1720 3770
rect 2560 3760 2600 3770
rect 2640 3760 2920 3770
rect 3280 3760 3320 3770
rect 4000 3760 4040 3770
rect 4080 3760 4120 3770
rect 5280 3760 5320 3770
rect 6000 3760 6320 3770
rect 8120 3760 8160 3770
rect 8320 3760 8360 3770
rect 9680 3760 9720 3770
rect 1640 3750 1720 3760
rect 2560 3750 2600 3760
rect 2640 3750 2920 3760
rect 3280 3750 3320 3760
rect 4000 3750 4040 3760
rect 4080 3750 4120 3760
rect 5280 3750 5320 3760
rect 6000 3750 6320 3760
rect 8120 3750 8160 3760
rect 8320 3750 8360 3760
rect 9680 3750 9720 3760
rect 1640 3740 1720 3750
rect 2560 3740 2600 3750
rect 2640 3740 2920 3750
rect 3280 3740 3320 3750
rect 4000 3740 4040 3750
rect 4080 3740 4120 3750
rect 5280 3740 5320 3750
rect 6000 3740 6320 3750
rect 8120 3740 8160 3750
rect 8320 3740 8360 3750
rect 9680 3740 9720 3750
rect 1600 3730 1720 3740
rect 2760 3730 2880 3740
rect 3960 3730 4040 3740
rect 5280 3730 5320 3740
rect 6040 3730 6440 3740
rect 1600 3720 1720 3730
rect 2760 3720 2880 3730
rect 3960 3720 4040 3730
rect 5280 3720 5320 3730
rect 6040 3720 6440 3730
rect 1600 3710 1720 3720
rect 2760 3710 2880 3720
rect 3960 3710 4040 3720
rect 5280 3710 5320 3720
rect 6040 3710 6440 3720
rect 1600 3700 1720 3710
rect 2760 3700 2880 3710
rect 3960 3700 4040 3710
rect 5280 3700 5320 3710
rect 6040 3700 6440 3710
rect 0 3690 40 3700
rect 1600 3690 1720 3700
rect 2880 3690 2960 3700
rect 3000 3690 3040 3700
rect 3320 3690 3360 3700
rect 6080 3690 6480 3700
rect 7000 3690 7040 3700
rect 8400 3690 8480 3700
rect 0 3680 40 3690
rect 1600 3680 1720 3690
rect 2880 3680 2960 3690
rect 3000 3680 3040 3690
rect 3320 3680 3360 3690
rect 6080 3680 6480 3690
rect 7000 3680 7040 3690
rect 8400 3680 8480 3690
rect 0 3670 40 3680
rect 1600 3670 1720 3680
rect 2880 3670 2960 3680
rect 3000 3670 3040 3680
rect 3320 3670 3360 3680
rect 6080 3670 6480 3680
rect 7000 3670 7040 3680
rect 8400 3670 8480 3680
rect 0 3660 40 3670
rect 1600 3660 1720 3670
rect 2880 3660 2960 3670
rect 3000 3660 3040 3670
rect 3320 3660 3360 3670
rect 6080 3660 6480 3670
rect 7000 3660 7040 3670
rect 8400 3660 8480 3670
rect 1680 3650 1720 3660
rect 3080 3650 3120 3660
rect 3320 3650 3360 3660
rect 3920 3650 3960 3660
rect 5320 3650 5360 3660
rect 6160 3650 6440 3660
rect 6960 3650 7000 3660
rect 8400 3650 8440 3660
rect 8480 3650 8520 3660
rect 1680 3640 1720 3650
rect 3080 3640 3120 3650
rect 3320 3640 3360 3650
rect 3920 3640 3960 3650
rect 5320 3640 5360 3650
rect 6160 3640 6440 3650
rect 6960 3640 7000 3650
rect 8400 3640 8440 3650
rect 8480 3640 8520 3650
rect 1680 3630 1720 3640
rect 3080 3630 3120 3640
rect 3320 3630 3360 3640
rect 3920 3630 3960 3640
rect 5320 3630 5360 3640
rect 6160 3630 6440 3640
rect 6960 3630 7000 3640
rect 8400 3630 8440 3640
rect 8480 3630 8520 3640
rect 1680 3620 1720 3630
rect 3080 3620 3120 3630
rect 3320 3620 3360 3630
rect 3920 3620 3960 3630
rect 5320 3620 5360 3630
rect 6160 3620 6440 3630
rect 6960 3620 7000 3630
rect 8400 3620 8440 3630
rect 8480 3620 8520 3630
rect 1680 3610 1720 3620
rect 3200 3610 3240 3620
rect 3360 3610 3400 3620
rect 5320 3610 5360 3620
rect 6160 3610 6440 3620
rect 8400 3610 8440 3620
rect 1680 3600 1720 3610
rect 3200 3600 3240 3610
rect 3360 3600 3400 3610
rect 5320 3600 5360 3610
rect 6160 3600 6440 3610
rect 8400 3600 8440 3610
rect 1680 3590 1720 3600
rect 3200 3590 3240 3600
rect 3360 3590 3400 3600
rect 5320 3590 5360 3600
rect 6160 3590 6440 3600
rect 8400 3590 8440 3600
rect 1680 3580 1720 3590
rect 3200 3580 3240 3590
rect 3360 3580 3400 3590
rect 5320 3580 5360 3590
rect 6160 3580 6440 3590
rect 8400 3580 8440 3590
rect 1440 3570 1480 3580
rect 1680 3570 1720 3580
rect 3880 3570 3920 3580
rect 5320 3570 5360 3580
rect 6160 3570 6360 3580
rect 8280 3570 8320 3580
rect 8440 3570 8480 3580
rect 9440 3570 9480 3580
rect 1440 3560 1480 3570
rect 1680 3560 1720 3570
rect 3880 3560 3920 3570
rect 5320 3560 5360 3570
rect 6160 3560 6360 3570
rect 8280 3560 8320 3570
rect 8440 3560 8480 3570
rect 9440 3560 9480 3570
rect 1440 3550 1480 3560
rect 1680 3550 1720 3560
rect 3880 3550 3920 3560
rect 5320 3550 5360 3560
rect 6160 3550 6360 3560
rect 8280 3550 8320 3560
rect 8440 3550 8480 3560
rect 9440 3550 9480 3560
rect 1440 3540 1480 3550
rect 1680 3540 1720 3550
rect 3880 3540 3920 3550
rect 5320 3540 5360 3550
rect 6160 3540 6360 3550
rect 8280 3540 8320 3550
rect 8440 3540 8480 3550
rect 9440 3540 9480 3550
rect 1440 3530 1480 3540
rect 2520 3530 2600 3540
rect 3400 3530 3440 3540
rect 5320 3530 5360 3540
rect 6160 3530 6360 3540
rect 8440 3530 8480 3540
rect 1440 3520 1480 3530
rect 2520 3520 2600 3530
rect 3400 3520 3440 3530
rect 5320 3520 5360 3530
rect 6160 3520 6360 3530
rect 8440 3520 8480 3530
rect 1440 3510 1480 3520
rect 2520 3510 2600 3520
rect 3400 3510 3440 3520
rect 5320 3510 5360 3520
rect 6160 3510 6360 3520
rect 8440 3510 8480 3520
rect 1440 3500 1480 3510
rect 2520 3500 2600 3510
rect 3400 3500 3440 3510
rect 5320 3500 5360 3510
rect 6160 3500 6360 3510
rect 8440 3500 8480 3510
rect 1400 3490 1480 3500
rect 2360 3490 2400 3500
rect 2760 3490 2840 3500
rect 3320 3490 3360 3500
rect 3920 3490 3960 3500
rect 4960 3490 5040 3500
rect 5320 3490 5360 3500
rect 6160 3490 6320 3500
rect 6840 3490 6880 3500
rect 8360 3490 8400 3500
rect 8480 3490 8520 3500
rect 9240 3490 9320 3500
rect 1400 3480 1480 3490
rect 2360 3480 2400 3490
rect 2760 3480 2840 3490
rect 3320 3480 3360 3490
rect 3920 3480 3960 3490
rect 4960 3480 5040 3490
rect 5320 3480 5360 3490
rect 6160 3480 6320 3490
rect 6840 3480 6880 3490
rect 8360 3480 8400 3490
rect 8480 3480 8520 3490
rect 9240 3480 9320 3490
rect 1400 3470 1480 3480
rect 2360 3470 2400 3480
rect 2760 3470 2840 3480
rect 3320 3470 3360 3480
rect 3920 3470 3960 3480
rect 4960 3470 5040 3480
rect 5320 3470 5360 3480
rect 6160 3470 6320 3480
rect 6840 3470 6880 3480
rect 8360 3470 8400 3480
rect 8480 3470 8520 3480
rect 9240 3470 9320 3480
rect 1400 3460 1480 3470
rect 2360 3460 2400 3470
rect 2760 3460 2840 3470
rect 3320 3460 3360 3470
rect 3920 3460 3960 3470
rect 4960 3460 5040 3470
rect 5320 3460 5360 3470
rect 6160 3460 6320 3470
rect 6840 3460 6880 3470
rect 8360 3460 8400 3470
rect 8480 3460 8520 3470
rect 9240 3460 9320 3470
rect 1400 3450 1440 3460
rect 2240 3450 2280 3460
rect 2920 3450 2960 3460
rect 3360 3450 3440 3460
rect 3920 3450 3960 3460
rect 4440 3450 4680 3460
rect 5320 3450 5360 3460
rect 5840 3450 6000 3460
rect 6120 3450 6280 3460
rect 6800 3450 6840 3460
rect 8440 3450 8520 3460
rect 9200 3450 9240 3460
rect 1400 3440 1440 3450
rect 2240 3440 2280 3450
rect 2920 3440 2960 3450
rect 3360 3440 3440 3450
rect 3920 3440 3960 3450
rect 4440 3440 4680 3450
rect 5320 3440 5360 3450
rect 5840 3440 6000 3450
rect 6120 3440 6280 3450
rect 6800 3440 6840 3450
rect 8440 3440 8520 3450
rect 9200 3440 9240 3450
rect 1400 3430 1440 3440
rect 2240 3430 2280 3440
rect 2920 3430 2960 3440
rect 3360 3430 3440 3440
rect 3920 3430 3960 3440
rect 4440 3430 4680 3440
rect 5320 3430 5360 3440
rect 5840 3430 6000 3440
rect 6120 3430 6280 3440
rect 6800 3430 6840 3440
rect 8440 3430 8520 3440
rect 9200 3430 9240 3440
rect 1400 3420 1440 3430
rect 2240 3420 2280 3430
rect 2920 3420 2960 3430
rect 3360 3420 3440 3430
rect 3920 3420 3960 3430
rect 4440 3420 4680 3430
rect 5320 3420 5360 3430
rect 5840 3420 6000 3430
rect 6120 3420 6280 3430
rect 6800 3420 6840 3430
rect 8440 3420 8520 3430
rect 9200 3420 9240 3430
rect 1360 3410 1440 3420
rect 3000 3410 3040 3420
rect 4280 3410 4320 3420
rect 4480 3410 4560 3420
rect 4840 3410 4920 3420
rect 5320 3410 5360 3420
rect 5680 3410 5720 3420
rect 5840 3410 6080 3420
rect 6120 3410 6200 3420
rect 6760 3410 6800 3420
rect 8480 3410 8520 3420
rect 9120 3410 9160 3420
rect 1360 3400 1440 3410
rect 3000 3400 3040 3410
rect 4280 3400 4320 3410
rect 4480 3400 4560 3410
rect 4840 3400 4920 3410
rect 5320 3400 5360 3410
rect 5680 3400 5720 3410
rect 5840 3400 6080 3410
rect 6120 3400 6200 3410
rect 6760 3400 6800 3410
rect 8480 3400 8520 3410
rect 9120 3400 9160 3410
rect 1360 3390 1440 3400
rect 3000 3390 3040 3400
rect 4280 3390 4320 3400
rect 4480 3390 4560 3400
rect 4840 3390 4920 3400
rect 5320 3390 5360 3400
rect 5680 3390 5720 3400
rect 5840 3390 6080 3400
rect 6120 3390 6200 3400
rect 6760 3390 6800 3400
rect 8480 3390 8520 3400
rect 9120 3390 9160 3400
rect 1360 3380 1440 3390
rect 3000 3380 3040 3390
rect 4280 3380 4320 3390
rect 4480 3380 4560 3390
rect 4840 3380 4920 3390
rect 5320 3380 5360 3390
rect 5680 3380 5720 3390
rect 5840 3380 6080 3390
rect 6120 3380 6200 3390
rect 6760 3380 6800 3390
rect 8480 3380 8520 3390
rect 9120 3380 9160 3390
rect 1360 3370 1440 3380
rect 2120 3370 2160 3380
rect 3480 3370 3520 3380
rect 3560 3370 3600 3380
rect 3960 3370 4000 3380
rect 4280 3370 4320 3380
rect 4720 3370 4800 3380
rect 4840 3370 4880 3380
rect 5320 3370 5360 3380
rect 5640 3370 5760 3380
rect 5840 3370 6080 3380
rect 6120 3370 6160 3380
rect 8480 3370 8520 3380
rect 9080 3370 9160 3380
rect 1360 3360 1440 3370
rect 2120 3360 2160 3370
rect 3480 3360 3520 3370
rect 3560 3360 3600 3370
rect 3960 3360 4000 3370
rect 4280 3360 4320 3370
rect 4720 3360 4800 3370
rect 4840 3360 4880 3370
rect 5320 3360 5360 3370
rect 5640 3360 5760 3370
rect 5840 3360 6080 3370
rect 6120 3360 6160 3370
rect 8480 3360 8520 3370
rect 9080 3360 9160 3370
rect 1360 3350 1440 3360
rect 2120 3350 2160 3360
rect 3480 3350 3520 3360
rect 3560 3350 3600 3360
rect 3960 3350 4000 3360
rect 4280 3350 4320 3360
rect 4720 3350 4800 3360
rect 4840 3350 4880 3360
rect 5320 3350 5360 3360
rect 5640 3350 5760 3360
rect 5840 3350 6080 3360
rect 6120 3350 6160 3360
rect 8480 3350 8520 3360
rect 9080 3350 9160 3360
rect 1360 3340 1440 3350
rect 2120 3340 2160 3350
rect 3480 3340 3520 3350
rect 3560 3340 3600 3350
rect 3960 3340 4000 3350
rect 4280 3340 4320 3350
rect 4720 3340 4800 3350
rect 4840 3340 4880 3350
rect 5320 3340 5360 3350
rect 5640 3340 5760 3350
rect 5840 3340 6080 3350
rect 6120 3340 6160 3350
rect 8480 3340 8520 3350
rect 9080 3340 9160 3350
rect 1320 3330 1400 3340
rect 2080 3330 2120 3340
rect 3480 3330 3520 3340
rect 3960 3330 4040 3340
rect 4240 3330 4320 3340
rect 4600 3330 4800 3340
rect 5600 3330 5800 3340
rect 5840 3330 6160 3340
rect 9080 3330 9120 3340
rect 1320 3320 1400 3330
rect 2080 3320 2120 3330
rect 3480 3320 3520 3330
rect 3960 3320 4040 3330
rect 4240 3320 4320 3330
rect 4600 3320 4800 3330
rect 5600 3320 5800 3330
rect 5840 3320 6160 3330
rect 9080 3320 9120 3330
rect 1320 3310 1400 3320
rect 2080 3310 2120 3320
rect 3480 3310 3520 3320
rect 3960 3310 4040 3320
rect 4240 3310 4320 3320
rect 4600 3310 4800 3320
rect 5600 3310 5800 3320
rect 5840 3310 6160 3320
rect 9080 3310 9120 3320
rect 1320 3300 1400 3310
rect 2080 3300 2120 3310
rect 3480 3300 3520 3310
rect 3960 3300 4040 3310
rect 4240 3300 4320 3310
rect 4600 3300 4800 3310
rect 5600 3300 5800 3310
rect 5840 3300 6160 3310
rect 9080 3300 9120 3310
rect 1320 3290 1400 3300
rect 3120 3290 3160 3300
rect 3520 3290 3600 3300
rect 4000 3290 4080 3300
rect 4240 3290 4320 3300
rect 4520 3290 4600 3300
rect 4680 3290 4720 3300
rect 5600 3290 6160 3300
rect 9640 3290 9680 3300
rect 1320 3280 1400 3290
rect 3120 3280 3160 3290
rect 3520 3280 3600 3290
rect 4000 3280 4080 3290
rect 4240 3280 4320 3290
rect 4520 3280 4600 3290
rect 4680 3280 4720 3290
rect 5600 3280 6160 3290
rect 9640 3280 9680 3290
rect 1320 3270 1400 3280
rect 3120 3270 3160 3280
rect 3520 3270 3600 3280
rect 4000 3270 4080 3280
rect 4240 3270 4320 3280
rect 4520 3270 4600 3280
rect 4680 3270 4720 3280
rect 5600 3270 6160 3280
rect 9640 3270 9680 3280
rect 1320 3260 1400 3270
rect 3120 3260 3160 3270
rect 3520 3260 3600 3270
rect 4000 3260 4080 3270
rect 4240 3260 4320 3270
rect 4520 3260 4600 3270
rect 4680 3260 4720 3270
rect 5600 3260 6160 3270
rect 9640 3260 9680 3270
rect 1280 3250 1400 3260
rect 2040 3250 2080 3260
rect 3600 3250 3640 3260
rect 4040 3250 4120 3260
rect 4280 3250 4360 3260
rect 4400 3250 4440 3260
rect 4600 3250 4640 3260
rect 5280 3250 5320 3260
rect 5640 3250 6200 3260
rect 6520 3250 6600 3260
rect 6640 3250 6680 3260
rect 9360 3250 9400 3260
rect 1280 3240 1400 3250
rect 2040 3240 2080 3250
rect 3600 3240 3640 3250
rect 4040 3240 4120 3250
rect 4280 3240 4360 3250
rect 4400 3240 4440 3250
rect 4600 3240 4640 3250
rect 5280 3240 5320 3250
rect 5640 3240 6200 3250
rect 6520 3240 6600 3250
rect 6640 3240 6680 3250
rect 9360 3240 9400 3250
rect 1280 3230 1400 3240
rect 2040 3230 2080 3240
rect 3600 3230 3640 3240
rect 4040 3230 4120 3240
rect 4280 3230 4360 3240
rect 4400 3230 4440 3240
rect 4600 3230 4640 3240
rect 5280 3230 5320 3240
rect 5640 3230 6200 3240
rect 6520 3230 6600 3240
rect 6640 3230 6680 3240
rect 9360 3230 9400 3240
rect 1280 3220 1400 3230
rect 2040 3220 2080 3230
rect 3600 3220 3640 3230
rect 4040 3220 4120 3230
rect 4280 3220 4360 3230
rect 4400 3220 4440 3230
rect 4600 3220 4640 3230
rect 5280 3220 5320 3230
rect 5640 3220 6200 3230
rect 6520 3220 6600 3230
rect 6640 3220 6680 3230
rect 9360 3220 9400 3230
rect 1280 3210 1360 3220
rect 2040 3210 2080 3220
rect 3160 3210 3200 3220
rect 3560 3210 3600 3220
rect 4040 3210 4160 3220
rect 4280 3210 4360 3220
rect 4480 3210 4520 3220
rect 4920 3210 4960 3220
rect 5280 3210 5320 3220
rect 5680 3210 6200 3220
rect 6440 3210 6480 3220
rect 6560 3210 6600 3220
rect 6640 3210 6680 3220
rect 9120 3210 9160 3220
rect 9520 3210 9600 3220
rect 1280 3200 1360 3210
rect 2040 3200 2080 3210
rect 3160 3200 3200 3210
rect 3560 3200 3600 3210
rect 4040 3200 4160 3210
rect 4280 3200 4360 3210
rect 4480 3200 4520 3210
rect 4920 3200 4960 3210
rect 5280 3200 5320 3210
rect 5680 3200 6200 3210
rect 6440 3200 6480 3210
rect 6560 3200 6600 3210
rect 6640 3200 6680 3210
rect 9120 3200 9160 3210
rect 9520 3200 9600 3210
rect 1280 3190 1360 3200
rect 2040 3190 2080 3200
rect 3160 3190 3200 3200
rect 3560 3190 3600 3200
rect 4040 3190 4160 3200
rect 4280 3190 4360 3200
rect 4480 3190 4520 3200
rect 4920 3190 4960 3200
rect 5280 3190 5320 3200
rect 5680 3190 6200 3200
rect 6440 3190 6480 3200
rect 6560 3190 6600 3200
rect 6640 3190 6680 3200
rect 9120 3190 9160 3200
rect 9520 3190 9600 3200
rect 1280 3180 1360 3190
rect 2040 3180 2080 3190
rect 3160 3180 3200 3190
rect 3560 3180 3600 3190
rect 4040 3180 4160 3190
rect 4280 3180 4360 3190
rect 4480 3180 4520 3190
rect 4920 3180 4960 3190
rect 5280 3180 5320 3190
rect 5680 3180 6200 3190
rect 6440 3180 6480 3190
rect 6560 3180 6600 3190
rect 6640 3180 6680 3190
rect 9120 3180 9160 3190
rect 9520 3180 9600 3190
rect 1240 3170 1360 3180
rect 4080 3170 4160 3180
rect 4400 3170 4480 3180
rect 4880 3170 4920 3180
rect 5720 3170 6240 3180
rect 6320 3170 6360 3180
rect 6560 3170 6600 3180
rect 9080 3170 9120 3180
rect 9240 3170 9280 3180
rect 9480 3170 9520 3180
rect 1240 3160 1360 3170
rect 4080 3160 4160 3170
rect 4400 3160 4480 3170
rect 4880 3160 4920 3170
rect 5720 3160 6240 3170
rect 6320 3160 6360 3170
rect 6560 3160 6600 3170
rect 9080 3160 9120 3170
rect 9240 3160 9280 3170
rect 9480 3160 9520 3170
rect 1240 3150 1360 3160
rect 4080 3150 4160 3160
rect 4400 3150 4480 3160
rect 4880 3150 4920 3160
rect 5720 3150 6240 3160
rect 6320 3150 6360 3160
rect 6560 3150 6600 3160
rect 9080 3150 9120 3160
rect 9240 3150 9280 3160
rect 9480 3150 9520 3160
rect 1240 3140 1360 3150
rect 4080 3140 4160 3150
rect 4400 3140 4480 3150
rect 4880 3140 4920 3150
rect 5720 3140 6240 3150
rect 6320 3140 6360 3150
rect 6560 3140 6600 3150
rect 9080 3140 9120 3150
rect 9240 3140 9280 3150
rect 9480 3140 9520 3150
rect 1240 3130 1360 3140
rect 2000 3130 2040 3140
rect 3760 3130 3920 3140
rect 4080 3130 4200 3140
rect 4480 3130 4520 3140
rect 4840 3130 4920 3140
rect 5880 3130 6120 3140
rect 6600 3130 6640 3140
rect 9080 3130 9120 3140
rect 9200 3130 9240 3140
rect 9440 3130 9520 3140
rect 1240 3120 1360 3130
rect 2000 3120 2040 3130
rect 3760 3120 3920 3130
rect 4080 3120 4200 3130
rect 4480 3120 4520 3130
rect 4840 3120 4920 3130
rect 5880 3120 6120 3130
rect 6600 3120 6640 3130
rect 9080 3120 9120 3130
rect 9200 3120 9240 3130
rect 9440 3120 9520 3130
rect 1240 3110 1360 3120
rect 2000 3110 2040 3120
rect 3760 3110 3920 3120
rect 4080 3110 4200 3120
rect 4480 3110 4520 3120
rect 4840 3110 4920 3120
rect 5880 3110 6120 3120
rect 6600 3110 6640 3120
rect 9080 3110 9120 3120
rect 9200 3110 9240 3120
rect 9440 3110 9520 3120
rect 1240 3100 1360 3110
rect 2000 3100 2040 3110
rect 3760 3100 3920 3110
rect 4080 3100 4200 3110
rect 4480 3100 4520 3110
rect 4840 3100 4920 3110
rect 5880 3100 6120 3110
rect 6600 3100 6640 3110
rect 9080 3100 9120 3110
rect 9200 3100 9240 3110
rect 9440 3100 9520 3110
rect 1240 3090 1320 3100
rect 2000 3090 2040 3100
rect 3760 3090 3880 3100
rect 4000 3090 4040 3100
rect 4120 3090 4240 3100
rect 4520 3090 4600 3100
rect 4760 3090 4880 3100
rect 6600 3090 6640 3100
rect 9040 3090 9120 3100
rect 9200 3090 9240 3100
rect 9360 3090 9480 3100
rect 1240 3080 1320 3090
rect 2000 3080 2040 3090
rect 3760 3080 3880 3090
rect 4000 3080 4040 3090
rect 4120 3080 4240 3090
rect 4520 3080 4600 3090
rect 4760 3080 4880 3090
rect 6600 3080 6640 3090
rect 9040 3080 9120 3090
rect 9200 3080 9240 3090
rect 9360 3080 9480 3090
rect 1240 3070 1320 3080
rect 2000 3070 2040 3080
rect 3760 3070 3880 3080
rect 4000 3070 4040 3080
rect 4120 3070 4240 3080
rect 4520 3070 4600 3080
rect 4760 3070 4880 3080
rect 6600 3070 6640 3080
rect 9040 3070 9120 3080
rect 9200 3070 9240 3080
rect 9360 3070 9480 3080
rect 1240 3060 1320 3070
rect 2000 3060 2040 3070
rect 3760 3060 3880 3070
rect 4000 3060 4040 3070
rect 4120 3060 4240 3070
rect 4520 3060 4600 3070
rect 4760 3060 4880 3070
rect 6600 3060 6640 3070
rect 9040 3060 9120 3070
rect 9200 3060 9240 3070
rect 9360 3060 9480 3070
rect 1200 3050 1320 3060
rect 3160 3050 3200 3060
rect 3720 3050 3760 3060
rect 4120 3050 4160 3060
rect 4200 3050 4280 3060
rect 4560 3050 4640 3060
rect 4720 3050 4840 3060
rect 6600 3050 6640 3060
rect 8320 3050 8360 3060
rect 9040 3050 9080 3060
rect 9240 3050 9480 3060
rect 1200 3040 1320 3050
rect 3160 3040 3200 3050
rect 3720 3040 3760 3050
rect 4120 3040 4160 3050
rect 4200 3040 4280 3050
rect 4560 3040 4640 3050
rect 4720 3040 4840 3050
rect 6600 3040 6640 3050
rect 8320 3040 8360 3050
rect 9040 3040 9080 3050
rect 9240 3040 9480 3050
rect 1200 3030 1320 3040
rect 3160 3030 3200 3040
rect 3720 3030 3760 3040
rect 4120 3030 4160 3040
rect 4200 3030 4280 3040
rect 4560 3030 4640 3040
rect 4720 3030 4840 3040
rect 6600 3030 6640 3040
rect 8320 3030 8360 3040
rect 9040 3030 9080 3040
rect 9240 3030 9480 3040
rect 1200 3020 1320 3030
rect 3160 3020 3200 3030
rect 3720 3020 3760 3030
rect 4120 3020 4160 3030
rect 4200 3020 4280 3030
rect 4560 3020 4640 3030
rect 4720 3020 4840 3030
rect 6600 3020 6640 3030
rect 8320 3020 8360 3030
rect 9040 3020 9080 3030
rect 9240 3020 9480 3030
rect 1200 3010 1320 3020
rect 3160 3010 3200 3020
rect 3720 3010 3880 3020
rect 4040 3010 4120 3020
rect 4160 3010 4320 3020
rect 4680 3010 4760 3020
rect 5200 3010 5240 3020
rect 6520 3010 6560 3020
rect 8400 3010 8440 3020
rect 9040 3010 9080 3020
rect 9120 3010 9400 3020
rect 1200 3000 1320 3010
rect 3160 3000 3200 3010
rect 3720 3000 3880 3010
rect 4040 3000 4120 3010
rect 4160 3000 4320 3010
rect 4680 3000 4760 3010
rect 5200 3000 5240 3010
rect 6520 3000 6560 3010
rect 8400 3000 8440 3010
rect 9040 3000 9080 3010
rect 9120 3000 9400 3010
rect 1200 2990 1320 3000
rect 3160 2990 3200 3000
rect 3720 2990 3880 3000
rect 4040 2990 4120 3000
rect 4160 2990 4320 3000
rect 4680 2990 4760 3000
rect 5200 2990 5240 3000
rect 6520 2990 6560 3000
rect 8400 2990 8440 3000
rect 9040 2990 9080 3000
rect 9120 2990 9400 3000
rect 1200 2980 1320 2990
rect 3160 2980 3200 2990
rect 3720 2980 3880 2990
rect 4040 2980 4120 2990
rect 4160 2980 4320 2990
rect 4680 2980 4760 2990
rect 5200 2980 5240 2990
rect 6520 2980 6560 2990
rect 8400 2980 8440 2990
rect 9040 2980 9080 2990
rect 9120 2980 9400 2990
rect 1160 2970 1280 2980
rect 3160 2970 3200 2980
rect 3840 2970 3880 2980
rect 4240 2970 4360 2980
rect 6520 2970 6600 2980
rect 8960 2970 9120 2980
rect 9200 2970 9280 2980
rect 1160 2960 1280 2970
rect 3160 2960 3200 2970
rect 3840 2960 3880 2970
rect 4240 2960 4360 2970
rect 6520 2960 6600 2970
rect 8960 2960 9120 2970
rect 9200 2960 9280 2970
rect 1160 2950 1280 2960
rect 3160 2950 3200 2960
rect 3840 2950 3880 2960
rect 4240 2950 4360 2960
rect 6520 2950 6600 2960
rect 8960 2950 9120 2960
rect 9200 2950 9280 2960
rect 1160 2940 1280 2950
rect 3160 2940 3200 2950
rect 3840 2940 3880 2950
rect 4240 2940 4360 2950
rect 6520 2940 6600 2950
rect 8960 2940 9120 2950
rect 9200 2940 9280 2950
rect 1160 2930 1280 2940
rect 3800 2930 3880 2940
rect 3960 2930 4000 2940
rect 4280 2930 4400 2940
rect 5160 2930 5200 2940
rect 6520 2930 6600 2940
rect 8960 2930 9120 2940
rect 9200 2930 9240 2940
rect 9360 2930 9400 2940
rect 1160 2920 1280 2930
rect 3800 2920 3880 2930
rect 3960 2920 4000 2930
rect 4280 2920 4400 2930
rect 5160 2920 5200 2930
rect 6520 2920 6600 2930
rect 8960 2920 9120 2930
rect 9200 2920 9240 2930
rect 9360 2920 9400 2930
rect 1160 2910 1280 2920
rect 3800 2910 3880 2920
rect 3960 2910 4000 2920
rect 4280 2910 4400 2920
rect 5160 2910 5200 2920
rect 6520 2910 6600 2920
rect 8960 2910 9120 2920
rect 9200 2910 9240 2920
rect 9360 2910 9400 2920
rect 1160 2900 1280 2910
rect 3800 2900 3880 2910
rect 3960 2900 4000 2910
rect 4280 2900 4400 2910
rect 5160 2900 5200 2910
rect 6520 2900 6600 2910
rect 8960 2900 9120 2910
rect 9200 2900 9240 2910
rect 9360 2900 9400 2910
rect 1160 2890 1240 2900
rect 3880 2890 3920 2900
rect 3960 2890 4000 2900
rect 4240 2890 4280 2900
rect 4360 2890 4440 2900
rect 6520 2890 6600 2900
rect 7480 2890 7520 2900
rect 9000 2890 9080 2900
rect 1160 2880 1240 2890
rect 3880 2880 3920 2890
rect 3960 2880 4000 2890
rect 4240 2880 4280 2890
rect 4360 2880 4440 2890
rect 6520 2880 6600 2890
rect 7480 2880 7520 2890
rect 9000 2880 9080 2890
rect 1160 2870 1240 2880
rect 3880 2870 3920 2880
rect 3960 2870 4000 2880
rect 4240 2870 4280 2880
rect 4360 2870 4440 2880
rect 6520 2870 6600 2880
rect 7480 2870 7520 2880
rect 9000 2870 9080 2880
rect 1160 2860 1240 2870
rect 3880 2860 3920 2870
rect 3960 2860 4000 2870
rect 4240 2860 4280 2870
rect 4360 2860 4440 2870
rect 6520 2860 6600 2870
rect 7480 2860 7520 2870
rect 9000 2860 9080 2870
rect 1120 2850 1240 2860
rect 1960 2850 2000 2860
rect 3880 2850 3960 2860
rect 4440 2850 4520 2860
rect 4640 2850 4680 2860
rect 5120 2850 5160 2860
rect 6520 2850 6560 2860
rect 8960 2850 9040 2860
rect 1120 2840 1240 2850
rect 1960 2840 2000 2850
rect 3880 2840 3960 2850
rect 4440 2840 4520 2850
rect 4640 2840 4680 2850
rect 5120 2840 5160 2850
rect 6520 2840 6560 2850
rect 8960 2840 9040 2850
rect 1120 2830 1240 2840
rect 1960 2830 2000 2840
rect 3880 2830 3960 2840
rect 4440 2830 4520 2840
rect 4640 2830 4680 2840
rect 5120 2830 5160 2840
rect 6520 2830 6560 2840
rect 8960 2830 9040 2840
rect 1120 2820 1240 2830
rect 1960 2820 2000 2830
rect 3880 2820 3960 2830
rect 4440 2820 4520 2830
rect 4640 2820 4680 2830
rect 5120 2820 5160 2830
rect 6520 2820 6560 2830
rect 8960 2820 9040 2830
rect 1120 2810 1240 2820
rect 1960 2810 2000 2820
rect 4480 2810 4760 2820
rect 5080 2810 5200 2820
rect 5720 2810 6120 2820
rect 6520 2810 6560 2820
rect 7120 2810 7160 2820
rect 8160 2810 8200 2820
rect 8880 2810 9000 2820
rect 1120 2800 1240 2810
rect 1960 2800 2000 2810
rect 4480 2800 4760 2810
rect 5080 2800 5200 2810
rect 5720 2800 6120 2810
rect 6520 2800 6560 2810
rect 7120 2800 7160 2810
rect 8160 2800 8200 2810
rect 8880 2800 9000 2810
rect 1120 2790 1240 2800
rect 1960 2790 2000 2800
rect 4480 2790 4760 2800
rect 5080 2790 5200 2800
rect 5720 2790 6120 2800
rect 6520 2790 6560 2800
rect 7120 2790 7160 2800
rect 8160 2790 8200 2800
rect 8880 2790 9000 2800
rect 1120 2780 1240 2790
rect 1960 2780 2000 2790
rect 4480 2780 4760 2790
rect 5080 2780 5200 2790
rect 5720 2780 6120 2790
rect 6520 2780 6560 2790
rect 7120 2780 7160 2790
rect 8160 2780 8200 2790
rect 8880 2780 9000 2790
rect 1080 2770 1200 2780
rect 1960 2770 2000 2780
rect 3880 2770 3920 2780
rect 4560 2770 4840 2780
rect 4920 2770 5040 2780
rect 5120 2770 5200 2780
rect 5520 2770 6040 2780
rect 6120 2770 6160 2780
rect 6520 2770 6560 2780
rect 8120 2770 8160 2780
rect 8720 2770 8760 2780
rect 8800 2770 8920 2780
rect 1080 2760 1200 2770
rect 1960 2760 2000 2770
rect 3880 2760 3920 2770
rect 4560 2760 4840 2770
rect 4920 2760 5040 2770
rect 5120 2760 5200 2770
rect 5520 2760 6040 2770
rect 6120 2760 6160 2770
rect 6520 2760 6560 2770
rect 8120 2760 8160 2770
rect 8720 2760 8760 2770
rect 8800 2760 8920 2770
rect 1080 2750 1200 2760
rect 1960 2750 2000 2760
rect 3880 2750 3920 2760
rect 4560 2750 4840 2760
rect 4920 2750 5040 2760
rect 5120 2750 5200 2760
rect 5520 2750 6040 2760
rect 6120 2750 6160 2760
rect 6520 2750 6560 2760
rect 8120 2750 8160 2760
rect 8720 2750 8760 2760
rect 8800 2750 8920 2760
rect 1080 2740 1200 2750
rect 1960 2740 2000 2750
rect 3880 2740 3920 2750
rect 4560 2740 4840 2750
rect 4920 2740 5040 2750
rect 5120 2740 5200 2750
rect 5520 2740 6040 2750
rect 6120 2740 6160 2750
rect 6520 2740 6560 2750
rect 8120 2740 8160 2750
rect 8720 2740 8760 2750
rect 8800 2740 8920 2750
rect 1080 2730 1160 2740
rect 1960 2730 2000 2740
rect 3880 2730 3920 2740
rect 4680 2730 5000 2740
rect 5120 2730 5200 2740
rect 5240 2730 5360 2740
rect 5480 2730 5960 2740
rect 6520 2730 6560 2740
rect 8680 2730 8840 2740
rect 8880 2730 8920 2740
rect 9960 2730 9990 2740
rect 1080 2720 1160 2730
rect 1960 2720 2000 2730
rect 3880 2720 3920 2730
rect 4680 2720 5000 2730
rect 5120 2720 5200 2730
rect 5240 2720 5360 2730
rect 5480 2720 5960 2730
rect 6520 2720 6560 2730
rect 8680 2720 8840 2730
rect 8880 2720 8920 2730
rect 9960 2720 9990 2730
rect 1080 2710 1160 2720
rect 1960 2710 2000 2720
rect 3880 2710 3920 2720
rect 4680 2710 5000 2720
rect 5120 2710 5200 2720
rect 5240 2710 5360 2720
rect 5480 2710 5960 2720
rect 6520 2710 6560 2720
rect 8680 2710 8840 2720
rect 8880 2710 8920 2720
rect 9960 2710 9990 2720
rect 1080 2700 1160 2710
rect 1960 2700 2000 2710
rect 3880 2700 3920 2710
rect 4680 2700 5000 2710
rect 5120 2700 5200 2710
rect 5240 2700 5360 2710
rect 5480 2700 5960 2710
rect 6520 2700 6560 2710
rect 8680 2700 8840 2710
rect 8880 2700 8920 2710
rect 9960 2700 9990 2710
rect 1040 2690 1120 2700
rect 1960 2690 2000 2700
rect 4840 2690 5000 2700
rect 5120 2690 5160 2700
rect 5200 2690 5400 2700
rect 5440 2690 5880 2700
rect 6520 2690 6560 2700
rect 7680 2690 7720 2700
rect 9000 2690 9080 2700
rect 9160 2690 9240 2700
rect 1040 2680 1120 2690
rect 1960 2680 2000 2690
rect 4840 2680 5000 2690
rect 5120 2680 5160 2690
rect 5200 2680 5400 2690
rect 5440 2680 5880 2690
rect 6520 2680 6560 2690
rect 7680 2680 7720 2690
rect 9000 2680 9080 2690
rect 9160 2680 9240 2690
rect 1040 2670 1120 2680
rect 1960 2670 2000 2680
rect 4840 2670 5000 2680
rect 5120 2670 5160 2680
rect 5200 2670 5400 2680
rect 5440 2670 5880 2680
rect 6520 2670 6560 2680
rect 7680 2670 7720 2680
rect 9000 2670 9080 2680
rect 9160 2670 9240 2680
rect 1040 2660 1120 2670
rect 1960 2660 2000 2670
rect 4840 2660 5000 2670
rect 5120 2660 5160 2670
rect 5200 2660 5400 2670
rect 5440 2660 5880 2670
rect 6520 2660 6560 2670
rect 7680 2660 7720 2670
rect 9000 2660 9080 2670
rect 9160 2660 9240 2670
rect 1040 2650 1120 2660
rect 2280 2650 2400 2660
rect 2880 2650 2920 2660
rect 3080 2650 3160 2660
rect 4800 2650 4960 2660
rect 5080 2650 5360 2660
rect 5400 2650 5840 2660
rect 6200 2650 6240 2660
rect 9040 2650 9120 2660
rect 9160 2650 9200 2660
rect 1040 2640 1120 2650
rect 2280 2640 2400 2650
rect 2880 2640 2920 2650
rect 3080 2640 3160 2650
rect 4800 2640 4960 2650
rect 5080 2640 5360 2650
rect 5400 2640 5840 2650
rect 6200 2640 6240 2650
rect 9040 2640 9120 2650
rect 9160 2640 9200 2650
rect 1040 2630 1120 2640
rect 2280 2630 2400 2640
rect 2880 2630 2920 2640
rect 3080 2630 3160 2640
rect 4800 2630 4960 2640
rect 5080 2630 5360 2640
rect 5400 2630 5840 2640
rect 6200 2630 6240 2640
rect 9040 2630 9120 2640
rect 9160 2630 9200 2640
rect 1040 2620 1120 2630
rect 2280 2620 2400 2630
rect 2880 2620 2920 2630
rect 3080 2620 3160 2630
rect 4800 2620 4960 2630
rect 5080 2620 5360 2630
rect 5400 2620 5840 2630
rect 6200 2620 6240 2630
rect 9040 2620 9120 2630
rect 9160 2620 9200 2630
rect 1000 2610 1080 2620
rect 1920 2610 1960 2620
rect 2080 2610 2280 2620
rect 2360 2610 2400 2620
rect 2840 2610 2880 2620
rect 3040 2610 3120 2620
rect 3880 2610 3920 2620
rect 4720 2610 5800 2620
rect 6240 2610 6280 2620
rect 9040 2610 9160 2620
rect 9920 2610 9990 2620
rect 1000 2600 1080 2610
rect 1920 2600 1960 2610
rect 2080 2600 2280 2610
rect 2360 2600 2400 2610
rect 2840 2600 2880 2610
rect 3040 2600 3120 2610
rect 3880 2600 3920 2610
rect 4720 2600 5800 2610
rect 6240 2600 6280 2610
rect 9040 2600 9160 2610
rect 9920 2600 9990 2610
rect 1000 2590 1080 2600
rect 1920 2590 1960 2600
rect 2080 2590 2280 2600
rect 2360 2590 2400 2600
rect 2840 2590 2880 2600
rect 3040 2590 3120 2600
rect 3880 2590 3920 2600
rect 4720 2590 5800 2600
rect 6240 2590 6280 2600
rect 9040 2590 9160 2600
rect 9920 2590 9990 2600
rect 1000 2580 1080 2590
rect 1920 2580 1960 2590
rect 2080 2580 2280 2590
rect 2360 2580 2400 2590
rect 2840 2580 2880 2590
rect 3040 2580 3120 2590
rect 3880 2580 3920 2590
rect 4720 2580 5800 2590
rect 6240 2580 6280 2590
rect 9040 2580 9160 2590
rect 9920 2580 9990 2590
rect 1000 2570 1080 2580
rect 2320 2570 2360 2580
rect 2880 2570 2920 2580
rect 3880 2570 3920 2580
rect 4240 2570 4280 2580
rect 4520 2570 4800 2580
rect 4840 2570 4880 2580
rect 4920 2570 5760 2580
rect 9040 2570 9160 2580
rect 1000 2560 1080 2570
rect 2320 2560 2360 2570
rect 2880 2560 2920 2570
rect 3880 2560 3920 2570
rect 4240 2560 4280 2570
rect 4520 2560 4800 2570
rect 4840 2560 4880 2570
rect 4920 2560 5760 2570
rect 9040 2560 9160 2570
rect 1000 2550 1080 2560
rect 2320 2550 2360 2560
rect 2880 2550 2920 2560
rect 3880 2550 3920 2560
rect 4240 2550 4280 2560
rect 4520 2550 4800 2560
rect 4840 2550 4880 2560
rect 4920 2550 5760 2560
rect 9040 2550 9160 2560
rect 1000 2540 1080 2550
rect 2320 2540 2360 2550
rect 2880 2540 2920 2550
rect 3880 2540 3920 2550
rect 4240 2540 4280 2550
rect 4520 2540 4800 2550
rect 4840 2540 4880 2550
rect 4920 2540 5760 2550
rect 9040 2540 9160 2550
rect 960 2530 1040 2540
rect 3920 2530 3960 2540
rect 4680 2530 5760 2540
rect 6280 2530 6320 2540
rect 6760 2530 6800 2540
rect 9080 2530 9120 2540
rect 960 2520 1040 2530
rect 3920 2520 3960 2530
rect 4680 2520 5760 2530
rect 6280 2520 6320 2530
rect 6760 2520 6800 2530
rect 9080 2520 9120 2530
rect 960 2510 1040 2520
rect 3920 2510 3960 2520
rect 4680 2510 5760 2520
rect 6280 2510 6320 2520
rect 6760 2510 6800 2520
rect 9080 2510 9120 2520
rect 960 2500 1040 2510
rect 3920 2500 3960 2510
rect 4680 2500 5760 2510
rect 6280 2500 6320 2510
rect 6760 2500 6800 2510
rect 9080 2500 9120 2510
rect 960 2490 1040 2500
rect 1880 2490 1920 2500
rect 3960 2490 4120 2500
rect 4600 2490 5600 2500
rect 5640 2490 5760 2500
rect 6320 2490 6360 2500
rect 7280 2490 7320 2500
rect 9320 2490 9600 2500
rect 960 2480 1040 2490
rect 1880 2480 1920 2490
rect 3960 2480 4120 2490
rect 4600 2480 5600 2490
rect 5640 2480 5760 2490
rect 6320 2480 6360 2490
rect 7280 2480 7320 2490
rect 9320 2480 9600 2490
rect 960 2470 1040 2480
rect 1880 2470 1920 2480
rect 3960 2470 4120 2480
rect 4600 2470 5600 2480
rect 5640 2470 5760 2480
rect 6320 2470 6360 2480
rect 7280 2470 7320 2480
rect 9320 2470 9600 2480
rect 960 2460 1040 2470
rect 1880 2460 1920 2470
rect 3960 2460 4120 2470
rect 4600 2460 5600 2470
rect 5640 2460 5760 2470
rect 6320 2460 6360 2470
rect 7280 2460 7320 2470
rect 9320 2460 9600 2470
rect 920 2450 1040 2460
rect 1880 2450 1920 2460
rect 3240 2450 3280 2460
rect 3960 2450 4080 2460
rect 4560 2450 5560 2460
rect 5640 2450 5720 2460
rect 6720 2450 6760 2460
rect 7320 2450 7360 2460
rect 9400 2450 9480 2460
rect 9560 2450 9640 2460
rect 920 2440 1040 2450
rect 1880 2440 1920 2450
rect 3240 2440 3280 2450
rect 3960 2440 4080 2450
rect 4560 2440 5560 2450
rect 5640 2440 5720 2450
rect 6720 2440 6760 2450
rect 7320 2440 7360 2450
rect 9400 2440 9480 2450
rect 9560 2440 9640 2450
rect 920 2430 1040 2440
rect 1880 2430 1920 2440
rect 3240 2430 3280 2440
rect 3960 2430 4080 2440
rect 4560 2430 5560 2440
rect 5640 2430 5720 2440
rect 6720 2430 6760 2440
rect 7320 2430 7360 2440
rect 9400 2430 9480 2440
rect 9560 2430 9640 2440
rect 920 2420 1040 2430
rect 1880 2420 1920 2430
rect 3240 2420 3280 2430
rect 3960 2420 4080 2430
rect 4560 2420 5560 2430
rect 5640 2420 5720 2430
rect 6720 2420 6760 2430
rect 7320 2420 7360 2430
rect 9400 2420 9480 2430
rect 9560 2420 9640 2430
rect 920 2410 1040 2420
rect 4560 2410 5560 2420
rect 5600 2410 5680 2420
rect 6360 2410 6400 2420
rect 6720 2410 6760 2420
rect 920 2400 1040 2410
rect 4560 2400 5560 2410
rect 5600 2400 5680 2410
rect 6360 2400 6400 2410
rect 6720 2400 6760 2410
rect 920 2390 1040 2400
rect 4560 2390 5560 2400
rect 5600 2390 5680 2400
rect 6360 2390 6400 2400
rect 6720 2390 6760 2400
rect 920 2380 1040 2390
rect 4560 2380 5560 2390
rect 5600 2380 5680 2390
rect 6360 2380 6400 2390
rect 6720 2380 6760 2390
rect 880 2370 1000 2380
rect 3280 2370 3320 2380
rect 4520 2370 5680 2380
rect 9680 2370 9760 2380
rect 880 2360 1000 2370
rect 3280 2360 3320 2370
rect 4520 2360 5680 2370
rect 9680 2360 9760 2370
rect 880 2350 1000 2360
rect 3280 2350 3320 2360
rect 4520 2350 5680 2360
rect 9680 2350 9760 2360
rect 880 2340 1000 2350
rect 3280 2340 3320 2350
rect 4520 2340 5680 2350
rect 9680 2340 9760 2350
rect 880 2330 1000 2340
rect 1840 2330 1880 2340
rect 3280 2330 3320 2340
rect 4480 2330 5640 2340
rect 6400 2330 6440 2340
rect 6840 2330 6920 2340
rect 8440 2330 8520 2340
rect 9240 2330 9280 2340
rect 9320 2330 9400 2340
rect 9600 2330 9760 2340
rect 880 2320 1000 2330
rect 1840 2320 1880 2330
rect 3280 2320 3320 2330
rect 4480 2320 5640 2330
rect 6400 2320 6440 2330
rect 6840 2320 6920 2330
rect 8440 2320 8520 2330
rect 9240 2320 9280 2330
rect 9320 2320 9400 2330
rect 9600 2320 9760 2330
rect 880 2310 1000 2320
rect 1840 2310 1880 2320
rect 3280 2310 3320 2320
rect 4480 2310 5640 2320
rect 6400 2310 6440 2320
rect 6840 2310 6920 2320
rect 8440 2310 8520 2320
rect 9240 2310 9280 2320
rect 9320 2310 9400 2320
rect 9600 2310 9760 2320
rect 880 2300 1000 2310
rect 1840 2300 1880 2310
rect 3280 2300 3320 2310
rect 4480 2300 5640 2310
rect 6400 2300 6440 2310
rect 6840 2300 6920 2310
rect 8440 2300 8520 2310
rect 9240 2300 9280 2310
rect 9320 2300 9400 2310
rect 9600 2300 9760 2310
rect 840 2290 1000 2300
rect 1840 2290 1880 2300
rect 4080 2290 5440 2300
rect 5520 2290 5640 2300
rect 6840 2290 6960 2300
rect 7080 2290 7120 2300
rect 9200 2290 9480 2300
rect 9600 2290 9640 2300
rect 9720 2290 9760 2300
rect 840 2280 1000 2290
rect 1840 2280 1880 2290
rect 4080 2280 5440 2290
rect 5520 2280 5640 2290
rect 6840 2280 6960 2290
rect 7080 2280 7120 2290
rect 9200 2280 9480 2290
rect 9600 2280 9640 2290
rect 9720 2280 9760 2290
rect 840 2270 1000 2280
rect 1840 2270 1880 2280
rect 4080 2270 5440 2280
rect 5520 2270 5640 2280
rect 6840 2270 6960 2280
rect 7080 2270 7120 2280
rect 9200 2270 9480 2280
rect 9600 2270 9640 2280
rect 9720 2270 9760 2280
rect 840 2260 1000 2270
rect 1840 2260 1880 2270
rect 4080 2260 5440 2270
rect 5520 2260 5640 2270
rect 6840 2260 6960 2270
rect 7080 2260 7120 2270
rect 9200 2260 9480 2270
rect 9600 2260 9640 2270
rect 9720 2260 9760 2270
rect 840 2250 1000 2260
rect 3320 2250 3360 2260
rect 4320 2250 5400 2260
rect 5520 2250 5600 2260
rect 6720 2250 6760 2260
rect 6840 2250 7160 2260
rect 7200 2250 7280 2260
rect 8600 2250 8640 2260
rect 9120 2250 9160 2260
rect 9360 2250 9640 2260
rect 9680 2250 9760 2260
rect 840 2240 1000 2250
rect 3320 2240 3360 2250
rect 4320 2240 5400 2250
rect 5520 2240 5600 2250
rect 6720 2240 6760 2250
rect 6840 2240 7160 2250
rect 7200 2240 7280 2250
rect 8600 2240 8640 2250
rect 9120 2240 9160 2250
rect 9360 2240 9640 2250
rect 9680 2240 9760 2250
rect 840 2230 1000 2240
rect 3320 2230 3360 2240
rect 4320 2230 5400 2240
rect 5520 2230 5600 2240
rect 6720 2230 6760 2240
rect 6840 2230 7160 2240
rect 7200 2230 7280 2240
rect 8600 2230 8640 2240
rect 9120 2230 9160 2240
rect 9360 2230 9640 2240
rect 9680 2230 9760 2240
rect 840 2220 1000 2230
rect 3320 2220 3360 2230
rect 4320 2220 5400 2230
rect 5520 2220 5600 2230
rect 6720 2220 6760 2230
rect 6840 2220 7160 2230
rect 7200 2220 7280 2230
rect 8600 2220 8640 2230
rect 9120 2220 9160 2230
rect 9360 2220 9640 2230
rect 9680 2220 9760 2230
rect 800 2210 1000 2220
rect 3320 2210 3360 2220
rect 4360 2210 5360 2220
rect 6720 2210 6760 2220
rect 6920 2210 7000 2220
rect 7280 2210 7360 2220
rect 9480 2210 9760 2220
rect 800 2200 1000 2210
rect 3320 2200 3360 2210
rect 4360 2200 5360 2210
rect 6720 2200 6760 2210
rect 6920 2200 7000 2210
rect 7280 2200 7360 2210
rect 9480 2200 9760 2210
rect 800 2190 1000 2200
rect 3320 2190 3360 2200
rect 4360 2190 5360 2200
rect 6720 2190 6760 2200
rect 6920 2190 7000 2200
rect 7280 2190 7360 2200
rect 9480 2190 9760 2200
rect 800 2180 1000 2190
rect 3320 2180 3360 2190
rect 4360 2180 5360 2190
rect 6720 2180 6760 2190
rect 6920 2180 7000 2190
rect 7280 2180 7360 2190
rect 9480 2180 9760 2190
rect 800 2170 1000 2180
rect 2440 2170 2520 2180
rect 2640 2170 2680 2180
rect 3320 2170 3360 2180
rect 4360 2170 5320 2180
rect 6480 2170 6520 2180
rect 6720 2170 6760 2180
rect 6960 2170 7080 2180
rect 7280 2170 7320 2180
rect 7360 2170 7400 2180
rect 7480 2170 7520 2180
rect 7680 2170 7720 2180
rect 9600 2170 9680 2180
rect 800 2160 1000 2170
rect 2440 2160 2520 2170
rect 2640 2160 2680 2170
rect 3320 2160 3360 2170
rect 4360 2160 5320 2170
rect 6480 2160 6520 2170
rect 6720 2160 6760 2170
rect 6960 2160 7080 2170
rect 7280 2160 7320 2170
rect 7360 2160 7400 2170
rect 7480 2160 7520 2170
rect 7680 2160 7720 2170
rect 9600 2160 9680 2170
rect 800 2150 1000 2160
rect 2440 2150 2520 2160
rect 2640 2150 2680 2160
rect 3320 2150 3360 2160
rect 4360 2150 5320 2160
rect 6480 2150 6520 2160
rect 6720 2150 6760 2160
rect 6960 2150 7080 2160
rect 7280 2150 7320 2160
rect 7360 2150 7400 2160
rect 7480 2150 7520 2160
rect 7680 2150 7720 2160
rect 9600 2150 9680 2160
rect 800 2140 1000 2150
rect 2440 2140 2520 2150
rect 2640 2140 2680 2150
rect 3320 2140 3360 2150
rect 4360 2140 5320 2150
rect 6480 2140 6520 2150
rect 6720 2140 6760 2150
rect 6960 2140 7080 2150
rect 7280 2140 7320 2150
rect 7360 2140 7400 2150
rect 7480 2140 7520 2150
rect 7680 2140 7720 2150
rect 9600 2140 9680 2150
rect 760 2130 960 2140
rect 3320 2130 3360 2140
rect 4360 2130 5280 2140
rect 6720 2130 6760 2140
rect 7000 2130 7280 2140
rect 7400 2130 7480 2140
rect 7720 2130 7840 2140
rect 9200 2130 9240 2140
rect 760 2120 960 2130
rect 3320 2120 3360 2130
rect 4360 2120 5280 2130
rect 6720 2120 6760 2130
rect 7000 2120 7280 2130
rect 7400 2120 7480 2130
rect 7720 2120 7840 2130
rect 9200 2120 9240 2130
rect 760 2110 960 2120
rect 3320 2110 3360 2120
rect 4360 2110 5280 2120
rect 6720 2110 6760 2120
rect 7000 2110 7280 2120
rect 7400 2110 7480 2120
rect 7720 2110 7840 2120
rect 9200 2110 9240 2120
rect 760 2100 960 2110
rect 3320 2100 3360 2110
rect 4360 2100 5280 2110
rect 6720 2100 6760 2110
rect 7000 2100 7280 2110
rect 7400 2100 7480 2110
rect 7720 2100 7840 2110
rect 9200 2100 9240 2110
rect 760 2090 960 2100
rect 3320 2090 3360 2100
rect 4320 2090 5280 2100
rect 6520 2090 6560 2100
rect 7080 2090 7240 2100
rect 7840 2090 7880 2100
rect 8440 2090 8480 2100
rect 9520 2090 9600 2100
rect 9640 2090 9680 2100
rect 760 2080 960 2090
rect 3320 2080 3360 2090
rect 4320 2080 5280 2090
rect 6520 2080 6560 2090
rect 7080 2080 7240 2090
rect 7840 2080 7880 2090
rect 8440 2080 8480 2090
rect 9520 2080 9600 2090
rect 9640 2080 9680 2090
rect 760 2070 960 2080
rect 3320 2070 3360 2080
rect 4320 2070 5280 2080
rect 6520 2070 6560 2080
rect 7080 2070 7240 2080
rect 7840 2070 7880 2080
rect 8440 2070 8480 2080
rect 9520 2070 9600 2080
rect 9640 2070 9680 2080
rect 760 2060 960 2070
rect 3320 2060 3360 2070
rect 4320 2060 5280 2070
rect 6520 2060 6560 2070
rect 7080 2060 7240 2070
rect 7840 2060 7880 2070
rect 8440 2060 8480 2070
rect 9520 2060 9600 2070
rect 9640 2060 9680 2070
rect 720 2050 960 2060
rect 3320 2050 3360 2060
rect 4360 2050 5120 2060
rect 5160 2050 5240 2060
rect 6520 2050 6560 2060
rect 7320 2050 7360 2060
rect 7720 2050 7800 2060
rect 7840 2050 7880 2060
rect 8520 2050 8560 2060
rect 9080 2050 9120 2060
rect 9240 2050 9280 2060
rect 9360 2050 9400 2060
rect 9440 2050 9480 2060
rect 720 2040 960 2050
rect 3320 2040 3360 2050
rect 4360 2040 5120 2050
rect 5160 2040 5240 2050
rect 6520 2040 6560 2050
rect 7320 2040 7360 2050
rect 7720 2040 7800 2050
rect 7840 2040 7880 2050
rect 8520 2040 8560 2050
rect 9080 2040 9120 2050
rect 9240 2040 9280 2050
rect 9360 2040 9400 2050
rect 9440 2040 9480 2050
rect 720 2030 960 2040
rect 3320 2030 3360 2040
rect 4360 2030 5120 2040
rect 5160 2030 5240 2040
rect 6520 2030 6560 2040
rect 7320 2030 7360 2040
rect 7720 2030 7800 2040
rect 7840 2030 7880 2040
rect 8520 2030 8560 2040
rect 9080 2030 9120 2040
rect 9240 2030 9280 2040
rect 9360 2030 9400 2040
rect 9440 2030 9480 2040
rect 720 2020 960 2030
rect 3320 2020 3360 2030
rect 4360 2020 5120 2030
rect 5160 2020 5240 2030
rect 6520 2020 6560 2030
rect 7320 2020 7360 2030
rect 7720 2020 7800 2030
rect 7840 2020 7880 2030
rect 8520 2020 8560 2030
rect 9080 2020 9120 2030
rect 9240 2020 9280 2030
rect 9360 2020 9400 2030
rect 9440 2020 9480 2030
rect 720 2010 960 2020
rect 3320 2010 3360 2020
rect 4320 2010 5120 2020
rect 6520 2010 6560 2020
rect 6760 2010 6800 2020
rect 7720 2010 7960 2020
rect 8600 2010 8680 2020
rect 720 2000 960 2010
rect 3320 2000 3360 2010
rect 4320 2000 5120 2010
rect 6520 2000 6560 2010
rect 6760 2000 6800 2010
rect 7720 2000 7960 2010
rect 8600 2000 8680 2010
rect 720 1990 960 2000
rect 3320 1990 3360 2000
rect 4320 1990 5120 2000
rect 6520 1990 6560 2000
rect 6760 1990 6800 2000
rect 7720 1990 7960 2000
rect 8600 1990 8680 2000
rect 720 1980 960 1990
rect 3320 1980 3360 1990
rect 4320 1980 5120 1990
rect 6520 1980 6560 1990
rect 6760 1980 6800 1990
rect 7720 1980 7960 1990
rect 8600 1980 8680 1990
rect 680 1970 960 1980
rect 3320 1970 3360 1980
rect 4360 1970 5040 1980
rect 6200 1970 6280 1980
rect 6520 1970 6560 1980
rect 6760 1970 6800 1980
rect 7720 1970 7760 1980
rect 7880 1970 7960 1980
rect 8760 1970 8800 1980
rect 680 1960 960 1970
rect 3320 1960 3360 1970
rect 4360 1960 5040 1970
rect 6200 1960 6280 1970
rect 6520 1960 6560 1970
rect 6760 1960 6800 1970
rect 7720 1960 7760 1970
rect 7880 1960 7960 1970
rect 8760 1960 8800 1970
rect 680 1950 960 1960
rect 3320 1950 3360 1960
rect 4360 1950 5040 1960
rect 6200 1950 6280 1960
rect 6520 1950 6560 1960
rect 6760 1950 6800 1960
rect 7720 1950 7760 1960
rect 7880 1950 7960 1960
rect 8760 1950 8800 1960
rect 680 1940 960 1950
rect 3320 1940 3360 1950
rect 4360 1940 5040 1950
rect 6200 1940 6280 1950
rect 6520 1940 6560 1950
rect 6760 1940 6800 1950
rect 7720 1940 7760 1950
rect 7880 1940 7960 1950
rect 8760 1940 8800 1950
rect 680 1930 920 1940
rect 3320 1930 3360 1940
rect 4360 1930 4480 1940
rect 4640 1930 4760 1940
rect 4880 1930 4960 1940
rect 6200 1930 6320 1940
rect 6520 1930 6560 1940
rect 6760 1930 6800 1940
rect 7720 1930 7760 1940
rect 680 1920 920 1930
rect 3320 1920 3360 1930
rect 4360 1920 4480 1930
rect 4640 1920 4760 1930
rect 4880 1920 4960 1930
rect 6200 1920 6320 1930
rect 6520 1920 6560 1930
rect 6760 1920 6800 1930
rect 7720 1920 7760 1930
rect 680 1910 920 1920
rect 3320 1910 3360 1920
rect 4360 1910 4480 1920
rect 4640 1910 4760 1920
rect 4880 1910 4960 1920
rect 6200 1910 6320 1920
rect 6520 1910 6560 1920
rect 6760 1910 6800 1920
rect 7720 1910 7760 1920
rect 680 1900 920 1910
rect 3320 1900 3360 1910
rect 4360 1900 4480 1910
rect 4640 1900 4760 1910
rect 4880 1900 4960 1910
rect 6200 1900 6320 1910
rect 6520 1900 6560 1910
rect 6760 1900 6800 1910
rect 7720 1900 7760 1910
rect 640 1890 920 1900
rect 2480 1890 2720 1900
rect 3320 1890 3360 1900
rect 4280 1890 4400 1900
rect 4440 1890 4480 1900
rect 4600 1890 4640 1900
rect 4680 1890 4760 1900
rect 4800 1890 4840 1900
rect 4920 1890 4960 1900
rect 6160 1890 6360 1900
rect 6480 1890 6600 1900
rect 6760 1890 6800 1900
rect 7720 1890 7800 1900
rect 640 1880 920 1890
rect 2480 1880 2720 1890
rect 3320 1880 3360 1890
rect 4280 1880 4400 1890
rect 4440 1880 4480 1890
rect 4600 1880 4640 1890
rect 4680 1880 4760 1890
rect 4800 1880 4840 1890
rect 4920 1880 4960 1890
rect 6160 1880 6360 1890
rect 6480 1880 6600 1890
rect 6760 1880 6800 1890
rect 7720 1880 7800 1890
rect 640 1870 920 1880
rect 2480 1870 2720 1880
rect 3320 1870 3360 1880
rect 4280 1870 4400 1880
rect 4440 1870 4480 1880
rect 4600 1870 4640 1880
rect 4680 1870 4760 1880
rect 4800 1870 4840 1880
rect 4920 1870 4960 1880
rect 6160 1870 6360 1880
rect 6480 1870 6600 1880
rect 6760 1870 6800 1880
rect 7720 1870 7800 1880
rect 640 1860 920 1870
rect 2480 1860 2720 1870
rect 3320 1860 3360 1870
rect 4280 1860 4400 1870
rect 4440 1860 4480 1870
rect 4600 1860 4640 1870
rect 4680 1860 4760 1870
rect 4800 1860 4840 1870
rect 4920 1860 4960 1870
rect 6160 1860 6360 1870
rect 6480 1860 6600 1870
rect 6760 1860 6800 1870
rect 7720 1860 7800 1870
rect 640 1850 920 1860
rect 2400 1850 2760 1860
rect 2800 1850 2840 1860
rect 3320 1850 3360 1860
rect 4280 1850 4480 1860
rect 4600 1850 4640 1860
rect 4680 1850 4720 1860
rect 4800 1850 4840 1860
rect 6120 1850 6280 1860
rect 6480 1850 6600 1860
rect 7720 1850 7800 1860
rect 640 1840 920 1850
rect 2400 1840 2760 1850
rect 2800 1840 2840 1850
rect 3320 1840 3360 1850
rect 4280 1840 4480 1850
rect 4600 1840 4640 1850
rect 4680 1840 4720 1850
rect 4800 1840 4840 1850
rect 6120 1840 6280 1850
rect 6480 1840 6600 1850
rect 7720 1840 7800 1850
rect 640 1830 920 1840
rect 2400 1830 2760 1840
rect 2800 1830 2840 1840
rect 3320 1830 3360 1840
rect 4280 1830 4480 1840
rect 4600 1830 4640 1840
rect 4680 1830 4720 1840
rect 4800 1830 4840 1840
rect 6120 1830 6280 1840
rect 6480 1830 6600 1840
rect 7720 1830 7800 1840
rect 640 1820 920 1830
rect 2400 1820 2760 1830
rect 2800 1820 2840 1830
rect 3320 1820 3360 1830
rect 4280 1820 4480 1830
rect 4600 1820 4640 1830
rect 4680 1820 4720 1830
rect 4800 1820 4840 1830
rect 6120 1820 6280 1830
rect 6480 1820 6600 1830
rect 7720 1820 7800 1830
rect 600 1810 920 1820
rect 2320 1810 2760 1820
rect 4280 1810 4360 1820
rect 4400 1810 4480 1820
rect 4520 1810 4560 1820
rect 4640 1810 4720 1820
rect 6080 1810 6280 1820
rect 6520 1810 6600 1820
rect 7760 1810 7800 1820
rect 9120 1810 9200 1820
rect 600 1800 920 1810
rect 2320 1800 2760 1810
rect 4280 1800 4360 1810
rect 4400 1800 4480 1810
rect 4520 1800 4560 1810
rect 4640 1800 4720 1810
rect 6080 1800 6280 1810
rect 6520 1800 6600 1810
rect 7760 1800 7800 1810
rect 9120 1800 9200 1810
rect 600 1790 920 1800
rect 2320 1790 2760 1800
rect 4280 1790 4360 1800
rect 4400 1790 4480 1800
rect 4520 1790 4560 1800
rect 4640 1790 4720 1800
rect 6080 1790 6280 1800
rect 6520 1790 6600 1800
rect 7760 1790 7800 1800
rect 9120 1790 9200 1800
rect 600 1780 920 1790
rect 2320 1780 2760 1790
rect 4280 1780 4360 1790
rect 4400 1780 4480 1790
rect 4520 1780 4560 1790
rect 4640 1780 4720 1790
rect 6080 1780 6280 1790
rect 6520 1780 6600 1790
rect 7760 1780 7800 1790
rect 9120 1780 9200 1790
rect 600 1770 920 1780
rect 1840 1770 1880 1780
rect 3280 1770 3320 1780
rect 4040 1770 4080 1780
rect 4280 1770 4360 1780
rect 4400 1770 4480 1780
rect 4560 1770 4600 1780
rect 4640 1770 4720 1780
rect 5200 1770 5240 1780
rect 6040 1770 6320 1780
rect 6560 1770 6640 1780
rect 7760 1770 7800 1780
rect 8360 1770 8400 1780
rect 9120 1770 9200 1780
rect 600 1760 920 1770
rect 1840 1760 1880 1770
rect 3280 1760 3320 1770
rect 4040 1760 4080 1770
rect 4280 1760 4360 1770
rect 4400 1760 4480 1770
rect 4560 1760 4600 1770
rect 4640 1760 4720 1770
rect 5200 1760 5240 1770
rect 6040 1760 6320 1770
rect 6560 1760 6640 1770
rect 7760 1760 7800 1770
rect 8360 1760 8400 1770
rect 9120 1760 9200 1770
rect 600 1750 920 1760
rect 1840 1750 1880 1760
rect 3280 1750 3320 1760
rect 4040 1750 4080 1760
rect 4280 1750 4360 1760
rect 4400 1750 4480 1760
rect 4560 1750 4600 1760
rect 4640 1750 4720 1760
rect 5200 1750 5240 1760
rect 6040 1750 6320 1760
rect 6560 1750 6640 1760
rect 7760 1750 7800 1760
rect 8360 1750 8400 1760
rect 9120 1750 9200 1760
rect 600 1740 920 1750
rect 1840 1740 1880 1750
rect 3280 1740 3320 1750
rect 4040 1740 4080 1750
rect 4280 1740 4360 1750
rect 4400 1740 4480 1750
rect 4560 1740 4600 1750
rect 4640 1740 4720 1750
rect 5200 1740 5240 1750
rect 6040 1740 6320 1750
rect 6560 1740 6640 1750
rect 7760 1740 7800 1750
rect 8360 1740 8400 1750
rect 9120 1740 9200 1750
rect 560 1730 880 1740
rect 3280 1730 3320 1740
rect 4280 1730 4320 1740
rect 4360 1730 4480 1740
rect 6040 1730 6320 1740
rect 6560 1730 6680 1740
rect 7760 1730 7800 1740
rect 9120 1730 9160 1740
rect 560 1720 880 1730
rect 3280 1720 3320 1730
rect 4280 1720 4320 1730
rect 4360 1720 4480 1730
rect 6040 1720 6320 1730
rect 6560 1720 6680 1730
rect 7760 1720 7800 1730
rect 9120 1720 9160 1730
rect 560 1710 880 1720
rect 3280 1710 3320 1720
rect 4280 1710 4320 1720
rect 4360 1710 4480 1720
rect 6040 1710 6320 1720
rect 6560 1710 6680 1720
rect 7760 1710 7800 1720
rect 9120 1710 9160 1720
rect 560 1700 880 1710
rect 3280 1700 3320 1710
rect 4280 1700 4320 1710
rect 4360 1700 4480 1710
rect 6040 1700 6320 1710
rect 6560 1700 6680 1710
rect 7760 1700 7800 1710
rect 9120 1700 9160 1710
rect 560 1690 880 1700
rect 3240 1690 3280 1700
rect 4040 1690 4080 1700
rect 4280 1690 4320 1700
rect 4360 1690 4400 1700
rect 4440 1690 4480 1700
rect 4520 1690 4560 1700
rect 6000 1690 6200 1700
rect 6240 1690 6320 1700
rect 6520 1690 6680 1700
rect 7760 1690 7800 1700
rect 8360 1690 8400 1700
rect 560 1680 880 1690
rect 3240 1680 3280 1690
rect 4040 1680 4080 1690
rect 4280 1680 4320 1690
rect 4360 1680 4400 1690
rect 4440 1680 4480 1690
rect 4520 1680 4560 1690
rect 6000 1680 6200 1690
rect 6240 1680 6320 1690
rect 6520 1680 6680 1690
rect 7760 1680 7800 1690
rect 8360 1680 8400 1690
rect 560 1670 880 1680
rect 3240 1670 3280 1680
rect 4040 1670 4080 1680
rect 4280 1670 4320 1680
rect 4360 1670 4400 1680
rect 4440 1670 4480 1680
rect 4520 1670 4560 1680
rect 6000 1670 6200 1680
rect 6240 1670 6320 1680
rect 6520 1670 6680 1680
rect 7760 1670 7800 1680
rect 8360 1670 8400 1680
rect 560 1660 880 1670
rect 3240 1660 3280 1670
rect 4040 1660 4080 1670
rect 4280 1660 4320 1670
rect 4360 1660 4400 1670
rect 4440 1660 4480 1670
rect 4520 1660 4560 1670
rect 6000 1660 6200 1670
rect 6240 1660 6320 1670
rect 6520 1660 6680 1670
rect 7760 1660 7800 1670
rect 8360 1660 8400 1670
rect 560 1650 880 1660
rect 1880 1650 1920 1660
rect 3240 1650 3280 1660
rect 4280 1650 4320 1660
rect 4360 1650 4400 1660
rect 4560 1650 4600 1660
rect 4640 1650 4720 1660
rect 4760 1650 4800 1660
rect 6000 1650 6200 1660
rect 6280 1650 6320 1660
rect 6520 1650 6680 1660
rect 7760 1650 7800 1660
rect 560 1640 880 1650
rect 1880 1640 1920 1650
rect 3240 1640 3280 1650
rect 4280 1640 4320 1650
rect 4360 1640 4400 1650
rect 4560 1640 4600 1650
rect 4640 1640 4720 1650
rect 4760 1640 4800 1650
rect 6000 1640 6200 1650
rect 6280 1640 6320 1650
rect 6520 1640 6680 1650
rect 7760 1640 7800 1650
rect 560 1630 880 1640
rect 1880 1630 1920 1640
rect 3240 1630 3280 1640
rect 4280 1630 4320 1640
rect 4360 1630 4400 1640
rect 4560 1630 4600 1640
rect 4640 1630 4720 1640
rect 4760 1630 4800 1640
rect 6000 1630 6200 1640
rect 6280 1630 6320 1640
rect 6520 1630 6680 1640
rect 7760 1630 7800 1640
rect 560 1620 880 1630
rect 1880 1620 1920 1630
rect 3240 1620 3280 1630
rect 4280 1620 4320 1630
rect 4360 1620 4400 1630
rect 4560 1620 4600 1630
rect 4640 1620 4720 1630
rect 4760 1620 4800 1630
rect 6000 1620 6200 1630
rect 6280 1620 6320 1630
rect 6520 1620 6680 1630
rect 7760 1620 7800 1630
rect 520 1610 880 1620
rect 3200 1610 3240 1620
rect 4080 1610 4120 1620
rect 4320 1610 4400 1620
rect 4440 1610 4840 1620
rect 5960 1610 6200 1620
rect 6280 1610 6320 1620
rect 6440 1610 6720 1620
rect 7360 1610 7400 1620
rect 7760 1610 7800 1620
rect 8320 1610 8360 1620
rect 520 1600 880 1610
rect 3200 1600 3240 1610
rect 4080 1600 4120 1610
rect 4320 1600 4400 1610
rect 4440 1600 4840 1610
rect 5960 1600 6200 1610
rect 6280 1600 6320 1610
rect 6440 1600 6720 1610
rect 7360 1600 7400 1610
rect 7760 1600 7800 1610
rect 8320 1600 8360 1610
rect 520 1590 880 1600
rect 3200 1590 3240 1600
rect 4080 1590 4120 1600
rect 4320 1590 4400 1600
rect 4440 1590 4840 1600
rect 5960 1590 6200 1600
rect 6280 1590 6320 1600
rect 6440 1590 6720 1600
rect 7360 1590 7400 1600
rect 7760 1590 7800 1600
rect 8320 1590 8360 1600
rect 520 1580 880 1590
rect 3200 1580 3240 1590
rect 4080 1580 4120 1590
rect 4320 1580 4400 1590
rect 4440 1580 4840 1590
rect 5960 1580 6200 1590
rect 6280 1580 6320 1590
rect 6440 1580 6720 1590
rect 7360 1580 7400 1590
rect 7760 1580 7800 1590
rect 8320 1580 8360 1590
rect 520 1570 840 1580
rect 1920 1570 1960 1580
rect 4080 1570 4120 1580
rect 4320 1570 4360 1580
rect 4480 1570 4800 1580
rect 5960 1570 6240 1580
rect 6280 1570 6320 1580
rect 6400 1570 6720 1580
rect 7360 1570 7400 1580
rect 7760 1570 7840 1580
rect 8320 1570 8400 1580
rect 520 1560 840 1570
rect 1920 1560 1960 1570
rect 4080 1560 4120 1570
rect 4320 1560 4360 1570
rect 4480 1560 4800 1570
rect 5960 1560 6240 1570
rect 6280 1560 6320 1570
rect 6400 1560 6720 1570
rect 7360 1560 7400 1570
rect 7760 1560 7840 1570
rect 8320 1560 8400 1570
rect 520 1550 840 1560
rect 1920 1550 1960 1560
rect 4080 1550 4120 1560
rect 4320 1550 4360 1560
rect 4480 1550 4800 1560
rect 5960 1550 6240 1560
rect 6280 1550 6320 1560
rect 6400 1550 6720 1560
rect 7360 1550 7400 1560
rect 7760 1550 7840 1560
rect 8320 1550 8400 1560
rect 520 1540 840 1550
rect 1920 1540 1960 1550
rect 4080 1540 4120 1550
rect 4320 1540 4360 1550
rect 4480 1540 4800 1550
rect 5960 1540 6240 1550
rect 6280 1540 6320 1550
rect 6400 1540 6720 1550
rect 7360 1540 7400 1550
rect 7760 1540 7840 1550
rect 8320 1540 8400 1550
rect 520 1530 840 1540
rect 1960 1530 2000 1540
rect 3160 1530 3200 1540
rect 4360 1530 4920 1540
rect 5960 1530 6240 1540
rect 6280 1530 6320 1540
rect 6400 1530 6800 1540
rect 7800 1530 7840 1540
rect 8320 1530 8360 1540
rect 9760 1530 9800 1540
rect 520 1520 840 1530
rect 1960 1520 2000 1530
rect 3160 1520 3200 1530
rect 4360 1520 4920 1530
rect 5960 1520 6240 1530
rect 6280 1520 6320 1530
rect 6400 1520 6800 1530
rect 7800 1520 7840 1530
rect 8320 1520 8360 1530
rect 9760 1520 9800 1530
rect 520 1510 840 1520
rect 1960 1510 2000 1520
rect 3160 1510 3200 1520
rect 4360 1510 4920 1520
rect 5960 1510 6240 1520
rect 6280 1510 6320 1520
rect 6400 1510 6800 1520
rect 7800 1510 7840 1520
rect 8320 1510 8360 1520
rect 9760 1510 9800 1520
rect 520 1500 840 1510
rect 1960 1500 2000 1510
rect 3160 1500 3200 1510
rect 4360 1500 4920 1510
rect 5960 1500 6240 1510
rect 6280 1500 6320 1510
rect 6400 1500 6800 1510
rect 7800 1500 7840 1510
rect 8320 1500 8360 1510
rect 9760 1500 9800 1510
rect 480 1490 840 1500
rect 920 1490 1000 1500
rect 3120 1490 3160 1500
rect 4360 1490 4440 1500
rect 4480 1490 5000 1500
rect 5880 1490 6200 1500
rect 6280 1490 6320 1500
rect 6360 1490 6800 1500
rect 7800 1490 7840 1500
rect 8320 1490 8360 1500
rect 9720 1490 9800 1500
rect 480 1480 840 1490
rect 920 1480 1000 1490
rect 3120 1480 3160 1490
rect 4360 1480 4440 1490
rect 4480 1480 5000 1490
rect 5880 1480 6200 1490
rect 6280 1480 6320 1490
rect 6360 1480 6800 1490
rect 7800 1480 7840 1490
rect 8320 1480 8360 1490
rect 9720 1480 9800 1490
rect 480 1470 840 1480
rect 920 1470 1000 1480
rect 3120 1470 3160 1480
rect 4360 1470 4440 1480
rect 4480 1470 5000 1480
rect 5880 1470 6200 1480
rect 6280 1470 6320 1480
rect 6360 1470 6800 1480
rect 7800 1470 7840 1480
rect 8320 1470 8360 1480
rect 9720 1470 9800 1480
rect 480 1460 840 1470
rect 920 1460 1000 1470
rect 3120 1460 3160 1470
rect 4360 1460 4440 1470
rect 4480 1460 5000 1470
rect 5880 1460 6200 1470
rect 6280 1460 6320 1470
rect 6360 1460 6800 1470
rect 7800 1460 7840 1470
rect 8320 1460 8360 1470
rect 9720 1460 9800 1470
rect 480 1450 880 1460
rect 1000 1450 1040 1460
rect 2000 1450 2040 1460
rect 3040 1450 3120 1460
rect 4120 1450 4160 1460
rect 4440 1450 5040 1460
rect 5880 1450 6200 1460
rect 6320 1450 6800 1460
rect 7800 1450 7840 1460
rect 8320 1450 8360 1460
rect 9720 1450 9760 1460
rect 480 1440 880 1450
rect 1000 1440 1040 1450
rect 2000 1440 2040 1450
rect 3040 1440 3120 1450
rect 4120 1440 4160 1450
rect 4440 1440 5040 1450
rect 5880 1440 6200 1450
rect 6320 1440 6800 1450
rect 7800 1440 7840 1450
rect 8320 1440 8360 1450
rect 9720 1440 9760 1450
rect 480 1430 880 1440
rect 1000 1430 1040 1440
rect 2000 1430 2040 1440
rect 3040 1430 3120 1440
rect 4120 1430 4160 1440
rect 4440 1430 5040 1440
rect 5880 1430 6200 1440
rect 6320 1430 6800 1440
rect 7800 1430 7840 1440
rect 8320 1430 8360 1440
rect 9720 1430 9760 1440
rect 480 1420 880 1430
rect 1000 1420 1040 1430
rect 2000 1420 2040 1430
rect 3040 1420 3120 1430
rect 4120 1420 4160 1430
rect 4440 1420 5040 1430
rect 5880 1420 6200 1430
rect 6320 1420 6800 1430
rect 7800 1420 7840 1430
rect 8320 1420 8360 1430
rect 9720 1420 9760 1430
rect 480 1410 840 1420
rect 1000 1410 1040 1420
rect 2040 1410 2080 1420
rect 3000 1410 3080 1420
rect 4440 1410 5120 1420
rect 5920 1410 6200 1420
rect 6320 1410 6800 1420
rect 7800 1410 7840 1420
rect 8280 1410 8360 1420
rect 9720 1410 9760 1420
rect 480 1400 840 1410
rect 1000 1400 1040 1410
rect 2040 1400 2080 1410
rect 3000 1400 3080 1410
rect 4440 1400 5120 1410
rect 5920 1400 6200 1410
rect 6320 1400 6800 1410
rect 7800 1400 7840 1410
rect 8280 1400 8360 1410
rect 9720 1400 9760 1410
rect 480 1390 840 1400
rect 1000 1390 1040 1400
rect 2040 1390 2080 1400
rect 3000 1390 3080 1400
rect 4440 1390 5120 1400
rect 5920 1390 6200 1400
rect 6320 1390 6800 1400
rect 7800 1390 7840 1400
rect 8280 1390 8360 1400
rect 9720 1390 9760 1400
rect 480 1380 840 1390
rect 1000 1380 1040 1390
rect 2040 1380 2080 1390
rect 3000 1380 3080 1390
rect 4440 1380 5120 1390
rect 5920 1380 6200 1390
rect 6320 1380 6800 1390
rect 7800 1380 7840 1390
rect 8280 1380 8360 1390
rect 9720 1380 9760 1390
rect 440 1370 840 1380
rect 960 1370 1040 1380
rect 2080 1370 2120 1380
rect 2960 1370 3000 1380
rect 3520 1370 3560 1380
rect 4400 1370 5120 1380
rect 5920 1370 6200 1380
rect 6320 1370 6800 1380
rect 8280 1370 8320 1380
rect 9680 1370 9720 1380
rect 440 1360 840 1370
rect 960 1360 1040 1370
rect 2080 1360 2120 1370
rect 2960 1360 3000 1370
rect 3520 1360 3560 1370
rect 4400 1360 5120 1370
rect 5920 1360 6200 1370
rect 6320 1360 6800 1370
rect 8280 1360 8320 1370
rect 9680 1360 9720 1370
rect 440 1350 840 1360
rect 960 1350 1040 1360
rect 2080 1350 2120 1360
rect 2960 1350 3000 1360
rect 3520 1350 3560 1360
rect 4400 1350 5120 1360
rect 5920 1350 6200 1360
rect 6320 1350 6800 1360
rect 8280 1350 8320 1360
rect 9680 1350 9720 1360
rect 440 1340 840 1350
rect 960 1340 1040 1350
rect 2080 1340 2120 1350
rect 2960 1340 3000 1350
rect 3520 1340 3560 1350
rect 4400 1340 5120 1350
rect 5920 1340 6200 1350
rect 6320 1340 6800 1350
rect 8280 1340 8320 1350
rect 9680 1340 9720 1350
rect 440 1330 840 1340
rect 920 1330 1040 1340
rect 2080 1330 2160 1340
rect 2800 1330 2960 1340
rect 3480 1330 3520 1340
rect 4160 1330 4200 1340
rect 4440 1330 5040 1340
rect 5200 1330 5240 1340
rect 5440 1330 5480 1340
rect 5920 1330 6200 1340
rect 6320 1330 6800 1340
rect 440 1320 840 1330
rect 920 1320 1040 1330
rect 2080 1320 2160 1330
rect 2800 1320 2960 1330
rect 3480 1320 3520 1330
rect 4160 1320 4200 1330
rect 4440 1320 5040 1330
rect 5200 1320 5240 1330
rect 5440 1320 5480 1330
rect 5920 1320 6200 1330
rect 6320 1320 6800 1330
rect 440 1310 840 1320
rect 920 1310 1040 1320
rect 2080 1310 2160 1320
rect 2800 1310 2960 1320
rect 3480 1310 3520 1320
rect 4160 1310 4200 1320
rect 4440 1310 5040 1320
rect 5200 1310 5240 1320
rect 5440 1310 5480 1320
rect 5920 1310 6200 1320
rect 6320 1310 6800 1320
rect 440 1300 840 1310
rect 920 1300 1040 1310
rect 2080 1300 2160 1310
rect 2800 1300 2960 1310
rect 3480 1300 3520 1310
rect 4160 1300 4200 1310
rect 4440 1300 5040 1310
rect 5200 1300 5240 1310
rect 5440 1300 5480 1310
rect 5920 1300 6200 1310
rect 6320 1300 6800 1310
rect 440 1290 800 1300
rect 920 1290 1000 1300
rect 2040 1290 2200 1300
rect 2720 1290 2880 1300
rect 3720 1290 3760 1300
rect 4440 1290 4960 1300
rect 5120 1290 5160 1300
rect 5200 1290 5240 1300
rect 5920 1290 6200 1300
rect 6320 1290 6800 1300
rect 7400 1290 7440 1300
rect 7840 1290 7880 1300
rect 9200 1290 9240 1300
rect 440 1280 800 1290
rect 920 1280 1000 1290
rect 2040 1280 2200 1290
rect 2720 1280 2880 1290
rect 3720 1280 3760 1290
rect 4440 1280 4960 1290
rect 5120 1280 5160 1290
rect 5200 1280 5240 1290
rect 5920 1280 6200 1290
rect 6320 1280 6800 1290
rect 7400 1280 7440 1290
rect 7840 1280 7880 1290
rect 9200 1280 9240 1290
rect 440 1270 800 1280
rect 920 1270 1000 1280
rect 2040 1270 2200 1280
rect 2720 1270 2880 1280
rect 3720 1270 3760 1280
rect 4440 1270 4960 1280
rect 5120 1270 5160 1280
rect 5200 1270 5240 1280
rect 5920 1270 6200 1280
rect 6320 1270 6800 1280
rect 7400 1270 7440 1280
rect 7840 1270 7880 1280
rect 9200 1270 9240 1280
rect 440 1260 800 1270
rect 920 1260 1000 1270
rect 2040 1260 2200 1270
rect 2720 1260 2880 1270
rect 3720 1260 3760 1270
rect 4440 1260 4960 1270
rect 5120 1260 5160 1270
rect 5200 1260 5240 1270
rect 5920 1260 6200 1270
rect 6320 1260 6800 1270
rect 7400 1260 7440 1270
rect 7840 1260 7880 1270
rect 9200 1260 9240 1270
rect 400 1250 800 1260
rect 920 1250 1000 1260
rect 2040 1250 2240 1260
rect 2640 1250 2840 1260
rect 3480 1250 3520 1260
rect 4440 1250 5000 1260
rect 5920 1250 6240 1260
rect 6320 1250 6760 1260
rect 7400 1250 7440 1260
rect 7840 1250 7880 1260
rect 9160 1250 9240 1260
rect 400 1240 800 1250
rect 920 1240 1000 1250
rect 2040 1240 2240 1250
rect 2640 1240 2840 1250
rect 3480 1240 3520 1250
rect 4440 1240 5000 1250
rect 5920 1240 6240 1250
rect 6320 1240 6760 1250
rect 7400 1240 7440 1250
rect 7840 1240 7880 1250
rect 9160 1240 9240 1250
rect 400 1230 800 1240
rect 920 1230 1000 1240
rect 2040 1230 2240 1240
rect 2640 1230 2840 1240
rect 3480 1230 3520 1240
rect 4440 1230 5000 1240
rect 5920 1230 6240 1240
rect 6320 1230 6760 1240
rect 7400 1230 7440 1240
rect 7840 1230 7880 1240
rect 9160 1230 9240 1240
rect 400 1220 800 1230
rect 920 1220 1000 1230
rect 2040 1220 2240 1230
rect 2640 1220 2840 1230
rect 3480 1220 3520 1230
rect 4440 1220 5000 1230
rect 5920 1220 6240 1230
rect 6320 1220 6760 1230
rect 7400 1220 7440 1230
rect 7840 1220 7880 1230
rect 9160 1220 9240 1230
rect 400 1210 800 1220
rect 880 1210 1000 1220
rect 2000 1210 2120 1220
rect 2240 1210 2320 1220
rect 2600 1210 2760 1220
rect 4480 1210 4720 1220
rect 4920 1210 4960 1220
rect 5920 1210 6240 1220
rect 6360 1210 6680 1220
rect 7400 1210 7440 1220
rect 7840 1210 7880 1220
rect 9200 1210 9240 1220
rect 9760 1210 9800 1220
rect 400 1200 800 1210
rect 880 1200 1000 1210
rect 2000 1200 2120 1210
rect 2240 1200 2320 1210
rect 2600 1200 2760 1210
rect 4480 1200 4720 1210
rect 4920 1200 4960 1210
rect 5920 1200 6240 1210
rect 6360 1200 6680 1210
rect 7400 1200 7440 1210
rect 7840 1200 7880 1210
rect 9200 1200 9240 1210
rect 9760 1200 9800 1210
rect 400 1190 800 1200
rect 880 1190 1000 1200
rect 2000 1190 2120 1200
rect 2240 1190 2320 1200
rect 2600 1190 2760 1200
rect 4480 1190 4720 1200
rect 4920 1190 4960 1200
rect 5920 1190 6240 1200
rect 6360 1190 6680 1200
rect 7400 1190 7440 1200
rect 7840 1190 7880 1200
rect 9200 1190 9240 1200
rect 9760 1190 9800 1200
rect 400 1180 800 1190
rect 880 1180 1000 1190
rect 2000 1180 2120 1190
rect 2240 1180 2320 1190
rect 2600 1180 2760 1190
rect 4480 1180 4720 1190
rect 4920 1180 4960 1190
rect 5920 1180 6240 1190
rect 6360 1180 6680 1190
rect 7400 1180 7440 1190
rect 7840 1180 7880 1190
rect 9200 1180 9240 1190
rect 9760 1180 9800 1190
rect 400 1170 760 1180
rect 880 1170 1000 1180
rect 2000 1170 2080 1180
rect 2280 1170 2880 1180
rect 4480 1170 4560 1180
rect 4920 1170 5000 1180
rect 5040 1170 5360 1180
rect 5920 1170 6280 1180
rect 6360 1170 6640 1180
rect 7400 1170 7440 1180
rect 7880 1170 7920 1180
rect 9200 1170 9240 1180
rect 9760 1170 9800 1180
rect 400 1160 760 1170
rect 880 1160 1000 1170
rect 2000 1160 2080 1170
rect 2280 1160 2880 1170
rect 4480 1160 4560 1170
rect 4920 1160 5000 1170
rect 5040 1160 5360 1170
rect 5920 1160 6280 1170
rect 6360 1160 6640 1170
rect 7400 1160 7440 1170
rect 7880 1160 7920 1170
rect 9200 1160 9240 1170
rect 9760 1160 9800 1170
rect 400 1150 760 1160
rect 880 1150 1000 1160
rect 2000 1150 2080 1160
rect 2280 1150 2880 1160
rect 4480 1150 4560 1160
rect 4920 1150 5000 1160
rect 5040 1150 5360 1160
rect 5920 1150 6280 1160
rect 6360 1150 6640 1160
rect 7400 1150 7440 1160
rect 7880 1150 7920 1160
rect 9200 1150 9240 1160
rect 9760 1150 9800 1160
rect 400 1140 760 1150
rect 880 1140 1000 1150
rect 2000 1140 2080 1150
rect 2280 1140 2880 1150
rect 4480 1140 4560 1150
rect 4920 1140 5000 1150
rect 5040 1140 5360 1150
rect 5920 1140 6280 1150
rect 6360 1140 6640 1150
rect 7400 1140 7440 1150
rect 7880 1140 7920 1150
rect 9200 1140 9240 1150
rect 9760 1140 9800 1150
rect 360 1130 640 1140
rect 880 1130 1000 1140
rect 1560 1130 1600 1140
rect 2000 1130 2040 1140
rect 2360 1130 2880 1140
rect 4480 1130 4560 1140
rect 4760 1130 5400 1140
rect 5680 1130 5720 1140
rect 5920 1130 6280 1140
rect 6400 1130 6560 1140
rect 7400 1130 7440 1140
rect 7880 1130 7920 1140
rect 9760 1130 9800 1140
rect 360 1120 640 1130
rect 880 1120 1000 1130
rect 1560 1120 1600 1130
rect 2000 1120 2040 1130
rect 2360 1120 2880 1130
rect 4480 1120 4560 1130
rect 4760 1120 5400 1130
rect 5680 1120 5720 1130
rect 5920 1120 6280 1130
rect 6400 1120 6560 1130
rect 7400 1120 7440 1130
rect 7880 1120 7920 1130
rect 9760 1120 9800 1130
rect 360 1110 640 1120
rect 880 1110 1000 1120
rect 1560 1110 1600 1120
rect 2000 1110 2040 1120
rect 2360 1110 2880 1120
rect 4480 1110 4560 1120
rect 4760 1110 5400 1120
rect 5680 1110 5720 1120
rect 5920 1110 6280 1120
rect 6400 1110 6560 1120
rect 7400 1110 7440 1120
rect 7880 1110 7920 1120
rect 9760 1110 9800 1120
rect 360 1100 640 1110
rect 880 1100 1000 1110
rect 1560 1100 1600 1110
rect 2000 1100 2040 1110
rect 2360 1100 2880 1110
rect 4480 1100 4560 1110
rect 4760 1100 5400 1110
rect 5680 1100 5720 1110
rect 5920 1100 6280 1110
rect 6400 1100 6560 1110
rect 7400 1100 7440 1110
rect 7880 1100 7920 1110
rect 9760 1100 9800 1110
rect 360 1090 640 1100
rect 720 1090 760 1100
rect 880 1090 1000 1100
rect 1480 1090 1520 1100
rect 1960 1090 2000 1100
rect 2840 1090 2920 1100
rect 4080 1090 4120 1100
rect 4480 1090 5480 1100
rect 5640 1090 5880 1100
rect 5960 1090 6280 1100
rect 6440 1090 6480 1100
rect 7400 1090 7440 1100
rect 7880 1090 7920 1100
rect 9760 1090 9800 1100
rect 360 1080 640 1090
rect 720 1080 760 1090
rect 880 1080 1000 1090
rect 1480 1080 1520 1090
rect 1960 1080 2000 1090
rect 2840 1080 2920 1090
rect 4080 1080 4120 1090
rect 4480 1080 5480 1090
rect 5640 1080 5880 1090
rect 5960 1080 6280 1090
rect 6440 1080 6480 1090
rect 7400 1080 7440 1090
rect 7880 1080 7920 1090
rect 9760 1080 9800 1090
rect 360 1070 640 1080
rect 720 1070 760 1080
rect 880 1070 1000 1080
rect 1480 1070 1520 1080
rect 1960 1070 2000 1080
rect 2840 1070 2920 1080
rect 4080 1070 4120 1080
rect 4480 1070 5480 1080
rect 5640 1070 5880 1080
rect 5960 1070 6280 1080
rect 6440 1070 6480 1080
rect 7400 1070 7440 1080
rect 7880 1070 7920 1080
rect 9760 1070 9800 1080
rect 360 1060 640 1070
rect 720 1060 760 1070
rect 880 1060 1000 1070
rect 1480 1060 1520 1070
rect 1960 1060 2000 1070
rect 2840 1060 2920 1070
rect 4080 1060 4120 1070
rect 4480 1060 5480 1070
rect 5640 1060 5880 1070
rect 5960 1060 6280 1070
rect 6440 1060 6480 1070
rect 7400 1060 7440 1070
rect 7880 1060 7920 1070
rect 9760 1060 9800 1070
rect 320 1050 640 1060
rect 840 1050 960 1060
rect 1440 1050 1480 1060
rect 1640 1050 1680 1060
rect 1960 1050 2000 1060
rect 2840 1050 2920 1060
rect 4080 1050 4120 1060
rect 4640 1050 5480 1060
rect 5520 1050 5840 1060
rect 5880 1050 6280 1060
rect 6400 1050 6440 1060
rect 7880 1050 7920 1060
rect 9760 1050 9800 1060
rect 320 1040 640 1050
rect 840 1040 960 1050
rect 1440 1040 1480 1050
rect 1640 1040 1680 1050
rect 1960 1040 2000 1050
rect 2840 1040 2920 1050
rect 4080 1040 4120 1050
rect 4640 1040 5480 1050
rect 5520 1040 5840 1050
rect 5880 1040 6280 1050
rect 6400 1040 6440 1050
rect 7880 1040 7920 1050
rect 9760 1040 9800 1050
rect 320 1030 640 1040
rect 840 1030 960 1040
rect 1440 1030 1480 1040
rect 1640 1030 1680 1040
rect 1960 1030 2000 1040
rect 2840 1030 2920 1040
rect 4080 1030 4120 1040
rect 4640 1030 5480 1040
rect 5520 1030 5840 1040
rect 5880 1030 6280 1040
rect 6400 1030 6440 1040
rect 7880 1030 7920 1040
rect 9760 1030 9800 1040
rect 320 1020 640 1030
rect 840 1020 960 1030
rect 1440 1020 1480 1030
rect 1640 1020 1680 1030
rect 1960 1020 2000 1030
rect 2840 1020 2920 1030
rect 4080 1020 4120 1030
rect 4640 1020 5480 1030
rect 5520 1020 5840 1030
rect 5880 1020 6280 1030
rect 6400 1020 6440 1030
rect 7880 1020 7920 1030
rect 9760 1020 9800 1030
rect 320 1010 680 1020
rect 840 1010 960 1020
rect 1400 1010 1440 1020
rect 1560 1010 1640 1020
rect 1960 1010 2000 1020
rect 2840 1010 2920 1020
rect 3680 1010 3720 1020
rect 4160 1010 4200 1020
rect 4720 1010 5440 1020
rect 5520 1010 5600 1020
rect 5640 1010 6320 1020
rect 6360 1010 6400 1020
rect 7880 1010 7920 1020
rect 9000 1010 9080 1020
rect 320 1000 680 1010
rect 840 1000 960 1010
rect 1400 1000 1440 1010
rect 1560 1000 1640 1010
rect 1960 1000 2000 1010
rect 2840 1000 2920 1010
rect 3680 1000 3720 1010
rect 4160 1000 4200 1010
rect 4720 1000 5440 1010
rect 5520 1000 5600 1010
rect 5640 1000 6320 1010
rect 6360 1000 6400 1010
rect 7880 1000 7920 1010
rect 9000 1000 9080 1010
rect 320 990 680 1000
rect 840 990 960 1000
rect 1400 990 1440 1000
rect 1560 990 1640 1000
rect 1960 990 2000 1000
rect 2840 990 2920 1000
rect 3680 990 3720 1000
rect 4160 990 4200 1000
rect 4720 990 5440 1000
rect 5520 990 5600 1000
rect 5640 990 6320 1000
rect 6360 990 6400 1000
rect 7880 990 7920 1000
rect 9000 990 9080 1000
rect 320 980 680 990
rect 840 980 960 990
rect 1400 980 1440 990
rect 1560 980 1640 990
rect 1960 980 2000 990
rect 2840 980 2920 990
rect 3680 980 3720 990
rect 4160 980 4200 990
rect 4720 980 5440 990
rect 5520 980 5600 990
rect 5640 980 6320 990
rect 6360 980 6400 990
rect 7880 980 7920 990
rect 9000 980 9080 990
rect 280 970 720 980
rect 800 970 960 980
rect 1520 970 1600 980
rect 1960 970 2000 980
rect 2840 970 2880 980
rect 4800 970 5320 980
rect 5960 970 6320 980
rect 6360 970 6400 980
rect 8160 970 8200 980
rect 8960 970 9080 980
rect 9480 970 9520 980
rect 280 960 720 970
rect 800 960 960 970
rect 1520 960 1600 970
rect 1960 960 2000 970
rect 2840 960 2880 970
rect 4800 960 5320 970
rect 5960 960 6320 970
rect 6360 960 6400 970
rect 8160 960 8200 970
rect 8960 960 9080 970
rect 9480 960 9520 970
rect 280 950 720 960
rect 800 950 960 960
rect 1520 950 1600 960
rect 1960 950 2000 960
rect 2840 950 2880 960
rect 4800 950 5320 960
rect 5960 950 6320 960
rect 6360 950 6400 960
rect 8160 950 8200 960
rect 8960 950 9080 960
rect 9480 950 9520 960
rect 280 940 720 950
rect 800 940 960 950
rect 1520 940 1600 950
rect 1960 940 2000 950
rect 2840 940 2880 950
rect 4800 940 5320 950
rect 5960 940 6320 950
rect 6360 940 6400 950
rect 8160 940 8200 950
rect 8960 940 9080 950
rect 9480 940 9520 950
rect 280 930 680 940
rect 800 930 960 940
rect 1480 930 1560 940
rect 1960 930 2000 940
rect 2760 930 2840 940
rect 4880 930 5160 940
rect 5200 930 5320 940
rect 6040 930 6200 940
rect 6280 930 6320 940
rect 6360 930 6400 940
rect 7920 930 7960 940
rect 8160 930 8200 940
rect 8920 930 9080 940
rect 280 920 680 930
rect 800 920 960 930
rect 1480 920 1560 930
rect 1960 920 2000 930
rect 2760 920 2840 930
rect 4880 920 5160 930
rect 5200 920 5320 930
rect 6040 920 6200 930
rect 6280 920 6320 930
rect 6360 920 6400 930
rect 7920 920 7960 930
rect 8160 920 8200 930
rect 8920 920 9080 930
rect 280 910 680 920
rect 800 910 960 920
rect 1480 910 1560 920
rect 1960 910 2000 920
rect 2760 910 2840 920
rect 4880 910 5160 920
rect 5200 910 5320 920
rect 6040 910 6200 920
rect 6280 910 6320 920
rect 6360 910 6400 920
rect 7920 910 7960 920
rect 8160 910 8200 920
rect 8920 910 9080 920
rect 280 900 680 910
rect 800 900 960 910
rect 1480 900 1560 910
rect 1960 900 2000 910
rect 2760 900 2840 910
rect 4880 900 5160 910
rect 5200 900 5320 910
rect 6040 900 6200 910
rect 6280 900 6320 910
rect 6360 900 6400 910
rect 7920 900 7960 910
rect 8160 900 8200 910
rect 8920 900 9080 910
rect 240 890 680 900
rect 920 890 960 900
rect 1240 890 1280 900
rect 1440 890 1520 900
rect 2720 890 2760 900
rect 3800 890 3840 900
rect 5080 890 5200 900
rect 5280 890 5320 900
rect 5680 890 5800 900
rect 6040 890 6200 900
rect 6280 890 6320 900
rect 6360 890 6400 900
rect 7920 890 7960 900
rect 8160 890 8200 900
rect 8880 890 9080 900
rect 240 880 680 890
rect 920 880 960 890
rect 1240 880 1280 890
rect 1440 880 1520 890
rect 2720 880 2760 890
rect 3800 880 3840 890
rect 5080 880 5200 890
rect 5280 880 5320 890
rect 5680 880 5800 890
rect 6040 880 6200 890
rect 6280 880 6320 890
rect 6360 880 6400 890
rect 7920 880 7960 890
rect 8160 880 8200 890
rect 8880 880 9080 890
rect 240 870 680 880
rect 920 870 960 880
rect 1240 870 1280 880
rect 1440 870 1520 880
rect 2720 870 2760 880
rect 3800 870 3840 880
rect 5080 870 5200 880
rect 5280 870 5320 880
rect 5680 870 5800 880
rect 6040 870 6200 880
rect 6280 870 6320 880
rect 6360 870 6400 880
rect 7920 870 7960 880
rect 8160 870 8200 880
rect 8880 870 9080 880
rect 240 860 680 870
rect 920 860 960 870
rect 1240 860 1280 870
rect 1440 860 1520 870
rect 2720 860 2760 870
rect 3800 860 3840 870
rect 5080 860 5200 870
rect 5280 860 5320 870
rect 5680 860 5800 870
rect 6040 860 6200 870
rect 6280 860 6320 870
rect 6360 860 6400 870
rect 7920 860 7960 870
rect 8160 860 8200 870
rect 8880 860 9080 870
rect 200 850 640 860
rect 1200 850 1240 860
rect 1400 850 1480 860
rect 2000 850 2040 860
rect 3840 850 3880 860
rect 4880 850 4920 860
rect 5200 850 5320 860
rect 5440 850 5760 860
rect 6040 850 6200 860
rect 6280 850 6320 860
rect 6400 850 6440 860
rect 7920 850 7960 860
rect 8160 850 8200 860
rect 8840 850 9080 860
rect 200 840 640 850
rect 1200 840 1240 850
rect 1400 840 1480 850
rect 2000 840 2040 850
rect 3840 840 3880 850
rect 4880 840 4920 850
rect 5200 840 5320 850
rect 5440 840 5760 850
rect 6040 840 6200 850
rect 6280 840 6320 850
rect 6400 840 6440 850
rect 7920 840 7960 850
rect 8160 840 8200 850
rect 8840 840 9080 850
rect 200 830 640 840
rect 1200 830 1240 840
rect 1400 830 1480 840
rect 2000 830 2040 840
rect 3840 830 3880 840
rect 4880 830 4920 840
rect 5200 830 5320 840
rect 5440 830 5760 840
rect 6040 830 6200 840
rect 6280 830 6320 840
rect 6400 830 6440 840
rect 7920 830 7960 840
rect 8160 830 8200 840
rect 8840 830 9080 840
rect 200 820 640 830
rect 1200 820 1240 830
rect 1400 820 1480 830
rect 2000 820 2040 830
rect 3840 820 3880 830
rect 4880 820 4920 830
rect 5200 820 5320 830
rect 5440 820 5760 830
rect 6040 820 6200 830
rect 6280 820 6320 830
rect 6400 820 6440 830
rect 7920 820 7960 830
rect 8160 820 8200 830
rect 8840 820 9080 830
rect 160 810 640 820
rect 840 810 920 820
rect 1360 810 1480 820
rect 2000 810 2040 820
rect 3880 810 3920 820
rect 5160 810 5480 820
rect 5520 810 5760 820
rect 6040 810 6160 820
rect 6280 810 6320 820
rect 6400 810 6440 820
rect 7400 810 7440 820
rect 7920 810 7960 820
rect 8160 810 8240 820
rect 8840 810 9160 820
rect 160 800 640 810
rect 840 800 920 810
rect 1360 800 1480 810
rect 2000 800 2040 810
rect 3880 800 3920 810
rect 5160 800 5480 810
rect 5520 800 5760 810
rect 6040 800 6160 810
rect 6280 800 6320 810
rect 6400 800 6440 810
rect 7400 800 7440 810
rect 7920 800 7960 810
rect 8160 800 8240 810
rect 8840 800 9160 810
rect 160 790 640 800
rect 840 790 920 800
rect 1360 790 1480 800
rect 2000 790 2040 800
rect 3880 790 3920 800
rect 5160 790 5480 800
rect 5520 790 5760 800
rect 6040 790 6160 800
rect 6280 790 6320 800
rect 6400 790 6440 800
rect 7400 790 7440 800
rect 7920 790 7960 800
rect 8160 790 8240 800
rect 8840 790 9160 800
rect 160 780 640 790
rect 840 780 920 790
rect 1360 780 1480 790
rect 2000 780 2040 790
rect 3880 780 3920 790
rect 5160 780 5480 790
rect 5520 780 5760 790
rect 6040 780 6160 790
rect 6280 780 6320 790
rect 6400 780 6440 790
rect 7400 780 7440 790
rect 7920 780 7960 790
rect 8160 780 8240 790
rect 8840 780 9160 790
rect 120 770 640 780
rect 800 770 920 780
rect 1080 770 1120 780
rect 1280 770 1440 780
rect 2520 770 2560 780
rect 3960 770 4000 780
rect 5320 770 5360 780
rect 5400 770 5760 780
rect 6280 770 6320 780
rect 6400 770 6480 780
rect 7400 770 7440 780
rect 8160 770 8240 780
rect 8800 770 9160 780
rect 120 760 640 770
rect 800 760 920 770
rect 1080 760 1120 770
rect 1280 760 1440 770
rect 2520 760 2560 770
rect 3960 760 4000 770
rect 5320 760 5360 770
rect 5400 760 5760 770
rect 6280 760 6320 770
rect 6400 760 6480 770
rect 7400 760 7440 770
rect 8160 760 8240 770
rect 8800 760 9160 770
rect 120 750 640 760
rect 800 750 920 760
rect 1080 750 1120 760
rect 1280 750 1440 760
rect 2520 750 2560 760
rect 3960 750 4000 760
rect 5320 750 5360 760
rect 5400 750 5760 760
rect 6280 750 6320 760
rect 6400 750 6480 760
rect 7400 750 7440 760
rect 8160 750 8240 760
rect 8800 750 9160 760
rect 120 740 640 750
rect 800 740 920 750
rect 1080 740 1120 750
rect 1280 740 1440 750
rect 2520 740 2560 750
rect 3960 740 4000 750
rect 5320 740 5360 750
rect 5400 740 5760 750
rect 6280 740 6320 750
rect 6400 740 6480 750
rect 7400 740 7440 750
rect 8160 740 8240 750
rect 8800 740 9160 750
rect 80 730 600 740
rect 760 730 920 740
rect 1040 730 1080 740
rect 1280 730 1400 740
rect 2040 730 2080 740
rect 2440 730 2480 740
rect 5120 730 5200 740
rect 5360 730 5400 740
rect 5440 730 5760 740
rect 6280 730 6320 740
rect 6440 730 6480 740
rect 7400 730 7440 740
rect 7960 730 8000 740
rect 8160 730 8240 740
rect 8760 730 9160 740
rect 80 720 600 730
rect 760 720 920 730
rect 1040 720 1080 730
rect 1280 720 1400 730
rect 2040 720 2080 730
rect 2440 720 2480 730
rect 5120 720 5200 730
rect 5360 720 5400 730
rect 5440 720 5760 730
rect 6280 720 6320 730
rect 6440 720 6480 730
rect 7400 720 7440 730
rect 7960 720 8000 730
rect 8160 720 8240 730
rect 8760 720 9160 730
rect 80 710 600 720
rect 760 710 920 720
rect 1040 710 1080 720
rect 1280 710 1400 720
rect 2040 710 2080 720
rect 2440 710 2480 720
rect 5120 710 5200 720
rect 5360 710 5400 720
rect 5440 710 5760 720
rect 6280 710 6320 720
rect 6440 710 6480 720
rect 7400 710 7440 720
rect 7960 710 8000 720
rect 8160 710 8240 720
rect 8760 710 9160 720
rect 80 700 600 710
rect 760 700 920 710
rect 1040 700 1080 710
rect 1280 700 1400 710
rect 2040 700 2080 710
rect 2440 700 2480 710
rect 5120 700 5200 710
rect 5360 700 5400 710
rect 5440 700 5760 710
rect 6280 700 6320 710
rect 6440 700 6480 710
rect 7400 700 7440 710
rect 7960 700 8000 710
rect 8160 700 8240 710
rect 8760 700 9160 710
rect 40 690 600 700
rect 760 690 1000 700
rect 1320 690 1360 700
rect 3280 690 3320 700
rect 4720 690 4760 700
rect 4920 690 4960 700
rect 5120 690 5200 700
rect 5400 690 5440 700
rect 5480 690 5520 700
rect 5640 690 5760 700
rect 6280 690 6360 700
rect 6440 690 6520 700
rect 7400 690 7440 700
rect 7960 690 8000 700
rect 8160 690 8280 700
rect 8760 690 9160 700
rect 40 680 600 690
rect 760 680 1000 690
rect 1320 680 1360 690
rect 3280 680 3320 690
rect 4720 680 4760 690
rect 4920 680 4960 690
rect 5120 680 5200 690
rect 5400 680 5440 690
rect 5480 680 5520 690
rect 5640 680 5760 690
rect 6280 680 6360 690
rect 6440 680 6520 690
rect 7400 680 7440 690
rect 7960 680 8000 690
rect 8160 680 8280 690
rect 8760 680 9160 690
rect 40 670 600 680
rect 760 670 1000 680
rect 1320 670 1360 680
rect 3280 670 3320 680
rect 4720 670 4760 680
rect 4920 670 4960 680
rect 5120 670 5200 680
rect 5400 670 5440 680
rect 5480 670 5520 680
rect 5640 670 5760 680
rect 6280 670 6360 680
rect 6440 670 6520 680
rect 7400 670 7440 680
rect 7960 670 8000 680
rect 8160 670 8280 680
rect 8760 670 9160 680
rect 40 660 600 670
rect 760 660 1000 670
rect 1320 660 1360 670
rect 3280 660 3320 670
rect 4720 660 4760 670
rect 4920 660 4960 670
rect 5120 660 5200 670
rect 5400 660 5440 670
rect 5480 660 5520 670
rect 5640 660 5760 670
rect 6280 660 6360 670
rect 6440 660 6520 670
rect 7400 660 7440 670
rect 7960 660 8000 670
rect 8160 660 8280 670
rect 8760 660 9160 670
rect 0 650 480 660
rect 1280 650 1360 660
rect 2080 650 2120 660
rect 3200 650 3240 660
rect 4720 650 4800 660
rect 5160 650 5200 660
rect 5280 650 5320 660
rect 5400 650 5440 660
rect 5480 650 5560 660
rect 5680 650 5760 660
rect 6280 650 6360 660
rect 6480 650 6520 660
rect 7400 650 7440 660
rect 8160 650 8320 660
rect 8720 650 9120 660
rect 0 640 480 650
rect 1280 640 1360 650
rect 2080 640 2120 650
rect 3200 640 3240 650
rect 4720 640 4800 650
rect 5160 640 5200 650
rect 5280 640 5320 650
rect 5400 640 5440 650
rect 5480 640 5560 650
rect 5680 640 5760 650
rect 6280 640 6360 650
rect 6480 640 6520 650
rect 7400 640 7440 650
rect 8160 640 8320 650
rect 8720 640 9120 650
rect 0 630 480 640
rect 1280 630 1360 640
rect 2080 630 2120 640
rect 3200 630 3240 640
rect 4720 630 4800 640
rect 5160 630 5200 640
rect 5280 630 5320 640
rect 5400 630 5440 640
rect 5480 630 5560 640
rect 5680 630 5760 640
rect 6280 630 6360 640
rect 6480 630 6520 640
rect 7400 630 7440 640
rect 8160 630 8320 640
rect 8720 630 9120 640
rect 0 620 480 630
rect 1280 620 1360 630
rect 2080 620 2120 630
rect 3200 620 3240 630
rect 4720 620 4800 630
rect 5160 620 5200 630
rect 5280 620 5320 630
rect 5400 620 5440 630
rect 5480 620 5560 630
rect 5680 620 5760 630
rect 6280 620 6360 630
rect 6480 620 6520 630
rect 7400 620 7440 630
rect 8160 620 8320 630
rect 8720 620 9120 630
rect 0 610 360 620
rect 1240 610 1320 620
rect 2240 610 2280 620
rect 4720 610 4760 620
rect 5560 610 5600 620
rect 5680 610 5840 620
rect 6320 610 6360 620
rect 6520 610 6560 620
rect 7400 610 7440 620
rect 8000 610 8040 620
rect 8160 610 8360 620
rect 8680 610 9080 620
rect 0 600 360 610
rect 1240 600 1320 610
rect 2240 600 2280 610
rect 4720 600 4760 610
rect 5560 600 5600 610
rect 5680 600 5840 610
rect 6320 600 6360 610
rect 6520 600 6560 610
rect 7400 600 7440 610
rect 8000 600 8040 610
rect 8160 600 8360 610
rect 8680 600 9080 610
rect 0 590 360 600
rect 1240 590 1320 600
rect 2240 590 2280 600
rect 4720 590 4760 600
rect 5560 590 5600 600
rect 5680 590 5840 600
rect 6320 590 6360 600
rect 6520 590 6560 600
rect 7400 590 7440 600
rect 8000 590 8040 600
rect 8160 590 8360 600
rect 8680 590 9080 600
rect 0 580 360 590
rect 1240 580 1320 590
rect 2240 580 2280 590
rect 4720 580 4760 590
rect 5560 580 5600 590
rect 5680 580 5840 590
rect 6320 580 6360 590
rect 6520 580 6560 590
rect 7400 580 7440 590
rect 8000 580 8040 590
rect 8160 580 8360 590
rect 8680 580 9080 590
rect 0 570 320 580
rect 1200 570 1240 580
rect 2120 570 2200 580
rect 4720 570 4760 580
rect 5560 570 5600 580
rect 5680 570 5880 580
rect 6320 570 6360 580
rect 6520 570 6560 580
rect 7360 570 7440 580
rect 8040 570 8080 580
rect 8120 570 8440 580
rect 8560 570 9040 580
rect 0 560 320 570
rect 1200 560 1240 570
rect 2120 560 2200 570
rect 4720 560 4760 570
rect 5560 560 5600 570
rect 5680 560 5880 570
rect 6320 560 6360 570
rect 6520 560 6560 570
rect 7360 560 7440 570
rect 8040 560 8080 570
rect 8120 560 8440 570
rect 8560 560 9040 570
rect 0 550 320 560
rect 1200 550 1240 560
rect 2120 550 2200 560
rect 4720 550 4760 560
rect 5560 550 5600 560
rect 5680 550 5880 560
rect 6320 550 6360 560
rect 6520 550 6560 560
rect 7360 550 7440 560
rect 8040 550 8080 560
rect 8120 550 8440 560
rect 8560 550 9040 560
rect 0 540 320 550
rect 1200 540 1240 550
rect 2120 540 2200 550
rect 4720 540 4760 550
rect 5560 540 5600 550
rect 5680 540 5880 550
rect 6320 540 6360 550
rect 6520 540 6560 550
rect 7360 540 7440 550
rect 8040 540 8080 550
rect 8120 540 8440 550
rect 8560 540 9040 550
rect 0 530 200 540
rect 680 530 720 540
rect 760 530 800 540
rect 840 530 880 540
rect 1080 530 1200 540
rect 2880 530 2920 540
rect 4480 530 4520 540
rect 4680 530 4720 540
rect 5360 530 5480 540
rect 5600 530 5920 540
rect 6320 530 6360 540
rect 6560 530 6600 540
rect 7360 530 7440 540
rect 8080 530 9160 540
rect 0 520 200 530
rect 680 520 720 530
rect 760 520 800 530
rect 840 520 880 530
rect 1080 520 1200 530
rect 2880 520 2920 530
rect 4480 520 4520 530
rect 4680 520 4720 530
rect 5360 520 5480 530
rect 5600 520 5920 530
rect 6320 520 6360 530
rect 6560 520 6600 530
rect 7360 520 7440 530
rect 8080 520 9160 530
rect 0 510 200 520
rect 680 510 720 520
rect 760 510 800 520
rect 840 510 880 520
rect 1080 510 1200 520
rect 2880 510 2920 520
rect 4480 510 4520 520
rect 4680 510 4720 520
rect 5360 510 5480 520
rect 5600 510 5920 520
rect 6320 510 6360 520
rect 6560 510 6600 520
rect 7360 510 7440 520
rect 8080 510 9160 520
rect 0 500 200 510
rect 680 500 720 510
rect 760 500 800 510
rect 840 500 880 510
rect 1080 500 1200 510
rect 2880 500 2920 510
rect 4480 500 4520 510
rect 4680 500 4720 510
rect 5360 500 5480 510
rect 5600 500 5920 510
rect 6320 500 6360 510
rect 6560 500 6600 510
rect 7360 500 7440 510
rect 8080 500 9160 510
rect 0 490 120 500
rect 640 490 920 500
rect 1080 490 1160 500
rect 2120 490 2160 500
rect 2760 490 2800 500
rect 4320 490 4480 500
rect 4520 490 4560 500
rect 4680 490 4720 500
rect 5360 490 5480 500
rect 5680 490 5800 500
rect 5840 490 5920 500
rect 6560 490 6600 500
rect 7360 490 7440 500
rect 8120 490 9080 500
rect 9200 490 9240 500
rect 0 480 120 490
rect 640 480 920 490
rect 1080 480 1160 490
rect 2120 480 2160 490
rect 2760 480 2800 490
rect 4320 480 4480 490
rect 4520 480 4560 490
rect 4680 480 4720 490
rect 5360 480 5480 490
rect 5680 480 5800 490
rect 5840 480 5920 490
rect 6560 480 6600 490
rect 7360 480 7440 490
rect 8120 480 9080 490
rect 9200 480 9240 490
rect 0 470 120 480
rect 640 470 920 480
rect 1080 470 1160 480
rect 2120 470 2160 480
rect 2760 470 2800 480
rect 4320 470 4480 480
rect 4520 470 4560 480
rect 4680 470 4720 480
rect 5360 470 5480 480
rect 5680 470 5800 480
rect 5840 470 5920 480
rect 6560 470 6600 480
rect 7360 470 7440 480
rect 8120 470 9080 480
rect 9200 470 9240 480
rect 0 460 120 470
rect 640 460 920 470
rect 1080 460 1160 470
rect 2120 460 2160 470
rect 2760 460 2800 470
rect 4320 460 4480 470
rect 4520 460 4560 470
rect 4680 460 4720 470
rect 5360 460 5480 470
rect 5680 460 5800 470
rect 5840 460 5920 470
rect 6560 460 6600 470
rect 7360 460 7440 470
rect 8120 460 9080 470
rect 9200 460 9240 470
rect 0 450 80 460
rect 560 450 600 460
rect 800 450 1120 460
rect 1800 450 1840 460
rect 4280 450 4320 460
rect 4440 450 4560 460
rect 4680 450 4720 460
rect 5680 450 5800 460
rect 5880 450 5960 460
rect 6280 450 6360 460
rect 6600 450 6640 460
rect 7360 450 7440 460
rect 8200 450 9000 460
rect 0 440 80 450
rect 560 440 600 450
rect 800 440 1120 450
rect 1800 440 1840 450
rect 4280 440 4320 450
rect 4440 440 4560 450
rect 4680 440 4720 450
rect 5680 440 5800 450
rect 5880 440 5960 450
rect 6280 440 6360 450
rect 6600 440 6640 450
rect 7360 440 7440 450
rect 8200 440 9000 450
rect 0 430 80 440
rect 560 430 600 440
rect 800 430 1120 440
rect 1800 430 1840 440
rect 4280 430 4320 440
rect 4440 430 4560 440
rect 4680 430 4720 440
rect 5680 430 5800 440
rect 5880 430 5960 440
rect 6280 430 6360 440
rect 6600 430 6640 440
rect 7360 430 7440 440
rect 8200 430 9000 440
rect 0 420 80 430
rect 560 420 600 430
rect 800 420 1120 430
rect 1800 420 1840 430
rect 4280 420 4320 430
rect 4440 420 4560 430
rect 4680 420 4720 430
rect 5680 420 5800 430
rect 5880 420 5960 430
rect 6280 420 6360 430
rect 6600 420 6640 430
rect 7360 420 7440 430
rect 8200 420 9000 430
rect 0 410 80 420
rect 400 410 440 420
rect 760 410 1080 420
rect 4280 410 4320 420
rect 4360 410 4720 420
rect 5200 410 5280 420
rect 5320 410 5360 420
rect 5720 410 6000 420
rect 6280 410 6360 420
rect 6600 410 6680 420
rect 7360 410 7440 420
rect 8280 410 9000 420
rect 9160 410 9200 420
rect 0 400 80 410
rect 400 400 440 410
rect 760 400 1080 410
rect 4280 400 4320 410
rect 4360 400 4720 410
rect 5200 400 5280 410
rect 5320 400 5360 410
rect 5720 400 6000 410
rect 6280 400 6360 410
rect 6600 400 6680 410
rect 7360 400 7440 410
rect 8280 400 9000 410
rect 9160 400 9200 410
rect 0 390 80 400
rect 400 390 440 400
rect 760 390 1080 400
rect 4280 390 4320 400
rect 4360 390 4720 400
rect 5200 390 5280 400
rect 5320 390 5360 400
rect 5720 390 6000 400
rect 6280 390 6360 400
rect 6600 390 6680 400
rect 7360 390 7440 400
rect 8280 390 9000 400
rect 9160 390 9200 400
rect 0 380 80 390
rect 400 380 440 390
rect 760 380 1080 390
rect 4280 380 4320 390
rect 4360 380 4720 390
rect 5200 380 5280 390
rect 5320 380 5360 390
rect 5720 380 6000 390
rect 6280 380 6360 390
rect 6600 380 6680 390
rect 7360 380 7440 390
rect 8280 380 9000 390
rect 9160 380 9200 390
rect 0 370 40 380
rect 400 370 440 380
rect 800 370 840 380
rect 920 370 1040 380
rect 4400 370 4560 380
rect 4600 370 4720 380
rect 5200 370 5280 380
rect 5320 370 5400 380
rect 5760 370 5800 380
rect 5840 370 6000 380
rect 6280 370 6360 380
rect 6640 370 6720 380
rect 7320 370 7440 380
rect 8280 370 8800 380
rect 8840 370 8960 380
rect 9040 370 9080 380
rect 9320 370 9360 380
rect 0 360 40 370
rect 400 360 440 370
rect 800 360 840 370
rect 920 360 1040 370
rect 4400 360 4560 370
rect 4600 360 4720 370
rect 5200 360 5280 370
rect 5320 360 5400 370
rect 5760 360 5800 370
rect 5840 360 6000 370
rect 6280 360 6360 370
rect 6640 360 6720 370
rect 7320 360 7440 370
rect 8280 360 8800 370
rect 8840 360 8960 370
rect 9040 360 9080 370
rect 9320 360 9360 370
rect 0 350 40 360
rect 400 350 440 360
rect 800 350 840 360
rect 920 350 1040 360
rect 4400 350 4560 360
rect 4600 350 4720 360
rect 5200 350 5280 360
rect 5320 350 5400 360
rect 5760 350 5800 360
rect 5840 350 6000 360
rect 6280 350 6360 360
rect 6640 350 6720 360
rect 7320 350 7440 360
rect 8280 350 8800 360
rect 8840 350 8960 360
rect 9040 350 9080 360
rect 9320 350 9360 360
rect 0 340 40 350
rect 400 340 440 350
rect 800 340 840 350
rect 920 340 1040 350
rect 4400 340 4560 350
rect 4600 340 4720 350
rect 5200 340 5280 350
rect 5320 340 5400 350
rect 5760 340 5800 350
rect 5840 340 6000 350
rect 6280 340 6360 350
rect 6640 340 6720 350
rect 7320 340 7440 350
rect 8280 340 8800 350
rect 8840 340 8960 350
rect 9040 340 9080 350
rect 9320 340 9360 350
rect 800 330 840 340
rect 880 330 1040 340
rect 4560 330 4680 340
rect 5720 330 6000 340
rect 6280 330 6360 340
rect 6680 330 6760 340
rect 7320 330 7440 340
rect 8320 330 9040 340
rect 9240 330 9360 340
rect 800 320 840 330
rect 880 320 1040 330
rect 4560 320 4680 330
rect 5720 320 6000 330
rect 6280 320 6360 330
rect 6680 320 6760 330
rect 7320 320 7440 330
rect 8320 320 9040 330
rect 9240 320 9360 330
rect 800 310 840 320
rect 880 310 1040 320
rect 4560 310 4680 320
rect 5720 310 6000 320
rect 6280 310 6360 320
rect 6680 310 6760 320
rect 7320 310 7440 320
rect 8320 310 9040 320
rect 9240 310 9360 320
rect 800 300 840 310
rect 880 300 1040 310
rect 4560 300 4680 310
rect 5720 300 6000 310
rect 6280 300 6360 310
rect 6680 300 6760 310
rect 7320 300 7440 310
rect 8320 300 9040 310
rect 9240 300 9360 310
rect 5720 290 5840 300
rect 5880 290 6000 300
rect 6040 290 6120 300
rect 6280 290 6360 300
rect 6720 290 6800 300
rect 7320 290 7440 300
rect 8360 290 8880 300
rect 8920 290 9040 300
rect 9240 290 9280 300
rect 5720 280 5840 290
rect 5880 280 6000 290
rect 6040 280 6120 290
rect 6280 280 6360 290
rect 6720 280 6800 290
rect 7320 280 7440 290
rect 8360 280 8880 290
rect 8920 280 9040 290
rect 9240 280 9280 290
rect 5720 270 5840 280
rect 5880 270 6000 280
rect 6040 270 6120 280
rect 6280 270 6360 280
rect 6720 270 6800 280
rect 7320 270 7440 280
rect 8360 270 8880 280
rect 8920 270 9040 280
rect 9240 270 9280 280
rect 5720 260 5840 270
rect 5880 260 6000 270
rect 6040 260 6120 270
rect 6280 260 6360 270
rect 6720 260 6800 270
rect 7320 260 7440 270
rect 8360 260 8880 270
rect 8920 260 9040 270
rect 9240 260 9280 270
rect 5720 250 5800 260
rect 5960 250 6120 260
rect 6280 250 6360 260
rect 6720 250 6840 260
rect 7320 250 7400 260
rect 8400 250 8880 260
rect 8960 250 9000 260
rect 5720 240 5800 250
rect 5960 240 6120 250
rect 6280 240 6360 250
rect 6720 240 6840 250
rect 7320 240 7400 250
rect 8400 240 8880 250
rect 8960 240 9000 250
rect 5720 230 5800 240
rect 5960 230 6120 240
rect 6280 230 6360 240
rect 6720 230 6840 240
rect 7320 230 7400 240
rect 8400 230 8880 240
rect 8960 230 9000 240
rect 5720 220 5800 230
rect 5960 220 6120 230
rect 6280 220 6360 230
rect 6720 220 6840 230
rect 7320 220 7400 230
rect 8400 220 8880 230
rect 8960 220 9000 230
rect 160 210 200 220
rect 6000 210 6080 220
rect 6320 210 6360 220
rect 6760 210 6880 220
rect 7320 210 7400 220
rect 8440 210 8600 220
rect 8640 210 8680 220
rect 8720 210 8840 220
rect 8960 210 9000 220
rect 160 200 200 210
rect 6000 200 6080 210
rect 6320 200 6360 210
rect 6760 200 6880 210
rect 7320 200 7400 210
rect 8440 200 8600 210
rect 8640 200 8680 210
rect 8720 200 8840 210
rect 8960 200 9000 210
rect 160 190 200 200
rect 6000 190 6080 200
rect 6320 190 6360 200
rect 6760 190 6880 200
rect 7320 190 7400 200
rect 8440 190 8600 200
rect 8640 190 8680 200
rect 8720 190 8840 200
rect 8960 190 9000 200
rect 160 180 200 190
rect 6000 180 6080 190
rect 6320 180 6360 190
rect 6760 180 6880 190
rect 7320 180 7400 190
rect 8440 180 8600 190
rect 8640 180 8680 190
rect 8720 180 8840 190
rect 8960 180 9000 190
rect 160 170 240 180
rect 360 170 440 180
rect 5360 170 5720 180
rect 5960 170 6080 180
rect 6320 170 6400 180
rect 6800 170 6960 180
rect 7320 170 7400 180
rect 8480 170 8560 180
rect 8760 170 8840 180
rect 9040 170 9080 180
rect 9200 170 9280 180
rect 9800 170 9840 180
rect 160 160 240 170
rect 360 160 440 170
rect 5360 160 5720 170
rect 5960 160 6080 170
rect 6320 160 6400 170
rect 6800 160 6960 170
rect 7320 160 7400 170
rect 8480 160 8560 170
rect 8760 160 8840 170
rect 9040 160 9080 170
rect 9200 160 9280 170
rect 9800 160 9840 170
rect 160 150 240 160
rect 360 150 440 160
rect 5360 150 5720 160
rect 5960 150 6080 160
rect 6320 150 6400 160
rect 6800 150 6960 160
rect 7320 150 7400 160
rect 8480 150 8560 160
rect 8760 150 8840 160
rect 9040 150 9080 160
rect 9200 150 9280 160
rect 9800 150 9840 160
rect 160 140 240 150
rect 360 140 440 150
rect 5360 140 5720 150
rect 5960 140 6080 150
rect 6320 140 6400 150
rect 6800 140 6960 150
rect 7320 140 7400 150
rect 8480 140 8560 150
rect 8760 140 8840 150
rect 9040 140 9080 150
rect 9200 140 9280 150
rect 9800 140 9840 150
rect 160 130 240 140
rect 320 130 400 140
rect 480 130 560 140
rect 4280 130 4440 140
rect 4880 130 4920 140
rect 5320 130 5960 140
rect 6000 130 6080 140
rect 6320 130 6400 140
rect 6800 130 7000 140
rect 7320 130 7400 140
rect 8520 130 8560 140
rect 8720 130 8800 140
rect 9040 130 9080 140
rect 9200 130 9320 140
rect 9760 130 9880 140
rect 160 120 240 130
rect 320 120 400 130
rect 480 120 560 130
rect 4280 120 4440 130
rect 4880 120 4920 130
rect 5320 120 5960 130
rect 6000 120 6080 130
rect 6320 120 6400 130
rect 6800 120 7000 130
rect 7320 120 7400 130
rect 8520 120 8560 130
rect 8720 120 8800 130
rect 9040 120 9080 130
rect 9200 120 9320 130
rect 9760 120 9880 130
rect 160 110 240 120
rect 320 110 400 120
rect 480 110 560 120
rect 4280 110 4440 120
rect 4880 110 4920 120
rect 5320 110 5960 120
rect 6000 110 6080 120
rect 6320 110 6400 120
rect 6800 110 7000 120
rect 7320 110 7400 120
rect 8520 110 8560 120
rect 8720 110 8800 120
rect 9040 110 9080 120
rect 9200 110 9320 120
rect 9760 110 9880 120
rect 160 100 240 110
rect 320 100 400 110
rect 480 100 560 110
rect 4280 100 4440 110
rect 4880 100 4920 110
rect 5320 100 5960 110
rect 6000 100 6080 110
rect 6320 100 6400 110
rect 6800 100 7000 110
rect 7320 100 7400 110
rect 8520 100 8560 110
rect 8720 100 8800 110
rect 9040 100 9080 110
rect 9200 100 9320 110
rect 9760 100 9880 110
rect 160 90 280 100
rect 320 90 360 100
rect 520 90 640 100
rect 680 90 840 100
rect 4320 90 4520 100
rect 4840 90 4880 100
rect 5360 90 5880 100
rect 6000 90 6080 100
rect 6400 90 6440 100
rect 6840 90 7040 100
rect 7320 90 7400 100
rect 8560 90 8600 100
rect 8720 90 8760 100
rect 8960 90 9000 100
rect 9200 90 9280 100
rect 9320 90 9360 100
rect 9800 90 9880 100
rect 160 80 280 90
rect 320 80 360 90
rect 520 80 640 90
rect 680 80 840 90
rect 4320 80 4520 90
rect 4840 80 4880 90
rect 5360 80 5880 90
rect 6000 80 6080 90
rect 6400 80 6440 90
rect 6840 80 7040 90
rect 7320 80 7400 90
rect 8560 80 8600 90
rect 8720 80 8760 90
rect 8960 80 9000 90
rect 9200 80 9280 90
rect 9320 80 9360 90
rect 9800 80 9880 90
rect 160 70 280 80
rect 320 70 360 80
rect 520 70 640 80
rect 680 70 840 80
rect 4320 70 4520 80
rect 4840 70 4880 80
rect 5360 70 5880 80
rect 6000 70 6080 80
rect 6400 70 6440 80
rect 6840 70 7040 80
rect 7320 70 7400 80
rect 8560 70 8600 80
rect 8720 70 8760 80
rect 8960 70 9000 80
rect 9200 70 9280 80
rect 9320 70 9360 80
rect 9800 70 9880 80
rect 160 60 280 70
rect 320 60 360 70
rect 520 60 640 70
rect 680 60 840 70
rect 4320 60 4520 70
rect 4840 60 4880 70
rect 5360 60 5880 70
rect 6000 60 6080 70
rect 6400 60 6440 70
rect 6840 60 7040 70
rect 7320 60 7400 70
rect 8560 60 8600 70
rect 8720 60 8760 70
rect 8960 60 9000 70
rect 9200 60 9280 70
rect 9320 60 9360 70
rect 9800 60 9880 70
rect 160 50 280 60
rect 320 50 360 60
rect 600 50 880 60
rect 4360 50 4520 60
rect 4560 50 4600 60
rect 4800 50 4840 60
rect 5360 50 5680 60
rect 5800 50 6080 60
rect 6440 50 6480 60
rect 6840 50 7120 60
rect 7320 50 7360 60
rect 8600 50 8720 60
rect 9200 50 9240 60
rect 9360 50 9440 60
rect 9800 50 9880 60
rect 160 40 280 50
rect 320 40 360 50
rect 600 40 880 50
rect 4360 40 4520 50
rect 4560 40 4600 50
rect 4800 40 4840 50
rect 5360 40 5680 50
rect 5800 40 6080 50
rect 6440 40 6480 50
rect 6840 40 7120 50
rect 7320 40 7360 50
rect 8600 40 8720 50
rect 9200 40 9240 50
rect 9360 40 9440 50
rect 9800 40 9880 50
rect 160 30 280 40
rect 320 30 360 40
rect 600 30 880 40
rect 4360 30 4520 40
rect 4560 30 4600 40
rect 4800 30 4840 40
rect 5360 30 5680 40
rect 5800 30 6080 40
rect 6440 30 6480 40
rect 6840 30 7120 40
rect 7320 30 7360 40
rect 8600 30 8720 40
rect 9200 30 9240 40
rect 9360 30 9440 40
rect 9800 30 9880 40
rect 160 20 280 30
rect 320 20 360 30
rect 600 20 880 30
rect 4360 20 4520 30
rect 4560 20 4600 30
rect 4800 20 4840 30
rect 5360 20 5680 30
rect 5800 20 6080 30
rect 6440 20 6480 30
rect 6840 20 7120 30
rect 7320 20 7360 30
rect 8600 20 8720 30
rect 9200 20 9240 30
rect 9360 20 9440 30
rect 9800 20 9880 30
rect 160 10 240 20
rect 320 10 360 20
rect 600 10 680 20
rect 720 10 920 20
rect 4400 10 4600 20
rect 5400 10 5640 20
rect 5840 10 6080 20
rect 6440 10 6480 20
rect 6880 10 7160 20
rect 7280 10 7360 20
rect 8680 10 8720 20
rect 9200 10 9240 20
rect 9400 10 9440 20
rect 9800 10 9920 20
rect 160 0 240 10
rect 320 0 360 10
rect 600 0 680 10
rect 720 0 920 10
rect 4400 0 4600 10
rect 5400 0 5640 10
rect 5840 0 6080 10
rect 6440 0 6480 10
rect 6880 0 7160 10
rect 7280 0 7360 10
rect 8680 0 8720 10
rect 9200 0 9240 10
rect 9400 0 9440 10
rect 9800 0 9920 10
<< metal2 >>
rect 2160 7490 2200 7500
rect 9760 7490 9800 7500
rect 2160 7480 2200 7490
rect 9760 7480 9800 7490
rect 2160 7470 2200 7480
rect 9760 7470 9800 7480
rect 2160 7460 2200 7470
rect 9760 7460 9800 7470
rect 2120 7450 2160 7460
rect 3560 7450 3600 7460
rect 9640 7450 9760 7460
rect 9960 7450 9990 7460
rect 2120 7440 2160 7450
rect 3560 7440 3600 7450
rect 9640 7440 9760 7450
rect 9960 7440 9990 7450
rect 2120 7430 2160 7440
rect 3560 7430 3600 7440
rect 9640 7430 9760 7440
rect 9960 7430 9990 7440
rect 2120 7420 2160 7430
rect 3560 7420 3600 7430
rect 9640 7420 9760 7430
rect 9960 7420 9990 7430
rect 2080 7410 2120 7420
rect 3600 7410 3640 7420
rect 9640 7410 9680 7420
rect 9920 7410 9990 7420
rect 2080 7400 2120 7410
rect 3600 7400 3640 7410
rect 9640 7400 9680 7410
rect 9920 7400 9990 7410
rect 2080 7390 2120 7400
rect 3600 7390 3640 7400
rect 9640 7390 9680 7400
rect 9920 7390 9990 7400
rect 2080 7380 2120 7390
rect 3600 7380 3640 7390
rect 9640 7380 9680 7390
rect 9920 7380 9990 7390
rect 2040 7370 2080 7380
rect 3320 7370 3360 7380
rect 2040 7360 2080 7370
rect 3320 7360 3360 7370
rect 2040 7350 2080 7360
rect 3320 7350 3360 7360
rect 2040 7340 2080 7350
rect 3320 7340 3360 7350
rect 9960 7330 9990 7340
rect 9960 7320 9990 7330
rect 9960 7310 9990 7320
rect 9960 7300 9990 7310
rect 2000 7290 2040 7300
rect 9640 7290 9840 7300
rect 9960 7290 9990 7300
rect 2000 7280 2040 7290
rect 9640 7280 9840 7290
rect 9960 7280 9990 7290
rect 2000 7270 2040 7280
rect 9640 7270 9840 7280
rect 9960 7270 9990 7280
rect 2000 7260 2040 7270
rect 9640 7260 9840 7270
rect 9960 7260 9990 7270
rect 3360 7250 3440 7260
rect 3840 7250 3880 7260
rect 9640 7250 9880 7260
rect 9960 7250 9990 7260
rect 3360 7240 3440 7250
rect 3840 7240 3880 7250
rect 9640 7240 9880 7250
rect 9960 7240 9990 7250
rect 3360 7230 3440 7240
rect 3840 7230 3880 7240
rect 9640 7230 9880 7240
rect 9960 7230 9990 7240
rect 3360 7220 3440 7230
rect 3840 7220 3880 7230
rect 9640 7220 9880 7230
rect 9960 7220 9990 7230
rect 1960 7210 2000 7220
rect 3880 7210 3920 7220
rect 9600 7210 9840 7220
rect 9960 7210 9990 7220
rect 1960 7200 2000 7210
rect 3880 7200 3920 7210
rect 9600 7200 9840 7210
rect 9960 7200 9990 7210
rect 1960 7190 2000 7200
rect 3880 7190 3920 7200
rect 9600 7190 9840 7200
rect 9960 7190 9990 7200
rect 1960 7180 2000 7190
rect 3880 7180 3920 7190
rect 9600 7180 9840 7190
rect 9960 7180 9990 7190
rect 1920 7170 1960 7180
rect 3880 7170 3920 7180
rect 9600 7170 9840 7180
rect 1920 7160 1960 7170
rect 3880 7160 3920 7170
rect 9600 7160 9840 7170
rect 1920 7150 1960 7160
rect 3880 7150 3920 7160
rect 9600 7150 9840 7160
rect 1920 7140 1960 7150
rect 3880 7140 3920 7150
rect 9600 7140 9840 7150
rect 1920 7130 1960 7140
rect 3400 7130 3440 7140
rect 3520 7130 3560 7140
rect 3640 7130 3720 7140
rect 3880 7130 3920 7140
rect 9600 7130 9680 7140
rect 9720 7130 9840 7140
rect 1920 7120 1960 7130
rect 3400 7120 3440 7130
rect 3520 7120 3560 7130
rect 3640 7120 3720 7130
rect 3880 7120 3920 7130
rect 9600 7120 9680 7130
rect 9720 7120 9840 7130
rect 1920 7110 1960 7120
rect 3400 7110 3440 7120
rect 3520 7110 3560 7120
rect 3640 7110 3720 7120
rect 3880 7110 3920 7120
rect 9600 7110 9680 7120
rect 9720 7110 9840 7120
rect 1920 7100 1960 7110
rect 3400 7100 3440 7110
rect 3520 7100 3560 7110
rect 3640 7100 3720 7110
rect 3880 7100 3920 7110
rect 9600 7100 9680 7110
rect 9720 7100 9840 7110
rect 2040 7090 2120 7100
rect 3480 7090 3520 7100
rect 3680 7090 3800 7100
rect 3840 7090 3920 7100
rect 9560 7090 9680 7100
rect 9720 7090 9800 7100
rect 2040 7080 2120 7090
rect 3480 7080 3520 7090
rect 3680 7080 3800 7090
rect 3840 7080 3920 7090
rect 9560 7080 9680 7090
rect 9720 7080 9800 7090
rect 2040 7070 2120 7080
rect 3480 7070 3520 7080
rect 3680 7070 3800 7080
rect 3840 7070 3920 7080
rect 9560 7070 9680 7080
rect 9720 7070 9800 7080
rect 2040 7060 2120 7070
rect 3480 7060 3520 7070
rect 3680 7060 3800 7070
rect 3840 7060 3920 7070
rect 9560 7060 9680 7070
rect 9720 7060 9800 7070
rect 1920 7050 1960 7060
rect 2000 7050 2080 7060
rect 3680 7050 3720 7060
rect 3840 7050 3920 7060
rect 9600 7050 9680 7060
rect 1920 7040 1960 7050
rect 2000 7040 2080 7050
rect 3680 7040 3720 7050
rect 3840 7040 3920 7050
rect 9600 7040 9680 7050
rect 1920 7030 1960 7040
rect 2000 7030 2080 7040
rect 3680 7030 3720 7040
rect 3840 7030 3920 7040
rect 9600 7030 9680 7040
rect 1920 7020 1960 7030
rect 2000 7020 2080 7030
rect 3680 7020 3720 7030
rect 3840 7020 3920 7030
rect 9600 7020 9680 7030
rect 1960 7010 2000 7020
rect 2240 7010 2440 7020
rect 2720 7010 3200 7020
rect 3560 7010 3600 7020
rect 3680 7010 3720 7020
rect 3840 7010 3920 7020
rect 9600 7010 9680 7020
rect 1960 7000 2000 7010
rect 2240 7000 2440 7010
rect 2720 7000 3200 7010
rect 3560 7000 3600 7010
rect 3680 7000 3720 7010
rect 3840 7000 3920 7010
rect 9600 7000 9680 7010
rect 1960 6990 2000 7000
rect 2240 6990 2440 7000
rect 2720 6990 3200 7000
rect 3560 6990 3600 7000
rect 3680 6990 3720 7000
rect 3840 6990 3920 7000
rect 9600 6990 9680 7000
rect 1960 6980 2000 6990
rect 2240 6980 2440 6990
rect 2720 6980 3200 6990
rect 3560 6980 3600 6990
rect 3680 6980 3720 6990
rect 3840 6980 3920 6990
rect 9600 6980 9680 6990
rect 1960 6970 2000 6980
rect 2280 6970 3160 6980
rect 3280 6970 3320 6980
rect 3640 6970 3680 6980
rect 3840 6970 3920 6980
rect 1960 6960 2000 6970
rect 2280 6960 3160 6970
rect 3280 6960 3320 6970
rect 3640 6960 3680 6970
rect 3840 6960 3920 6970
rect 1960 6950 2000 6960
rect 2280 6950 3160 6960
rect 3280 6950 3320 6960
rect 3640 6950 3680 6960
rect 3840 6950 3920 6960
rect 1960 6940 2000 6950
rect 2280 6940 3160 6950
rect 3280 6940 3320 6950
rect 3640 6940 3680 6950
rect 3840 6940 3920 6950
rect 2320 6930 2480 6940
rect 2560 6930 3200 6940
rect 3720 6930 3800 6940
rect 9600 6930 9680 6940
rect 2320 6920 2480 6930
rect 2560 6920 3200 6930
rect 3720 6920 3800 6930
rect 9600 6920 9680 6930
rect 2320 6910 2480 6920
rect 2560 6910 3200 6920
rect 3720 6910 3800 6920
rect 9600 6910 9680 6920
rect 2320 6900 2480 6910
rect 2560 6900 3200 6910
rect 3720 6900 3800 6910
rect 9600 6900 9680 6910
rect 1880 6890 1920 6900
rect 2400 6890 2520 6900
rect 2640 6890 2920 6900
rect 2960 6890 3080 6900
rect 3120 6890 3160 6900
rect 3760 6890 3880 6900
rect 9600 6890 9680 6900
rect 1880 6880 1920 6890
rect 2400 6880 2520 6890
rect 2640 6880 2920 6890
rect 2960 6880 3080 6890
rect 3120 6880 3160 6890
rect 3760 6880 3880 6890
rect 9600 6880 9680 6890
rect 1880 6870 1920 6880
rect 2400 6870 2520 6880
rect 2640 6870 2920 6880
rect 2960 6870 3080 6880
rect 3120 6870 3160 6880
rect 3760 6870 3880 6880
rect 9600 6870 9680 6880
rect 1880 6860 1920 6870
rect 2400 6860 2520 6870
rect 2640 6860 2920 6870
rect 2960 6860 3080 6870
rect 3120 6860 3160 6870
rect 3760 6860 3880 6870
rect 9600 6860 9680 6870
rect 1880 6850 1920 6860
rect 2480 6850 2560 6860
rect 2800 6850 3040 6860
rect 3800 6850 3880 6860
rect 9600 6850 9680 6860
rect 1880 6840 1920 6850
rect 2480 6840 2560 6850
rect 2800 6840 3040 6850
rect 3800 6840 3880 6850
rect 9600 6840 9680 6850
rect 1880 6830 1920 6840
rect 2480 6830 2560 6840
rect 2800 6830 3040 6840
rect 3800 6830 3880 6840
rect 9600 6830 9680 6840
rect 1880 6820 1920 6830
rect 2480 6820 2560 6830
rect 2800 6820 3040 6830
rect 3800 6820 3880 6830
rect 9600 6820 9680 6830
rect 2560 6810 2760 6820
rect 3640 6810 3680 6820
rect 3840 6810 3880 6820
rect 9600 6810 9680 6820
rect 2560 6800 2760 6810
rect 3640 6800 3680 6810
rect 3840 6800 3880 6810
rect 9600 6800 9680 6810
rect 2560 6790 2760 6800
rect 3640 6790 3680 6800
rect 3840 6790 3880 6800
rect 9600 6790 9680 6800
rect 2560 6780 2760 6790
rect 3640 6780 3680 6790
rect 3840 6780 3880 6790
rect 9600 6780 9680 6790
rect 1960 6770 2000 6780
rect 2280 6770 2440 6780
rect 2840 6770 3040 6780
rect 3840 6770 3920 6780
rect 9640 6770 9680 6780
rect 1960 6760 2000 6770
rect 2280 6760 2440 6770
rect 2840 6760 3040 6770
rect 3840 6760 3920 6770
rect 9640 6760 9680 6770
rect 1960 6750 2000 6760
rect 2280 6750 2440 6760
rect 2840 6750 3040 6760
rect 3840 6750 3920 6760
rect 9640 6750 9680 6760
rect 1960 6740 2000 6750
rect 2280 6740 2440 6750
rect 2840 6740 3040 6750
rect 3840 6740 3920 6750
rect 9640 6740 9680 6750
rect 2240 6730 2280 6740
rect 2480 6730 2520 6740
rect 3160 6730 3280 6740
rect 3760 6730 3800 6740
rect 3880 6730 3920 6740
rect 9640 6730 9680 6740
rect 2240 6720 2280 6730
rect 2480 6720 2520 6730
rect 3160 6720 3280 6730
rect 3760 6720 3800 6730
rect 3880 6720 3920 6730
rect 9640 6720 9680 6730
rect 2240 6710 2280 6720
rect 2480 6710 2520 6720
rect 3160 6710 3280 6720
rect 3760 6710 3800 6720
rect 3880 6710 3920 6720
rect 9640 6710 9680 6720
rect 2240 6700 2280 6710
rect 2480 6700 2520 6710
rect 3160 6700 3280 6710
rect 3760 6700 3800 6710
rect 3880 6700 3920 6710
rect 9640 6700 9680 6710
rect 2520 6690 2560 6700
rect 3400 6690 3440 6700
rect 3800 6690 3840 6700
rect 3920 6690 3960 6700
rect 9520 6690 9560 6700
rect 9640 6690 9680 6700
rect 9920 6690 9960 6700
rect 2520 6680 2560 6690
rect 3400 6680 3440 6690
rect 3800 6680 3840 6690
rect 3920 6680 3960 6690
rect 9520 6680 9560 6690
rect 9640 6680 9680 6690
rect 9920 6680 9960 6690
rect 2520 6670 2560 6680
rect 3400 6670 3440 6680
rect 3800 6670 3840 6680
rect 3920 6670 3960 6680
rect 9520 6670 9560 6680
rect 9640 6670 9680 6680
rect 9920 6670 9960 6680
rect 2520 6660 2560 6670
rect 3400 6660 3440 6670
rect 3800 6660 3840 6670
rect 3920 6660 3960 6670
rect 9520 6660 9560 6670
rect 9640 6660 9680 6670
rect 9920 6660 9960 6670
rect 2200 6650 2240 6660
rect 2560 6650 2600 6660
rect 3520 6650 3560 6660
rect 3920 6650 3960 6660
rect 9600 6650 9680 6660
rect 2200 6640 2240 6650
rect 2560 6640 2600 6650
rect 3520 6640 3560 6650
rect 3920 6640 3960 6650
rect 9600 6640 9680 6650
rect 2200 6630 2240 6640
rect 2560 6630 2600 6640
rect 3520 6630 3560 6640
rect 3920 6630 3960 6640
rect 9600 6630 9680 6640
rect 2200 6620 2240 6630
rect 2560 6620 2600 6630
rect 3520 6620 3560 6630
rect 3920 6620 3960 6630
rect 9600 6620 9680 6630
rect 1600 6610 1640 6620
rect 2160 6610 2200 6620
rect 2600 6610 2640 6620
rect 3640 6610 3680 6620
rect 9480 6610 9520 6620
rect 9640 6610 9680 6620
rect 1600 6600 1640 6610
rect 2160 6600 2200 6610
rect 2600 6600 2640 6610
rect 3640 6600 3680 6610
rect 9480 6600 9520 6610
rect 9640 6600 9680 6610
rect 1600 6590 1640 6600
rect 2160 6590 2200 6600
rect 2600 6590 2640 6600
rect 3640 6590 3680 6600
rect 9480 6590 9520 6600
rect 9640 6590 9680 6600
rect 1600 6580 1640 6590
rect 2160 6580 2200 6590
rect 2600 6580 2640 6590
rect 3640 6580 3680 6590
rect 9480 6580 9520 6590
rect 9640 6580 9680 6590
rect 1520 6570 1560 6580
rect 1600 6570 1640 6580
rect 2040 6570 2080 6580
rect 2600 6570 2640 6580
rect 3720 6570 3760 6580
rect 3920 6570 4000 6580
rect 1520 6560 1560 6570
rect 1600 6560 1640 6570
rect 2040 6560 2080 6570
rect 2600 6560 2640 6570
rect 3720 6560 3760 6570
rect 3920 6560 4000 6570
rect 1520 6550 1560 6560
rect 1600 6550 1640 6560
rect 2040 6550 2080 6560
rect 2600 6550 2640 6560
rect 3720 6550 3760 6560
rect 3920 6550 4000 6560
rect 1520 6540 1560 6550
rect 1600 6540 1640 6550
rect 2040 6540 2080 6550
rect 2600 6540 2640 6550
rect 3720 6540 3760 6550
rect 3920 6540 4000 6550
rect 1360 6530 1440 6540
rect 1760 6530 1840 6540
rect 2040 6530 2080 6540
rect 2560 6530 2600 6540
rect 3800 6530 3840 6540
rect 6320 6530 6560 6540
rect 1360 6520 1440 6530
rect 1760 6520 1840 6530
rect 2040 6520 2080 6530
rect 2560 6520 2600 6530
rect 3800 6520 3840 6530
rect 6320 6520 6560 6530
rect 1360 6510 1440 6520
rect 1760 6510 1840 6520
rect 2040 6510 2080 6520
rect 2560 6510 2600 6520
rect 3800 6510 3840 6520
rect 6320 6510 6560 6520
rect 1360 6500 1440 6510
rect 1760 6500 1840 6510
rect 2040 6500 2080 6510
rect 2560 6500 2600 6510
rect 3800 6500 3840 6510
rect 6320 6500 6560 6510
rect 1320 6490 1360 6500
rect 1680 6490 1760 6500
rect 1800 6490 1840 6500
rect 2520 6490 2560 6500
rect 3880 6490 3920 6500
rect 6080 6490 6400 6500
rect 6520 6490 6600 6500
rect 1320 6480 1360 6490
rect 1680 6480 1760 6490
rect 1800 6480 1840 6490
rect 2520 6480 2560 6490
rect 3880 6480 3920 6490
rect 6080 6480 6400 6490
rect 6520 6480 6600 6490
rect 1320 6470 1360 6480
rect 1680 6470 1760 6480
rect 1800 6470 1840 6480
rect 2520 6470 2560 6480
rect 3880 6470 3920 6480
rect 6080 6470 6400 6480
rect 6520 6470 6600 6480
rect 1320 6460 1360 6470
rect 1680 6460 1760 6470
rect 1800 6460 1840 6470
rect 2520 6460 2560 6470
rect 3880 6460 3920 6470
rect 6080 6460 6400 6470
rect 6520 6460 6600 6470
rect 1280 6450 1320 6460
rect 1640 6450 1680 6460
rect 1760 6450 1960 6460
rect 2080 6450 2120 6460
rect 6080 6450 6120 6460
rect 6200 6450 6400 6460
rect 6560 6450 6600 6460
rect 9680 6450 9760 6460
rect 1280 6440 1320 6450
rect 1640 6440 1680 6450
rect 1760 6440 1960 6450
rect 2080 6440 2120 6450
rect 6080 6440 6120 6450
rect 6200 6440 6400 6450
rect 6560 6440 6600 6450
rect 9680 6440 9760 6450
rect 1280 6430 1320 6440
rect 1640 6430 1680 6440
rect 1760 6430 1960 6440
rect 2080 6430 2120 6440
rect 6080 6430 6120 6440
rect 6200 6430 6400 6440
rect 6560 6430 6600 6440
rect 9680 6430 9760 6440
rect 1280 6420 1320 6430
rect 1640 6420 1680 6430
rect 1760 6420 1960 6430
rect 2080 6420 2120 6430
rect 6080 6420 6120 6430
rect 6200 6420 6400 6430
rect 6560 6420 6600 6430
rect 9680 6420 9760 6430
rect 1360 6410 1480 6420
rect 1600 6410 1640 6420
rect 1960 6410 2040 6420
rect 4000 6410 4040 6420
rect 6120 6410 6400 6420
rect 6600 6410 6720 6420
rect 9920 6410 9990 6420
rect 1360 6400 1480 6410
rect 1600 6400 1640 6410
rect 1960 6400 2040 6410
rect 4000 6400 4040 6410
rect 6120 6400 6400 6410
rect 6600 6400 6720 6410
rect 9920 6400 9990 6410
rect 1360 6390 1480 6400
rect 1600 6390 1640 6400
rect 1960 6390 2040 6400
rect 4000 6390 4040 6400
rect 6120 6390 6400 6400
rect 6600 6390 6720 6400
rect 9920 6390 9990 6400
rect 1360 6380 1480 6390
rect 1600 6380 1640 6390
rect 1960 6380 2040 6390
rect 4000 6380 4040 6390
rect 6120 6380 6400 6390
rect 6600 6380 6720 6390
rect 9920 6380 9990 6390
rect 1400 6370 1440 6380
rect 5800 6370 5840 6380
rect 6360 6370 6440 6380
rect 6600 6370 6800 6380
rect 1400 6360 1440 6370
rect 5800 6360 5840 6370
rect 6360 6360 6440 6370
rect 6600 6360 6800 6370
rect 1400 6350 1440 6360
rect 5800 6350 5840 6360
rect 6360 6350 6440 6360
rect 6600 6350 6800 6360
rect 1400 6340 1440 6350
rect 5800 6340 5840 6350
rect 6360 6340 6440 6350
rect 6600 6340 6800 6350
rect 1400 6330 1440 6340
rect 1560 6330 1600 6340
rect 1640 6330 1680 6340
rect 2400 6330 2480 6340
rect 5480 6330 5640 6340
rect 5680 6330 5800 6340
rect 6440 6330 6520 6340
rect 6720 6330 6800 6340
rect 1400 6320 1440 6330
rect 1560 6320 1600 6330
rect 1640 6320 1680 6330
rect 2400 6320 2480 6330
rect 5480 6320 5640 6330
rect 5680 6320 5800 6330
rect 6440 6320 6520 6330
rect 6720 6320 6800 6330
rect 1400 6310 1440 6320
rect 1560 6310 1600 6320
rect 1640 6310 1680 6320
rect 2400 6310 2480 6320
rect 5480 6310 5640 6320
rect 5680 6310 5800 6320
rect 6440 6310 6520 6320
rect 6720 6310 6800 6320
rect 1400 6300 1440 6310
rect 1560 6300 1600 6310
rect 1640 6300 1680 6310
rect 2400 6300 2480 6310
rect 5480 6300 5640 6310
rect 5680 6300 5800 6310
rect 6440 6300 6520 6310
rect 6720 6300 6800 6310
rect 1240 6290 1280 6300
rect 1400 6290 1440 6300
rect 1560 6290 1640 6300
rect 1800 6290 1840 6300
rect 2400 6290 2480 6300
rect 5360 6290 5400 6300
rect 5520 6290 5640 6300
rect 6520 6290 6600 6300
rect 6760 6290 6800 6300
rect 9840 6290 9960 6300
rect 1240 6280 1280 6290
rect 1400 6280 1440 6290
rect 1560 6280 1640 6290
rect 1800 6280 1840 6290
rect 2400 6280 2480 6290
rect 5360 6280 5400 6290
rect 5520 6280 5640 6290
rect 6520 6280 6600 6290
rect 6760 6280 6800 6290
rect 9840 6280 9960 6290
rect 1240 6270 1280 6280
rect 1400 6270 1440 6280
rect 1560 6270 1640 6280
rect 1800 6270 1840 6280
rect 2400 6270 2480 6280
rect 5360 6270 5400 6280
rect 5520 6270 5640 6280
rect 6520 6270 6600 6280
rect 6760 6270 6800 6280
rect 9840 6270 9960 6280
rect 1240 6260 1280 6270
rect 1400 6260 1440 6270
rect 1560 6260 1640 6270
rect 1800 6260 1840 6270
rect 2400 6260 2480 6270
rect 5360 6260 5400 6270
rect 5520 6260 5640 6270
rect 6520 6260 6600 6270
rect 6760 6260 6800 6270
rect 9840 6260 9960 6270
rect 1400 6250 1440 6260
rect 1560 6250 1600 6260
rect 2400 6250 2440 6260
rect 5320 6250 5360 6260
rect 5520 6250 5560 6260
rect 6560 6250 6640 6260
rect 6760 6250 6840 6260
rect 9400 6250 9440 6260
rect 9480 6250 9520 6260
rect 9640 6250 9680 6260
rect 1400 6240 1440 6250
rect 1560 6240 1600 6250
rect 2400 6240 2440 6250
rect 5320 6240 5360 6250
rect 5520 6240 5560 6250
rect 6560 6240 6640 6250
rect 6760 6240 6840 6250
rect 9400 6240 9440 6250
rect 9480 6240 9520 6250
rect 9640 6240 9680 6250
rect 1400 6230 1440 6240
rect 1560 6230 1600 6240
rect 2400 6230 2440 6240
rect 5320 6230 5360 6240
rect 5520 6230 5560 6240
rect 6560 6230 6640 6240
rect 6760 6230 6840 6240
rect 9400 6230 9440 6240
rect 9480 6230 9520 6240
rect 9640 6230 9680 6240
rect 1400 6220 1440 6230
rect 1560 6220 1600 6230
rect 2400 6220 2440 6230
rect 5320 6220 5360 6230
rect 5520 6220 5560 6230
rect 6560 6220 6640 6230
rect 6760 6220 6840 6230
rect 9400 6220 9440 6230
rect 9480 6220 9520 6230
rect 9640 6220 9680 6230
rect 1320 6210 1440 6220
rect 1600 6210 1640 6220
rect 1720 6210 1760 6220
rect 2400 6210 2440 6220
rect 5480 6210 5520 6220
rect 6640 6210 6680 6220
rect 6760 6210 6800 6220
rect 6840 6210 6880 6220
rect 9320 6210 9400 6220
rect 1320 6200 1440 6210
rect 1600 6200 1640 6210
rect 1720 6200 1760 6210
rect 2400 6200 2440 6210
rect 5480 6200 5520 6210
rect 6640 6200 6680 6210
rect 6760 6200 6800 6210
rect 6840 6200 6880 6210
rect 9320 6200 9400 6210
rect 1320 6190 1440 6200
rect 1600 6190 1640 6200
rect 1720 6190 1760 6200
rect 2400 6190 2440 6200
rect 5480 6190 5520 6200
rect 6640 6190 6680 6200
rect 6760 6190 6800 6200
rect 6840 6190 6880 6200
rect 9320 6190 9400 6200
rect 1320 6180 1440 6190
rect 1600 6180 1640 6190
rect 1720 6180 1760 6190
rect 2400 6180 2440 6190
rect 5480 6180 5520 6190
rect 6640 6180 6680 6190
rect 6760 6180 6800 6190
rect 6840 6180 6880 6190
rect 9320 6180 9400 6190
rect 1280 6170 1440 6180
rect 1600 6170 1680 6180
rect 1720 6170 1760 6180
rect 2400 6170 2440 6180
rect 5280 6170 5320 6180
rect 6760 6170 6880 6180
rect 9240 6170 9280 6180
rect 9600 6170 9680 6180
rect 9800 6170 9840 6180
rect 1280 6160 1440 6170
rect 1600 6160 1680 6170
rect 1720 6160 1760 6170
rect 2400 6160 2440 6170
rect 5280 6160 5320 6170
rect 6760 6160 6880 6170
rect 9240 6160 9280 6170
rect 9600 6160 9680 6170
rect 9800 6160 9840 6170
rect 1280 6150 1440 6160
rect 1600 6150 1680 6160
rect 1720 6150 1760 6160
rect 2400 6150 2440 6160
rect 5280 6150 5320 6160
rect 6760 6150 6880 6160
rect 9240 6150 9280 6160
rect 9600 6150 9680 6160
rect 9800 6150 9840 6160
rect 1280 6140 1440 6150
rect 1600 6140 1680 6150
rect 1720 6140 1760 6150
rect 2400 6140 2440 6150
rect 5280 6140 5320 6150
rect 6760 6140 6880 6150
rect 9240 6140 9280 6150
rect 9600 6140 9680 6150
rect 9800 6140 9840 6150
rect 1280 6130 1360 6140
rect 1400 6130 1440 6140
rect 3920 6130 3960 6140
rect 6680 6130 6720 6140
rect 6840 6130 6920 6140
rect 9160 6130 9200 6140
rect 9400 6130 9440 6140
rect 1280 6120 1360 6130
rect 1400 6120 1440 6130
rect 3920 6120 3960 6130
rect 6680 6120 6720 6130
rect 6840 6120 6920 6130
rect 9160 6120 9200 6130
rect 9400 6120 9440 6130
rect 1280 6110 1360 6120
rect 1400 6110 1440 6120
rect 3920 6110 3960 6120
rect 6680 6110 6720 6120
rect 6840 6110 6920 6120
rect 9160 6110 9200 6120
rect 9400 6110 9440 6120
rect 1280 6100 1360 6110
rect 1400 6100 1440 6110
rect 3920 6100 3960 6110
rect 6680 6100 6720 6110
rect 6840 6100 6920 6110
rect 9160 6100 9200 6110
rect 9400 6100 9440 6110
rect 1280 6090 1320 6100
rect 1640 6090 1680 6100
rect 1760 6090 1800 6100
rect 2440 6090 2480 6100
rect 3840 6090 3880 6100
rect 3960 6090 4000 6100
rect 5240 6090 5280 6100
rect 5360 6090 5400 6100
rect 6720 6090 6760 6100
rect 6840 6090 6960 6100
rect 9080 6090 9120 6100
rect 9320 6090 9360 6100
rect 9480 6090 9520 6100
rect 1280 6080 1320 6090
rect 1640 6080 1680 6090
rect 1760 6080 1800 6090
rect 2440 6080 2480 6090
rect 3840 6080 3880 6090
rect 3960 6080 4000 6090
rect 5240 6080 5280 6090
rect 5360 6080 5400 6090
rect 6720 6080 6760 6090
rect 6840 6080 6960 6090
rect 9080 6080 9120 6090
rect 9320 6080 9360 6090
rect 9480 6080 9520 6090
rect 1280 6070 1320 6080
rect 1640 6070 1680 6080
rect 1760 6070 1800 6080
rect 2440 6070 2480 6080
rect 3840 6070 3880 6080
rect 3960 6070 4000 6080
rect 5240 6070 5280 6080
rect 5360 6070 5400 6080
rect 6720 6070 6760 6080
rect 6840 6070 6960 6080
rect 9080 6070 9120 6080
rect 9320 6070 9360 6080
rect 9480 6070 9520 6080
rect 1280 6060 1320 6070
rect 1640 6060 1680 6070
rect 1760 6060 1800 6070
rect 2440 6060 2480 6070
rect 3840 6060 3880 6070
rect 3960 6060 4000 6070
rect 5240 6060 5280 6070
rect 5360 6060 5400 6070
rect 6720 6060 6760 6070
rect 6840 6060 6960 6070
rect 9080 6060 9120 6070
rect 9320 6060 9360 6070
rect 9480 6060 9520 6070
rect 1200 6050 1240 6060
rect 1280 6050 1320 6060
rect 1600 6050 1720 6060
rect 3760 6050 3800 6060
rect 4000 6050 4040 6060
rect 6720 6050 6760 6060
rect 6800 6050 6960 6060
rect 8920 6050 9040 6060
rect 9160 6050 9200 6060
rect 9320 6050 9360 6060
rect 9400 6050 9440 6060
rect 9480 6050 9520 6060
rect 9840 6050 9880 6060
rect 1200 6040 1240 6050
rect 1280 6040 1320 6050
rect 1600 6040 1720 6050
rect 3760 6040 3800 6050
rect 4000 6040 4040 6050
rect 6720 6040 6760 6050
rect 6800 6040 6960 6050
rect 8920 6040 9040 6050
rect 9160 6040 9200 6050
rect 9320 6040 9360 6050
rect 9400 6040 9440 6050
rect 9480 6040 9520 6050
rect 9840 6040 9880 6050
rect 1200 6030 1240 6040
rect 1280 6030 1320 6040
rect 1600 6030 1720 6040
rect 3760 6030 3800 6040
rect 4000 6030 4040 6040
rect 6720 6030 6760 6040
rect 6800 6030 6960 6040
rect 8920 6030 9040 6040
rect 9160 6030 9200 6040
rect 9320 6030 9360 6040
rect 9400 6030 9440 6040
rect 9480 6030 9520 6040
rect 9840 6030 9880 6040
rect 1200 6020 1240 6030
rect 1280 6020 1320 6030
rect 1600 6020 1720 6030
rect 3760 6020 3800 6030
rect 4000 6020 4040 6030
rect 6720 6020 6760 6030
rect 6800 6020 6960 6030
rect 8920 6020 9040 6030
rect 9160 6020 9200 6030
rect 9320 6020 9360 6030
rect 9400 6020 9440 6030
rect 9480 6020 9520 6030
rect 9840 6020 9880 6030
rect 840 6010 960 6020
rect 1120 6010 1200 6020
rect 1680 6010 1720 6020
rect 3200 6010 3240 6020
rect 3760 6010 3800 6020
rect 4040 6010 4080 6020
rect 4320 6010 4360 6020
rect 6760 6010 6800 6020
rect 6840 6010 6960 6020
rect 8760 6010 8840 6020
rect 9040 6010 9080 6020
rect 840 6000 960 6010
rect 1120 6000 1200 6010
rect 1680 6000 1720 6010
rect 3200 6000 3240 6010
rect 3760 6000 3800 6010
rect 4040 6000 4080 6010
rect 4320 6000 4360 6010
rect 6760 6000 6800 6010
rect 6840 6000 6960 6010
rect 8760 6000 8840 6010
rect 9040 6000 9080 6010
rect 840 5990 960 6000
rect 1120 5990 1200 6000
rect 1680 5990 1720 6000
rect 3200 5990 3240 6000
rect 3760 5990 3800 6000
rect 4040 5990 4080 6000
rect 4320 5990 4360 6000
rect 6760 5990 6800 6000
rect 6840 5990 6960 6000
rect 8760 5990 8840 6000
rect 9040 5990 9080 6000
rect 840 5980 960 5990
rect 1120 5980 1200 5990
rect 1680 5980 1720 5990
rect 3200 5980 3240 5990
rect 3760 5980 3800 5990
rect 4040 5980 4080 5990
rect 4320 5980 4360 5990
rect 6760 5980 6800 5990
rect 6840 5980 6960 5990
rect 8760 5980 8840 5990
rect 9040 5980 9080 5990
rect 920 5970 1120 5980
rect 1160 5970 1200 5980
rect 1680 5970 1720 5980
rect 2520 5970 2560 5980
rect 3160 5970 3240 5980
rect 4120 5970 4160 5980
rect 4320 5970 4360 5980
rect 5160 5970 5200 5980
rect 5320 5970 5360 5980
rect 6760 5970 6840 5980
rect 6960 5970 7000 5980
rect 8640 5970 8680 5980
rect 9160 5970 9200 5980
rect 9880 5970 9920 5980
rect 920 5960 1120 5970
rect 1160 5960 1200 5970
rect 1680 5960 1720 5970
rect 2520 5960 2560 5970
rect 3160 5960 3240 5970
rect 4120 5960 4160 5970
rect 4320 5960 4360 5970
rect 5160 5960 5200 5970
rect 5320 5960 5360 5970
rect 6760 5960 6840 5970
rect 6960 5960 7000 5970
rect 8640 5960 8680 5970
rect 9160 5960 9200 5970
rect 9880 5960 9920 5970
rect 920 5950 1120 5960
rect 1160 5950 1200 5960
rect 1680 5950 1720 5960
rect 2520 5950 2560 5960
rect 3160 5950 3240 5960
rect 4120 5950 4160 5960
rect 4320 5950 4360 5960
rect 5160 5950 5200 5960
rect 5320 5950 5360 5960
rect 6760 5950 6840 5960
rect 6960 5950 7000 5960
rect 8640 5950 8680 5960
rect 9160 5950 9200 5960
rect 9880 5950 9920 5960
rect 920 5940 1120 5950
rect 1160 5940 1200 5950
rect 1680 5940 1720 5950
rect 2520 5940 2560 5950
rect 3160 5940 3240 5950
rect 4120 5940 4160 5950
rect 4320 5940 4360 5950
rect 5160 5940 5200 5950
rect 5320 5940 5360 5950
rect 6760 5940 6840 5950
rect 6960 5940 7000 5950
rect 8640 5940 8680 5950
rect 9160 5940 9200 5950
rect 9880 5940 9920 5950
rect 720 5930 760 5940
rect 1680 5930 1720 5940
rect 3120 5930 3160 5940
rect 3200 5930 3280 5940
rect 5320 5930 5360 5940
rect 6800 5930 6840 5940
rect 6960 5930 7000 5940
rect 8520 5930 8560 5940
rect 9160 5930 9200 5940
rect 9480 5930 9520 5940
rect 720 5920 760 5930
rect 1680 5920 1720 5930
rect 3120 5920 3160 5930
rect 3200 5920 3280 5930
rect 5320 5920 5360 5930
rect 6800 5920 6840 5930
rect 6960 5920 7000 5930
rect 8520 5920 8560 5930
rect 9160 5920 9200 5930
rect 9480 5920 9520 5930
rect 720 5910 760 5920
rect 1680 5910 1720 5920
rect 3120 5910 3160 5920
rect 3200 5910 3280 5920
rect 5320 5910 5360 5920
rect 6800 5910 6840 5920
rect 6960 5910 7000 5920
rect 8520 5910 8560 5920
rect 9160 5910 9200 5920
rect 9480 5910 9520 5920
rect 720 5900 760 5910
rect 1680 5900 1720 5910
rect 3120 5900 3160 5910
rect 3200 5900 3280 5910
rect 5320 5900 5360 5910
rect 6800 5900 6840 5910
rect 6960 5900 7000 5910
rect 8520 5900 8560 5910
rect 9160 5900 9200 5910
rect 9480 5900 9520 5910
rect 680 5890 800 5900
rect 960 5890 1000 5900
rect 1760 5890 1840 5900
rect 3080 5890 3120 5900
rect 5120 5890 5160 5900
rect 6800 5890 6840 5900
rect 6960 5890 7000 5900
rect 8400 5890 8440 5900
rect 8600 5890 8640 5900
rect 8840 5890 8880 5900
rect 9160 5890 9200 5900
rect 680 5880 800 5890
rect 960 5880 1000 5890
rect 1760 5880 1840 5890
rect 3080 5880 3120 5890
rect 5120 5880 5160 5890
rect 6800 5880 6840 5890
rect 6960 5880 7000 5890
rect 8400 5880 8440 5890
rect 8600 5880 8640 5890
rect 8840 5880 8880 5890
rect 9160 5880 9200 5890
rect 680 5870 800 5880
rect 960 5870 1000 5880
rect 1760 5870 1840 5880
rect 3080 5870 3120 5880
rect 5120 5870 5160 5880
rect 6800 5870 6840 5880
rect 6960 5870 7000 5880
rect 8400 5870 8440 5880
rect 8600 5870 8640 5880
rect 8840 5870 8880 5880
rect 9160 5870 9200 5880
rect 680 5860 800 5870
rect 960 5860 1000 5870
rect 1760 5860 1840 5870
rect 3080 5860 3120 5870
rect 5120 5860 5160 5870
rect 6800 5860 6840 5870
rect 6960 5860 7000 5870
rect 8400 5860 8440 5870
rect 8600 5860 8640 5870
rect 8840 5860 8880 5870
rect 9160 5860 9200 5870
rect 640 5850 680 5860
rect 720 5850 800 5860
rect 880 5850 920 5860
rect 2320 5850 2360 5860
rect 2600 5850 2680 5860
rect 2960 5850 3040 5860
rect 3240 5850 3280 5860
rect 3720 5850 3760 5860
rect 6800 5850 6840 5860
rect 6960 5850 7000 5860
rect 8240 5850 8280 5860
rect 8600 5850 8640 5860
rect 8840 5850 8920 5860
rect 8960 5850 9000 5860
rect 9080 5850 9120 5860
rect 9160 5850 9280 5860
rect 640 5840 680 5850
rect 720 5840 800 5850
rect 880 5840 920 5850
rect 2320 5840 2360 5850
rect 2600 5840 2680 5850
rect 2960 5840 3040 5850
rect 3240 5840 3280 5850
rect 3720 5840 3760 5850
rect 6800 5840 6840 5850
rect 6960 5840 7000 5850
rect 8240 5840 8280 5850
rect 8600 5840 8640 5850
rect 8840 5840 8920 5850
rect 8960 5840 9000 5850
rect 9080 5840 9120 5850
rect 9160 5840 9280 5850
rect 640 5830 680 5840
rect 720 5830 800 5840
rect 880 5830 920 5840
rect 2320 5830 2360 5840
rect 2600 5830 2680 5840
rect 2960 5830 3040 5840
rect 3240 5830 3280 5840
rect 3720 5830 3760 5840
rect 6800 5830 6840 5840
rect 6960 5830 7000 5840
rect 8240 5830 8280 5840
rect 8600 5830 8640 5840
rect 8840 5830 8920 5840
rect 8960 5830 9000 5840
rect 9080 5830 9120 5840
rect 9160 5830 9280 5840
rect 640 5820 680 5830
rect 720 5820 800 5830
rect 880 5820 920 5830
rect 2320 5820 2360 5830
rect 2600 5820 2680 5830
rect 2960 5820 3040 5830
rect 3240 5820 3280 5830
rect 3720 5820 3760 5830
rect 6800 5820 6840 5830
rect 6960 5820 7000 5830
rect 8240 5820 8280 5830
rect 8600 5820 8640 5830
rect 8840 5820 8920 5830
rect 8960 5820 9000 5830
rect 9080 5820 9120 5830
rect 9160 5820 9280 5830
rect 560 5810 600 5820
rect 640 5810 720 5820
rect 800 5810 840 5820
rect 1840 5810 1880 5820
rect 2280 5810 2360 5820
rect 2600 5810 2680 5820
rect 2840 5810 2960 5820
rect 3240 5810 3280 5820
rect 3760 5810 3840 5820
rect 6800 5810 6840 5820
rect 6960 5810 7000 5820
rect 8400 5810 8440 5820
rect 8720 5810 8760 5820
rect 8880 5810 8920 5820
rect 560 5800 600 5810
rect 640 5800 720 5810
rect 800 5800 840 5810
rect 1840 5800 1880 5810
rect 2280 5800 2360 5810
rect 2600 5800 2680 5810
rect 2840 5800 2960 5810
rect 3240 5800 3280 5810
rect 3760 5800 3840 5810
rect 6800 5800 6840 5810
rect 6960 5800 7000 5810
rect 8400 5800 8440 5810
rect 8720 5800 8760 5810
rect 8880 5800 8920 5810
rect 560 5790 600 5800
rect 640 5790 720 5800
rect 800 5790 840 5800
rect 1840 5790 1880 5800
rect 2280 5790 2360 5800
rect 2600 5790 2680 5800
rect 2840 5790 2960 5800
rect 3240 5790 3280 5800
rect 3760 5790 3840 5800
rect 6800 5790 6840 5800
rect 6960 5790 7000 5800
rect 8400 5790 8440 5800
rect 8720 5790 8760 5800
rect 8880 5790 8920 5800
rect 560 5780 600 5790
rect 640 5780 720 5790
rect 800 5780 840 5790
rect 1840 5780 1880 5790
rect 2280 5780 2360 5790
rect 2600 5780 2680 5790
rect 2840 5780 2960 5790
rect 3240 5780 3280 5790
rect 3760 5780 3840 5790
rect 6800 5780 6840 5790
rect 6960 5780 7000 5790
rect 8400 5780 8440 5790
rect 8720 5780 8760 5790
rect 8880 5780 8920 5790
rect 2240 5770 2320 5780
rect 2600 5770 2640 5780
rect 2800 5770 2960 5780
rect 3240 5770 3280 5780
rect 3880 5770 3920 5780
rect 5080 5770 5120 5780
rect 5280 5770 5320 5780
rect 6960 5770 7000 5780
rect 8000 5770 8040 5780
rect 8240 5770 8280 5780
rect 8360 5770 8400 5780
rect 8800 5770 8840 5780
rect 9920 5770 9960 5780
rect 2240 5760 2320 5770
rect 2600 5760 2640 5770
rect 2800 5760 2960 5770
rect 3240 5760 3280 5770
rect 3880 5760 3920 5770
rect 5080 5760 5120 5770
rect 5280 5760 5320 5770
rect 6960 5760 7000 5770
rect 8000 5760 8040 5770
rect 8240 5760 8280 5770
rect 8360 5760 8400 5770
rect 8800 5760 8840 5770
rect 9920 5760 9960 5770
rect 2240 5750 2320 5760
rect 2600 5750 2640 5760
rect 2800 5750 2960 5760
rect 3240 5750 3280 5760
rect 3880 5750 3920 5760
rect 5080 5750 5120 5760
rect 5280 5750 5320 5760
rect 6960 5750 7000 5760
rect 8000 5750 8040 5760
rect 8240 5750 8280 5760
rect 8360 5750 8400 5760
rect 8800 5750 8840 5760
rect 9920 5750 9960 5760
rect 2240 5740 2320 5750
rect 2600 5740 2640 5750
rect 2800 5740 2960 5750
rect 3240 5740 3280 5750
rect 3880 5740 3920 5750
rect 5080 5740 5120 5750
rect 5280 5740 5320 5750
rect 6960 5740 7000 5750
rect 8000 5740 8040 5750
rect 8240 5740 8280 5750
rect 8360 5740 8400 5750
rect 8800 5740 8840 5750
rect 9920 5740 9960 5750
rect 1880 5730 1920 5740
rect 2200 5730 2240 5740
rect 2520 5730 2600 5740
rect 2760 5730 2840 5740
rect 3240 5730 3280 5740
rect 3760 5730 3840 5740
rect 6920 5730 6960 5740
rect 7880 5730 7920 5740
rect 8120 5730 8200 5740
rect 8280 5730 8320 5740
rect 8360 5730 8400 5740
rect 1880 5720 1920 5730
rect 2200 5720 2240 5730
rect 2520 5720 2600 5730
rect 2760 5720 2840 5730
rect 3240 5720 3280 5730
rect 3760 5720 3840 5730
rect 6920 5720 6960 5730
rect 7880 5720 7920 5730
rect 8120 5720 8200 5730
rect 8280 5720 8320 5730
rect 8360 5720 8400 5730
rect 1880 5710 1920 5720
rect 2200 5710 2240 5720
rect 2520 5710 2600 5720
rect 2760 5710 2840 5720
rect 3240 5710 3280 5720
rect 3760 5710 3840 5720
rect 6920 5710 6960 5720
rect 7880 5710 7920 5720
rect 8120 5710 8200 5720
rect 8280 5710 8320 5720
rect 8360 5710 8400 5720
rect 1880 5700 1920 5710
rect 2200 5700 2240 5710
rect 2520 5700 2600 5710
rect 2760 5700 2840 5710
rect 3240 5700 3280 5710
rect 3760 5700 3840 5710
rect 6920 5700 6960 5710
rect 7880 5700 7920 5710
rect 8120 5700 8200 5710
rect 8280 5700 8320 5710
rect 8360 5700 8400 5710
rect 800 5690 840 5700
rect 1080 5690 1160 5700
rect 1880 5690 1920 5700
rect 2200 5690 2280 5700
rect 2480 5690 2560 5700
rect 2680 5690 2800 5700
rect 3240 5690 3280 5700
rect 3720 5690 3760 5700
rect 3880 5690 3920 5700
rect 5080 5690 5120 5700
rect 6840 5690 6880 5700
rect 6920 5690 6960 5700
rect 7720 5690 7760 5700
rect 7800 5690 7920 5700
rect 8000 5690 8120 5700
rect 8280 5690 8320 5700
rect 8440 5690 8480 5700
rect 800 5680 840 5690
rect 1080 5680 1160 5690
rect 1880 5680 1920 5690
rect 2200 5680 2280 5690
rect 2480 5680 2560 5690
rect 2680 5680 2800 5690
rect 3240 5680 3280 5690
rect 3720 5680 3760 5690
rect 3880 5680 3920 5690
rect 5080 5680 5120 5690
rect 6840 5680 6880 5690
rect 6920 5680 6960 5690
rect 7720 5680 7760 5690
rect 7800 5680 7920 5690
rect 8000 5680 8120 5690
rect 8280 5680 8320 5690
rect 8440 5680 8480 5690
rect 800 5670 840 5680
rect 1080 5670 1160 5680
rect 1880 5670 1920 5680
rect 2200 5670 2280 5680
rect 2480 5670 2560 5680
rect 2680 5670 2800 5680
rect 3240 5670 3280 5680
rect 3720 5670 3760 5680
rect 3880 5670 3920 5680
rect 5080 5670 5120 5680
rect 6840 5670 6880 5680
rect 6920 5670 6960 5680
rect 7720 5670 7760 5680
rect 7800 5670 7920 5680
rect 8000 5670 8120 5680
rect 8280 5670 8320 5680
rect 8440 5670 8480 5680
rect 800 5660 840 5670
rect 1080 5660 1160 5670
rect 1880 5660 1920 5670
rect 2200 5660 2280 5670
rect 2480 5660 2560 5670
rect 2680 5660 2800 5670
rect 3240 5660 3280 5670
rect 3720 5660 3760 5670
rect 3880 5660 3920 5670
rect 5080 5660 5120 5670
rect 6840 5660 6880 5670
rect 6920 5660 6960 5670
rect 7720 5660 7760 5670
rect 7800 5660 7920 5670
rect 8000 5660 8120 5670
rect 8280 5660 8320 5670
rect 8440 5660 8480 5670
rect 760 5650 800 5660
rect 1880 5650 1960 5660
rect 2480 5650 2520 5660
rect 2640 5650 2720 5660
rect 3240 5650 3280 5660
rect 3720 5650 3760 5660
rect 3840 5650 3880 5660
rect 6840 5650 6880 5660
rect 7640 5650 7720 5660
rect 7800 5650 7920 5660
rect 8000 5650 8040 5660
rect 8520 5650 8560 5660
rect 9960 5650 9990 5660
rect 760 5640 800 5650
rect 1880 5640 1960 5650
rect 2480 5640 2520 5650
rect 2640 5640 2720 5650
rect 3240 5640 3280 5650
rect 3720 5640 3760 5650
rect 3840 5640 3880 5650
rect 6840 5640 6880 5650
rect 7640 5640 7720 5650
rect 7800 5640 7920 5650
rect 8000 5640 8040 5650
rect 8520 5640 8560 5650
rect 9960 5640 9990 5650
rect 760 5630 800 5640
rect 1880 5630 1960 5640
rect 2480 5630 2520 5640
rect 2640 5630 2720 5640
rect 3240 5630 3280 5640
rect 3720 5630 3760 5640
rect 3840 5630 3880 5640
rect 6840 5630 6880 5640
rect 7640 5630 7720 5640
rect 7800 5630 7920 5640
rect 8000 5630 8040 5640
rect 8520 5630 8560 5640
rect 9960 5630 9990 5640
rect 760 5620 800 5630
rect 1880 5620 1960 5630
rect 2480 5620 2520 5630
rect 2640 5620 2720 5630
rect 3240 5620 3280 5630
rect 3720 5620 3760 5630
rect 3840 5620 3880 5630
rect 6840 5620 6880 5630
rect 7640 5620 7720 5630
rect 7800 5620 7920 5630
rect 8000 5620 8040 5630
rect 8520 5620 8560 5630
rect 9960 5620 9990 5630
rect 1920 5610 1960 5620
rect 2160 5610 2200 5620
rect 2440 5610 2480 5620
rect 2640 5610 2720 5620
rect 3240 5610 3280 5620
rect 3680 5610 3720 5620
rect 3760 5610 3800 5620
rect 5560 5610 5600 5620
rect 5800 5610 5840 5620
rect 7440 5610 7680 5620
rect 7720 5610 7800 5620
rect 7920 5610 7960 5620
rect 8000 5610 8040 5620
rect 8400 5610 8480 5620
rect 8960 5610 9000 5620
rect 9960 5610 9990 5620
rect 1920 5600 1960 5610
rect 2160 5600 2200 5610
rect 2440 5600 2480 5610
rect 2640 5600 2720 5610
rect 3240 5600 3280 5610
rect 3680 5600 3720 5610
rect 3760 5600 3800 5610
rect 5560 5600 5600 5610
rect 5800 5600 5840 5610
rect 7440 5600 7680 5610
rect 7720 5600 7800 5610
rect 7920 5600 7960 5610
rect 8000 5600 8040 5610
rect 8400 5600 8480 5610
rect 8960 5600 9000 5610
rect 9960 5600 9990 5610
rect 1920 5590 1960 5600
rect 2160 5590 2200 5600
rect 2440 5590 2480 5600
rect 2640 5590 2720 5600
rect 3240 5590 3280 5600
rect 3680 5590 3720 5600
rect 3760 5590 3800 5600
rect 5560 5590 5600 5600
rect 5800 5590 5840 5600
rect 7440 5590 7680 5600
rect 7720 5590 7800 5600
rect 7920 5590 7960 5600
rect 8000 5590 8040 5600
rect 8400 5590 8480 5600
rect 8960 5590 9000 5600
rect 9960 5590 9990 5600
rect 1920 5580 1960 5590
rect 2160 5580 2200 5590
rect 2440 5580 2480 5590
rect 2640 5580 2720 5590
rect 3240 5580 3280 5590
rect 3680 5580 3720 5590
rect 3760 5580 3800 5590
rect 5560 5580 5600 5590
rect 5800 5580 5840 5590
rect 7440 5580 7680 5590
rect 7720 5580 7800 5590
rect 7920 5580 7960 5590
rect 8000 5580 8040 5590
rect 8400 5580 8480 5590
rect 8960 5580 9000 5590
rect 9960 5580 9990 5590
rect 640 5570 680 5580
rect 1920 5570 1960 5580
rect 2160 5570 2200 5580
rect 2400 5570 2440 5580
rect 2600 5570 2680 5580
rect 2880 5570 2920 5580
rect 3240 5570 3280 5580
rect 3440 5570 3480 5580
rect 3640 5570 3760 5580
rect 5240 5570 5280 5580
rect 5520 5570 5640 5580
rect 5880 5570 5920 5580
rect 6200 5570 6280 5580
rect 6440 5570 6560 5580
rect 6880 5570 6920 5580
rect 7360 5570 7400 5580
rect 7600 5570 7640 5580
rect 7760 5570 7800 5580
rect 7920 5570 7960 5580
rect 8000 5570 8040 5580
rect 8240 5570 8360 5580
rect 8840 5570 8880 5580
rect 8920 5570 8960 5580
rect 9080 5570 9120 5580
rect 640 5560 680 5570
rect 1920 5560 1960 5570
rect 2160 5560 2200 5570
rect 2400 5560 2440 5570
rect 2600 5560 2680 5570
rect 2880 5560 2920 5570
rect 3240 5560 3280 5570
rect 3440 5560 3480 5570
rect 3640 5560 3760 5570
rect 5240 5560 5280 5570
rect 5520 5560 5640 5570
rect 5880 5560 5920 5570
rect 6200 5560 6280 5570
rect 6440 5560 6560 5570
rect 6880 5560 6920 5570
rect 7360 5560 7400 5570
rect 7600 5560 7640 5570
rect 7760 5560 7800 5570
rect 7920 5560 7960 5570
rect 8000 5560 8040 5570
rect 8240 5560 8360 5570
rect 8840 5560 8880 5570
rect 8920 5560 8960 5570
rect 9080 5560 9120 5570
rect 640 5550 680 5560
rect 1920 5550 1960 5560
rect 2160 5550 2200 5560
rect 2400 5550 2440 5560
rect 2600 5550 2680 5560
rect 2880 5550 2920 5560
rect 3240 5550 3280 5560
rect 3440 5550 3480 5560
rect 3640 5550 3760 5560
rect 5240 5550 5280 5560
rect 5520 5550 5640 5560
rect 5880 5550 5920 5560
rect 6200 5550 6280 5560
rect 6440 5550 6560 5560
rect 6880 5550 6920 5560
rect 7360 5550 7400 5560
rect 7600 5550 7640 5560
rect 7760 5550 7800 5560
rect 7920 5550 7960 5560
rect 8000 5550 8040 5560
rect 8240 5550 8360 5560
rect 8840 5550 8880 5560
rect 8920 5550 8960 5560
rect 9080 5550 9120 5560
rect 640 5540 680 5550
rect 1920 5540 1960 5550
rect 2160 5540 2200 5550
rect 2400 5540 2440 5550
rect 2600 5540 2680 5550
rect 2880 5540 2920 5550
rect 3240 5540 3280 5550
rect 3440 5540 3480 5550
rect 3640 5540 3760 5550
rect 5240 5540 5280 5550
rect 5520 5540 5640 5550
rect 5880 5540 5920 5550
rect 6200 5540 6280 5550
rect 6440 5540 6560 5550
rect 6880 5540 6920 5550
rect 7360 5540 7400 5550
rect 7600 5540 7640 5550
rect 7760 5540 7800 5550
rect 7920 5540 7960 5550
rect 8000 5540 8040 5550
rect 8240 5540 8360 5550
rect 8840 5540 8880 5550
rect 8920 5540 8960 5550
rect 9080 5540 9120 5550
rect 520 5530 640 5540
rect 920 5530 960 5540
rect 2160 5530 2200 5540
rect 2600 5530 2680 5540
rect 2840 5530 3000 5540
rect 3200 5530 3240 5540
rect 5640 5530 5720 5540
rect 5920 5530 5960 5540
rect 6160 5530 6240 5540
rect 6520 5530 6600 5540
rect 6880 5530 6960 5540
rect 7480 5530 7520 5540
rect 7720 5530 7760 5540
rect 7840 5530 7880 5540
rect 8680 5530 8720 5540
rect 8840 5530 8880 5540
rect 8920 5530 8960 5540
rect 9040 5530 9080 5540
rect 520 5520 640 5530
rect 920 5520 960 5530
rect 2160 5520 2200 5530
rect 2600 5520 2680 5530
rect 2840 5520 3000 5530
rect 3200 5520 3240 5530
rect 5640 5520 5720 5530
rect 5920 5520 5960 5530
rect 6160 5520 6240 5530
rect 6520 5520 6600 5530
rect 6880 5520 6960 5530
rect 7480 5520 7520 5530
rect 7720 5520 7760 5530
rect 7840 5520 7880 5530
rect 8680 5520 8720 5530
rect 8840 5520 8880 5530
rect 8920 5520 8960 5530
rect 9040 5520 9080 5530
rect 520 5510 640 5520
rect 920 5510 960 5520
rect 2160 5510 2200 5520
rect 2600 5510 2680 5520
rect 2840 5510 3000 5520
rect 3200 5510 3240 5520
rect 5640 5510 5720 5520
rect 5920 5510 5960 5520
rect 6160 5510 6240 5520
rect 6520 5510 6600 5520
rect 6880 5510 6960 5520
rect 7480 5510 7520 5520
rect 7720 5510 7760 5520
rect 7840 5510 7880 5520
rect 8680 5510 8720 5520
rect 8840 5510 8880 5520
rect 8920 5510 8960 5520
rect 9040 5510 9080 5520
rect 520 5500 640 5510
rect 920 5500 960 5510
rect 2160 5500 2200 5510
rect 2600 5500 2680 5510
rect 2840 5500 3000 5510
rect 3200 5500 3240 5510
rect 5640 5500 5720 5510
rect 5920 5500 5960 5510
rect 6160 5500 6240 5510
rect 6520 5500 6600 5510
rect 6880 5500 6960 5510
rect 7480 5500 7520 5510
rect 7720 5500 7760 5510
rect 7840 5500 7880 5510
rect 8680 5500 8720 5510
rect 8840 5500 8880 5510
rect 8920 5500 8960 5510
rect 9040 5500 9080 5510
rect 1960 5490 2000 5500
rect 2160 5490 2200 5500
rect 2360 5490 2400 5500
rect 2560 5490 2600 5500
rect 2760 5490 3000 5500
rect 3200 5490 3240 5500
rect 5520 5490 5720 5500
rect 5920 5490 5960 5500
rect 6160 5490 6200 5500
rect 6440 5490 6520 5500
rect 6920 5490 6960 5500
rect 7480 5490 7520 5500
rect 8640 5490 8680 5500
rect 8920 5490 8960 5500
rect 9000 5490 9040 5500
rect 1960 5480 2000 5490
rect 2160 5480 2200 5490
rect 2360 5480 2400 5490
rect 2560 5480 2600 5490
rect 2760 5480 3000 5490
rect 3200 5480 3240 5490
rect 5520 5480 5720 5490
rect 5920 5480 5960 5490
rect 6160 5480 6200 5490
rect 6440 5480 6520 5490
rect 6920 5480 6960 5490
rect 7480 5480 7520 5490
rect 8640 5480 8680 5490
rect 8920 5480 8960 5490
rect 9000 5480 9040 5490
rect 1960 5470 2000 5480
rect 2160 5470 2200 5480
rect 2360 5470 2400 5480
rect 2560 5470 2600 5480
rect 2760 5470 3000 5480
rect 3200 5470 3240 5480
rect 5520 5470 5720 5480
rect 5920 5470 5960 5480
rect 6160 5470 6200 5480
rect 6440 5470 6520 5480
rect 6920 5470 6960 5480
rect 7480 5470 7520 5480
rect 8640 5470 8680 5480
rect 8920 5470 8960 5480
rect 9000 5470 9040 5480
rect 1960 5460 2000 5470
rect 2160 5460 2200 5470
rect 2360 5460 2400 5470
rect 2560 5460 2600 5470
rect 2760 5460 3000 5470
rect 3200 5460 3240 5470
rect 5520 5460 5720 5470
rect 5920 5460 5960 5470
rect 6160 5460 6200 5470
rect 6440 5460 6520 5470
rect 6920 5460 6960 5470
rect 7480 5460 7520 5470
rect 8640 5460 8680 5470
rect 8920 5460 8960 5470
rect 9000 5460 9040 5470
rect 440 5450 480 5460
rect 1960 5450 2000 5460
rect 2160 5450 2240 5460
rect 2360 5450 2400 5460
rect 2600 5450 2680 5460
rect 2760 5450 2880 5460
rect 2920 5450 3040 5460
rect 3160 5450 3240 5460
rect 3560 5450 3600 5460
rect 5440 5450 5480 5460
rect 5600 5450 5640 5460
rect 5920 5450 5960 5460
rect 6160 5450 6200 5460
rect 6480 5450 6560 5460
rect 6920 5450 6960 5460
rect 7240 5450 7400 5460
rect 7640 5450 7680 5460
rect 7920 5450 7960 5460
rect 8400 5450 8480 5460
rect 9560 5450 9600 5460
rect 440 5440 480 5450
rect 1960 5440 2000 5450
rect 2160 5440 2240 5450
rect 2360 5440 2400 5450
rect 2600 5440 2680 5450
rect 2760 5440 2880 5450
rect 2920 5440 3040 5450
rect 3160 5440 3240 5450
rect 3560 5440 3600 5450
rect 5440 5440 5480 5450
rect 5600 5440 5640 5450
rect 5920 5440 5960 5450
rect 6160 5440 6200 5450
rect 6480 5440 6560 5450
rect 6920 5440 6960 5450
rect 7240 5440 7400 5450
rect 7640 5440 7680 5450
rect 7920 5440 7960 5450
rect 8400 5440 8480 5450
rect 9560 5440 9600 5450
rect 440 5430 480 5440
rect 1960 5430 2000 5440
rect 2160 5430 2240 5440
rect 2360 5430 2400 5440
rect 2600 5430 2680 5440
rect 2760 5430 2880 5440
rect 2920 5430 3040 5440
rect 3160 5430 3240 5440
rect 3560 5430 3600 5440
rect 5440 5430 5480 5440
rect 5600 5430 5640 5440
rect 5920 5430 5960 5440
rect 6160 5430 6200 5440
rect 6480 5430 6560 5440
rect 6920 5430 6960 5440
rect 7240 5430 7400 5440
rect 7640 5430 7680 5440
rect 7920 5430 7960 5440
rect 8400 5430 8480 5440
rect 9560 5430 9600 5440
rect 440 5420 480 5430
rect 1960 5420 2000 5430
rect 2160 5420 2240 5430
rect 2360 5420 2400 5430
rect 2600 5420 2680 5430
rect 2760 5420 2880 5430
rect 2920 5420 3040 5430
rect 3160 5420 3240 5430
rect 3560 5420 3600 5430
rect 5440 5420 5480 5430
rect 5600 5420 5640 5430
rect 5920 5420 5960 5430
rect 6160 5420 6200 5430
rect 6480 5420 6560 5430
rect 6920 5420 6960 5430
rect 7240 5420 7400 5430
rect 7640 5420 7680 5430
rect 7920 5420 7960 5430
rect 8400 5420 8480 5430
rect 9560 5420 9600 5430
rect 1960 5410 2040 5420
rect 2160 5410 2240 5420
rect 2360 5410 2400 5420
rect 2680 5410 2880 5420
rect 3080 5410 3160 5420
rect 5080 5410 5120 5420
rect 5400 5410 5440 5420
rect 6160 5410 6200 5420
rect 6600 5410 6680 5420
rect 7320 5410 7400 5420
rect 7640 5410 7680 5420
rect 7760 5410 7800 5420
rect 7880 5410 7960 5420
rect 8320 5410 8360 5420
rect 8480 5410 8520 5420
rect 8840 5410 8880 5420
rect 9400 5410 9440 5420
rect 1960 5400 2040 5410
rect 2160 5400 2240 5410
rect 2360 5400 2400 5410
rect 2680 5400 2880 5410
rect 3080 5400 3160 5410
rect 5080 5400 5120 5410
rect 5400 5400 5440 5410
rect 6160 5400 6200 5410
rect 6600 5400 6680 5410
rect 7320 5400 7400 5410
rect 7640 5400 7680 5410
rect 7760 5400 7800 5410
rect 7880 5400 7960 5410
rect 8320 5400 8360 5410
rect 8480 5400 8520 5410
rect 8840 5400 8880 5410
rect 9400 5400 9440 5410
rect 1960 5390 2040 5400
rect 2160 5390 2240 5400
rect 2360 5390 2400 5400
rect 2680 5390 2880 5400
rect 3080 5390 3160 5400
rect 5080 5390 5120 5400
rect 5400 5390 5440 5400
rect 6160 5390 6200 5400
rect 6600 5390 6680 5400
rect 7320 5390 7400 5400
rect 7640 5390 7680 5400
rect 7760 5390 7800 5400
rect 7880 5390 7960 5400
rect 8320 5390 8360 5400
rect 8480 5390 8520 5400
rect 8840 5390 8880 5400
rect 9400 5390 9440 5400
rect 1960 5380 2040 5390
rect 2160 5380 2240 5390
rect 2360 5380 2400 5390
rect 2680 5380 2880 5390
rect 3080 5380 3160 5390
rect 5080 5380 5120 5390
rect 5400 5380 5440 5390
rect 6160 5380 6200 5390
rect 6600 5380 6680 5390
rect 7320 5380 7400 5390
rect 7640 5380 7680 5390
rect 7760 5380 7800 5390
rect 7880 5380 7960 5390
rect 8320 5380 8360 5390
rect 8480 5380 8520 5390
rect 8840 5380 8880 5390
rect 9400 5380 9440 5390
rect 400 5370 440 5380
rect 2000 5370 2040 5380
rect 2160 5370 2240 5380
rect 2360 5370 2400 5380
rect 2600 5370 2720 5380
rect 5080 5370 5120 5380
rect 5200 5370 5240 5380
rect 5400 5370 5600 5380
rect 5880 5370 5920 5380
rect 6160 5370 6200 5380
rect 6680 5370 6720 5380
rect 7320 5370 7400 5380
rect 7560 5370 7640 5380
rect 7880 5370 7960 5380
rect 8120 5370 8160 5380
rect 8200 5370 8240 5380
rect 8280 5370 8360 5380
rect 8400 5370 8440 5380
rect 8480 5370 8520 5380
rect 8760 5370 8800 5380
rect 8880 5370 8960 5380
rect 9440 5370 9520 5380
rect 9560 5370 9600 5380
rect 400 5360 440 5370
rect 2000 5360 2040 5370
rect 2160 5360 2240 5370
rect 2360 5360 2400 5370
rect 2600 5360 2720 5370
rect 5080 5360 5120 5370
rect 5200 5360 5240 5370
rect 5400 5360 5600 5370
rect 5880 5360 5920 5370
rect 6160 5360 6200 5370
rect 6680 5360 6720 5370
rect 7320 5360 7400 5370
rect 7560 5360 7640 5370
rect 7880 5360 7960 5370
rect 8120 5360 8160 5370
rect 8200 5360 8240 5370
rect 8280 5360 8360 5370
rect 8400 5360 8440 5370
rect 8480 5360 8520 5370
rect 8760 5360 8800 5370
rect 8880 5360 8960 5370
rect 9440 5360 9520 5370
rect 9560 5360 9600 5370
rect 400 5350 440 5360
rect 2000 5350 2040 5360
rect 2160 5350 2240 5360
rect 2360 5350 2400 5360
rect 2600 5350 2720 5360
rect 5080 5350 5120 5360
rect 5200 5350 5240 5360
rect 5400 5350 5600 5360
rect 5880 5350 5920 5360
rect 6160 5350 6200 5360
rect 6680 5350 6720 5360
rect 7320 5350 7400 5360
rect 7560 5350 7640 5360
rect 7880 5350 7960 5360
rect 8120 5350 8160 5360
rect 8200 5350 8240 5360
rect 8280 5350 8360 5360
rect 8400 5350 8440 5360
rect 8480 5350 8520 5360
rect 8760 5350 8800 5360
rect 8880 5350 8960 5360
rect 9440 5350 9520 5360
rect 9560 5350 9600 5360
rect 400 5340 440 5350
rect 2000 5340 2040 5350
rect 2160 5340 2240 5350
rect 2360 5340 2400 5350
rect 2600 5340 2720 5350
rect 5080 5340 5120 5350
rect 5200 5340 5240 5350
rect 5400 5340 5600 5350
rect 5880 5340 5920 5350
rect 6160 5340 6200 5350
rect 6680 5340 6720 5350
rect 7320 5340 7400 5350
rect 7560 5340 7640 5350
rect 7880 5340 7960 5350
rect 8120 5340 8160 5350
rect 8200 5340 8240 5350
rect 8280 5340 8360 5350
rect 8400 5340 8440 5350
rect 8480 5340 8520 5350
rect 8760 5340 8800 5350
rect 8880 5340 8960 5350
rect 9440 5340 9520 5350
rect 9560 5340 9600 5350
rect 240 5330 320 5340
rect 2000 5330 2120 5340
rect 2160 5330 2240 5340
rect 2360 5330 2400 5340
rect 2480 5330 2520 5340
rect 2600 5330 2720 5340
rect 3520 5330 3560 5340
rect 5120 5330 5160 5340
rect 5680 5330 5760 5340
rect 5800 5330 5880 5340
rect 6160 5330 6200 5340
rect 6560 5330 6640 5340
rect 6720 5330 6760 5340
rect 7280 5330 7360 5340
rect 7880 5330 8040 5340
rect 8160 5330 8240 5340
rect 8600 5330 8640 5340
rect 9120 5330 9160 5340
rect 9320 5330 9360 5340
rect 240 5320 320 5330
rect 2000 5320 2120 5330
rect 2160 5320 2240 5330
rect 2360 5320 2400 5330
rect 2480 5320 2520 5330
rect 2600 5320 2720 5330
rect 3520 5320 3560 5330
rect 5120 5320 5160 5330
rect 5680 5320 5760 5330
rect 5800 5320 5880 5330
rect 6160 5320 6200 5330
rect 6560 5320 6640 5330
rect 6720 5320 6760 5330
rect 7280 5320 7360 5330
rect 7880 5320 8040 5330
rect 8160 5320 8240 5330
rect 8600 5320 8640 5330
rect 9120 5320 9160 5330
rect 9320 5320 9360 5330
rect 240 5310 320 5320
rect 2000 5310 2120 5320
rect 2160 5310 2240 5320
rect 2360 5310 2400 5320
rect 2480 5310 2520 5320
rect 2600 5310 2720 5320
rect 3520 5310 3560 5320
rect 5120 5310 5160 5320
rect 5680 5310 5760 5320
rect 5800 5310 5880 5320
rect 6160 5310 6200 5320
rect 6560 5310 6640 5320
rect 6720 5310 6760 5320
rect 7280 5310 7360 5320
rect 7880 5310 8040 5320
rect 8160 5310 8240 5320
rect 8600 5310 8640 5320
rect 9120 5310 9160 5320
rect 9320 5310 9360 5320
rect 240 5300 320 5310
rect 2000 5300 2120 5310
rect 2160 5300 2240 5310
rect 2360 5300 2400 5310
rect 2480 5300 2520 5310
rect 2600 5300 2720 5310
rect 3520 5300 3560 5310
rect 5120 5300 5160 5310
rect 5680 5300 5760 5310
rect 5800 5300 5880 5310
rect 6160 5300 6200 5310
rect 6560 5300 6640 5310
rect 6720 5300 6760 5310
rect 7280 5300 7360 5310
rect 7880 5300 8040 5310
rect 8160 5300 8240 5310
rect 8600 5300 8640 5310
rect 9120 5300 9160 5310
rect 9320 5300 9360 5310
rect 2000 5290 2160 5300
rect 2200 5290 2240 5300
rect 2360 5290 2400 5300
rect 2440 5290 2480 5300
rect 2560 5290 2600 5300
rect 2640 5290 2800 5300
rect 5080 5290 5200 5300
rect 5680 5290 5840 5300
rect 6200 5290 6320 5300
rect 6360 5290 6440 5300
rect 7280 5290 7320 5300
rect 7920 5290 8000 5300
rect 8320 5290 8360 5300
rect 8520 5290 8560 5300
rect 9160 5290 9200 5300
rect 9240 5290 9280 5300
rect 9560 5290 9640 5300
rect 9840 5290 9880 5300
rect 9920 5290 9960 5300
rect 2000 5280 2160 5290
rect 2200 5280 2240 5290
rect 2360 5280 2400 5290
rect 2440 5280 2480 5290
rect 2560 5280 2600 5290
rect 2640 5280 2800 5290
rect 5080 5280 5200 5290
rect 5680 5280 5840 5290
rect 6200 5280 6320 5290
rect 6360 5280 6440 5290
rect 7280 5280 7320 5290
rect 7920 5280 8000 5290
rect 8320 5280 8360 5290
rect 8520 5280 8560 5290
rect 9160 5280 9200 5290
rect 9240 5280 9280 5290
rect 9560 5280 9640 5290
rect 9840 5280 9880 5290
rect 9920 5280 9960 5290
rect 2000 5270 2160 5280
rect 2200 5270 2240 5280
rect 2360 5270 2400 5280
rect 2440 5270 2480 5280
rect 2560 5270 2600 5280
rect 2640 5270 2800 5280
rect 5080 5270 5200 5280
rect 5680 5270 5840 5280
rect 6200 5270 6320 5280
rect 6360 5270 6440 5280
rect 7280 5270 7320 5280
rect 7920 5270 8000 5280
rect 8320 5270 8360 5280
rect 8520 5270 8560 5280
rect 9160 5270 9200 5280
rect 9240 5270 9280 5280
rect 9560 5270 9640 5280
rect 9840 5270 9880 5280
rect 9920 5270 9960 5280
rect 2000 5260 2160 5270
rect 2200 5260 2240 5270
rect 2360 5260 2400 5270
rect 2440 5260 2480 5270
rect 2560 5260 2600 5270
rect 2640 5260 2800 5270
rect 5080 5260 5200 5270
rect 5680 5260 5840 5270
rect 6200 5260 6320 5270
rect 6360 5260 6440 5270
rect 7280 5260 7320 5270
rect 7920 5260 8000 5270
rect 8320 5260 8360 5270
rect 8520 5260 8560 5270
rect 9160 5260 9200 5270
rect 9240 5260 9280 5270
rect 9560 5260 9640 5270
rect 9840 5260 9880 5270
rect 9920 5260 9960 5270
rect 600 5250 640 5260
rect 2040 5250 2160 5260
rect 2200 5250 2240 5260
rect 2400 5250 2480 5260
rect 2600 5250 2640 5260
rect 2680 5250 2720 5260
rect 2800 5250 2880 5260
rect 3480 5250 3520 5260
rect 5080 5250 5200 5260
rect 5680 5250 5720 5260
rect 6320 5250 6560 5260
rect 7280 5250 7360 5260
rect 7920 5250 8000 5260
rect 8360 5250 8400 5260
rect 8480 5250 8520 5260
rect 8840 5250 8880 5260
rect 9440 5250 9480 5260
rect 9800 5250 9840 5260
rect 9920 5250 9960 5260
rect 600 5240 640 5250
rect 2040 5240 2160 5250
rect 2200 5240 2240 5250
rect 2400 5240 2480 5250
rect 2600 5240 2640 5250
rect 2680 5240 2720 5250
rect 2800 5240 2880 5250
rect 3480 5240 3520 5250
rect 5080 5240 5200 5250
rect 5680 5240 5720 5250
rect 6320 5240 6560 5250
rect 7280 5240 7360 5250
rect 7920 5240 8000 5250
rect 8360 5240 8400 5250
rect 8480 5240 8520 5250
rect 8840 5240 8880 5250
rect 9440 5240 9480 5250
rect 9800 5240 9840 5250
rect 9920 5240 9960 5250
rect 600 5230 640 5240
rect 2040 5230 2160 5240
rect 2200 5230 2240 5240
rect 2400 5230 2480 5240
rect 2600 5230 2640 5240
rect 2680 5230 2720 5240
rect 2800 5230 2880 5240
rect 3480 5230 3520 5240
rect 5080 5230 5200 5240
rect 5680 5230 5720 5240
rect 6320 5230 6560 5240
rect 7280 5230 7360 5240
rect 7920 5230 8000 5240
rect 8360 5230 8400 5240
rect 8480 5230 8520 5240
rect 8840 5230 8880 5240
rect 9440 5230 9480 5240
rect 9800 5230 9840 5240
rect 9920 5230 9960 5240
rect 600 5220 640 5230
rect 2040 5220 2160 5230
rect 2200 5220 2240 5230
rect 2400 5220 2480 5230
rect 2600 5220 2640 5230
rect 2680 5220 2720 5230
rect 2800 5220 2880 5230
rect 3480 5220 3520 5230
rect 5080 5220 5200 5230
rect 5680 5220 5720 5230
rect 6320 5220 6560 5230
rect 7280 5220 7360 5230
rect 7920 5220 8000 5230
rect 8360 5220 8400 5230
rect 8480 5220 8520 5230
rect 8840 5220 8880 5230
rect 9440 5220 9480 5230
rect 9800 5220 9840 5230
rect 9920 5220 9960 5230
rect 600 5210 680 5220
rect 2040 5210 2240 5220
rect 2400 5210 2440 5220
rect 2720 5210 2760 5220
rect 2880 5210 2920 5220
rect 5160 5210 5200 5220
rect 7280 5210 7360 5220
rect 7960 5210 8000 5220
rect 8680 5210 8760 5220
rect 9000 5210 9040 5220
rect 9280 5210 9360 5220
rect 9520 5210 9600 5220
rect 9680 5210 9720 5220
rect 9840 5210 9880 5220
rect 600 5200 680 5210
rect 2040 5200 2240 5210
rect 2400 5200 2440 5210
rect 2720 5200 2760 5210
rect 2880 5200 2920 5210
rect 5160 5200 5200 5210
rect 7280 5200 7360 5210
rect 7960 5200 8000 5210
rect 8680 5200 8760 5210
rect 9000 5200 9040 5210
rect 9280 5200 9360 5210
rect 9520 5200 9600 5210
rect 9680 5200 9720 5210
rect 9840 5200 9880 5210
rect 600 5190 680 5200
rect 2040 5190 2240 5200
rect 2400 5190 2440 5200
rect 2720 5190 2760 5200
rect 2880 5190 2920 5200
rect 5160 5190 5200 5200
rect 7280 5190 7360 5200
rect 7960 5190 8000 5200
rect 8680 5190 8760 5200
rect 9000 5190 9040 5200
rect 9280 5190 9360 5200
rect 9520 5190 9600 5200
rect 9680 5190 9720 5200
rect 9840 5190 9880 5200
rect 600 5180 680 5190
rect 2040 5180 2240 5190
rect 2400 5180 2440 5190
rect 2720 5180 2760 5190
rect 2880 5180 2920 5190
rect 5160 5180 5200 5190
rect 7280 5180 7360 5190
rect 7960 5180 8000 5190
rect 8680 5180 8760 5190
rect 9000 5180 9040 5190
rect 9280 5180 9360 5190
rect 9520 5180 9600 5190
rect 9680 5180 9720 5190
rect 9840 5180 9880 5190
rect 600 5170 680 5180
rect 2040 5170 2200 5180
rect 2400 5170 2440 5180
rect 2840 5170 3000 5180
rect 3440 5170 3480 5180
rect 5080 5170 5120 5180
rect 5160 5170 5200 5180
rect 7320 5170 7360 5180
rect 7960 5170 8000 5180
rect 8120 5170 8160 5180
rect 9040 5170 9080 5180
rect 9160 5170 9200 5180
rect 9480 5170 9520 5180
rect 600 5160 680 5170
rect 2040 5160 2200 5170
rect 2400 5160 2440 5170
rect 2840 5160 3000 5170
rect 3440 5160 3480 5170
rect 5080 5160 5120 5170
rect 5160 5160 5200 5170
rect 7320 5160 7360 5170
rect 7960 5160 8000 5170
rect 8120 5160 8160 5170
rect 9040 5160 9080 5170
rect 9160 5160 9200 5170
rect 9480 5160 9520 5170
rect 600 5150 680 5160
rect 2040 5150 2200 5160
rect 2400 5150 2440 5160
rect 2840 5150 3000 5160
rect 3440 5150 3480 5160
rect 5080 5150 5120 5160
rect 5160 5150 5200 5160
rect 7320 5150 7360 5160
rect 7960 5150 8000 5160
rect 8120 5150 8160 5160
rect 9040 5150 9080 5160
rect 9160 5150 9200 5160
rect 9480 5150 9520 5160
rect 600 5140 680 5150
rect 2040 5140 2200 5150
rect 2400 5140 2440 5150
rect 2840 5140 3000 5150
rect 3440 5140 3480 5150
rect 5080 5140 5120 5150
rect 5160 5140 5200 5150
rect 7320 5140 7360 5150
rect 7960 5140 8000 5150
rect 8120 5140 8160 5150
rect 9040 5140 9080 5150
rect 9160 5140 9200 5150
rect 9480 5140 9520 5150
rect 520 5130 600 5140
rect 2080 5130 2200 5140
rect 2760 5130 2800 5140
rect 2920 5130 2960 5140
rect 5120 5130 5200 5140
rect 7960 5130 8000 5140
rect 8040 5130 8080 5140
rect 8400 5130 8440 5140
rect 8640 5130 8680 5140
rect 8880 5130 8920 5140
rect 8960 5130 9040 5140
rect 9240 5130 9280 5140
rect 9320 5130 9360 5140
rect 9840 5130 9920 5140
rect 520 5120 600 5130
rect 2080 5120 2200 5130
rect 2760 5120 2800 5130
rect 2920 5120 2960 5130
rect 5120 5120 5200 5130
rect 7960 5120 8000 5130
rect 8040 5120 8080 5130
rect 8400 5120 8440 5130
rect 8640 5120 8680 5130
rect 8880 5120 8920 5130
rect 8960 5120 9040 5130
rect 9240 5120 9280 5130
rect 9320 5120 9360 5130
rect 9840 5120 9920 5130
rect 520 5110 600 5120
rect 2080 5110 2200 5120
rect 2760 5110 2800 5120
rect 2920 5110 2960 5120
rect 5120 5110 5200 5120
rect 7960 5110 8000 5120
rect 8040 5110 8080 5120
rect 8400 5110 8440 5120
rect 8640 5110 8680 5120
rect 8880 5110 8920 5120
rect 8960 5110 9040 5120
rect 9240 5110 9280 5120
rect 9320 5110 9360 5120
rect 9840 5110 9920 5120
rect 520 5100 600 5110
rect 2080 5100 2200 5110
rect 2760 5100 2800 5110
rect 2920 5100 2960 5110
rect 5120 5100 5200 5110
rect 7960 5100 8000 5110
rect 8040 5100 8080 5110
rect 8400 5100 8440 5110
rect 8640 5100 8680 5110
rect 8880 5100 8920 5110
rect 8960 5100 9040 5110
rect 9240 5100 9280 5110
rect 9320 5100 9360 5110
rect 9840 5100 9920 5110
rect 440 5090 600 5100
rect 2080 5090 2280 5100
rect 2440 5090 2480 5100
rect 2800 5090 2840 5100
rect 8000 5090 8040 5100
rect 8400 5090 8440 5100
rect 8800 5090 8840 5100
rect 9080 5090 9120 5100
rect 9760 5090 9840 5100
rect 440 5080 600 5090
rect 2080 5080 2280 5090
rect 2440 5080 2480 5090
rect 2800 5080 2840 5090
rect 8000 5080 8040 5090
rect 8400 5080 8440 5090
rect 8800 5080 8840 5090
rect 9080 5080 9120 5090
rect 9760 5080 9840 5090
rect 440 5070 600 5080
rect 2080 5070 2280 5080
rect 2440 5070 2480 5080
rect 2800 5070 2840 5080
rect 8000 5070 8040 5080
rect 8400 5070 8440 5080
rect 8800 5070 8840 5080
rect 9080 5070 9120 5080
rect 9760 5070 9840 5080
rect 440 5060 600 5070
rect 2080 5060 2280 5070
rect 2440 5060 2480 5070
rect 2800 5060 2840 5070
rect 8000 5060 8040 5070
rect 8400 5060 8440 5070
rect 8800 5060 8840 5070
rect 9080 5060 9120 5070
rect 9760 5060 9840 5070
rect 360 5050 400 5060
rect 2080 5050 2280 5060
rect 2440 5050 2520 5060
rect 2640 5050 2880 5060
rect 5160 5050 5200 5060
rect 8000 5050 8040 5060
rect 8320 5050 8360 5060
rect 8480 5050 8520 5060
rect 8960 5050 9000 5060
rect 9080 5050 9120 5060
rect 9440 5050 9520 5060
rect 9600 5050 9640 5060
rect 360 5040 400 5050
rect 2080 5040 2280 5050
rect 2440 5040 2520 5050
rect 2640 5040 2880 5050
rect 5160 5040 5200 5050
rect 8000 5040 8040 5050
rect 8320 5040 8360 5050
rect 8480 5040 8520 5050
rect 8960 5040 9000 5050
rect 9080 5040 9120 5050
rect 9440 5040 9520 5050
rect 9600 5040 9640 5050
rect 360 5030 400 5040
rect 2080 5030 2280 5040
rect 2440 5030 2520 5040
rect 2640 5030 2880 5040
rect 5160 5030 5200 5040
rect 8000 5030 8040 5040
rect 8320 5030 8360 5040
rect 8480 5030 8520 5040
rect 8960 5030 9000 5040
rect 9080 5030 9120 5040
rect 9440 5030 9520 5040
rect 9600 5030 9640 5040
rect 360 5020 400 5030
rect 2080 5020 2280 5030
rect 2440 5020 2520 5030
rect 2640 5020 2880 5030
rect 5160 5020 5200 5030
rect 8000 5020 8040 5030
rect 8320 5020 8360 5030
rect 8480 5020 8520 5030
rect 8960 5020 9000 5030
rect 9080 5020 9120 5030
rect 9440 5020 9520 5030
rect 9600 5020 9640 5030
rect 360 5010 400 5020
rect 2120 5010 2320 5020
rect 2440 5010 2760 5020
rect 3360 5010 3400 5020
rect 5720 5010 5760 5020
rect 8040 5010 8080 5020
rect 8200 5010 8240 5020
rect 8760 5010 8840 5020
rect 8920 5010 8960 5020
rect 9000 5010 9040 5020
rect 9120 5010 9160 5020
rect 9320 5010 9360 5020
rect 9480 5010 9520 5020
rect 360 5000 400 5010
rect 2120 5000 2320 5010
rect 2440 5000 2760 5010
rect 3360 5000 3400 5010
rect 5720 5000 5760 5010
rect 8040 5000 8080 5010
rect 8200 5000 8240 5010
rect 8760 5000 8840 5010
rect 8920 5000 8960 5010
rect 9000 5000 9040 5010
rect 9120 5000 9160 5010
rect 9320 5000 9360 5010
rect 9480 5000 9520 5010
rect 360 4990 400 5000
rect 2120 4990 2320 5000
rect 2440 4990 2760 5000
rect 3360 4990 3400 5000
rect 5720 4990 5760 5000
rect 8040 4990 8080 5000
rect 8200 4990 8240 5000
rect 8760 4990 8840 5000
rect 8920 4990 8960 5000
rect 9000 4990 9040 5000
rect 9120 4990 9160 5000
rect 9320 4990 9360 5000
rect 9480 4990 9520 5000
rect 360 4980 400 4990
rect 2120 4980 2320 4990
rect 2440 4980 2760 4990
rect 3360 4980 3400 4990
rect 5720 4980 5760 4990
rect 8040 4980 8080 4990
rect 8200 4980 8240 4990
rect 8760 4980 8840 4990
rect 8920 4980 8960 4990
rect 9000 4980 9040 4990
rect 9120 4980 9160 4990
rect 9320 4980 9360 4990
rect 9480 4980 9520 4990
rect 240 4970 280 4980
rect 360 4970 400 4980
rect 2160 4970 2320 4980
rect 2480 4970 2680 4980
rect 2720 4970 2760 4980
rect 4040 4970 4080 4980
rect 4280 4970 4320 4980
rect 5640 4970 5760 4980
rect 6320 4970 6400 4980
rect 7920 4970 7960 4980
rect 8200 4970 8240 4980
rect 8280 4970 8320 4980
rect 8400 4970 8440 4980
rect 8840 4970 8880 4980
rect 9080 4970 9120 4980
rect 9200 4970 9240 4980
rect 9600 4970 9640 4980
rect 240 4960 280 4970
rect 360 4960 400 4970
rect 2160 4960 2320 4970
rect 2480 4960 2680 4970
rect 2720 4960 2760 4970
rect 4040 4960 4080 4970
rect 4280 4960 4320 4970
rect 5640 4960 5760 4970
rect 6320 4960 6400 4970
rect 7920 4960 7960 4970
rect 8200 4960 8240 4970
rect 8280 4960 8320 4970
rect 8400 4960 8440 4970
rect 8840 4960 8880 4970
rect 9080 4960 9120 4970
rect 9200 4960 9240 4970
rect 9600 4960 9640 4970
rect 240 4950 280 4960
rect 360 4950 400 4960
rect 2160 4950 2320 4960
rect 2480 4950 2680 4960
rect 2720 4950 2760 4960
rect 4040 4950 4080 4960
rect 4280 4950 4320 4960
rect 5640 4950 5760 4960
rect 6320 4950 6400 4960
rect 7920 4950 7960 4960
rect 8200 4950 8240 4960
rect 8280 4950 8320 4960
rect 8400 4950 8440 4960
rect 8840 4950 8880 4960
rect 9080 4950 9120 4960
rect 9200 4950 9240 4960
rect 9600 4950 9640 4960
rect 240 4940 280 4950
rect 360 4940 400 4950
rect 2160 4940 2320 4950
rect 2480 4940 2680 4950
rect 2720 4940 2760 4950
rect 4040 4940 4080 4950
rect 4280 4940 4320 4950
rect 5640 4940 5760 4950
rect 6320 4940 6400 4950
rect 7920 4940 7960 4950
rect 8200 4940 8240 4950
rect 8280 4940 8320 4950
rect 8400 4940 8440 4950
rect 8840 4940 8880 4950
rect 9080 4940 9120 4950
rect 9200 4940 9240 4950
rect 9600 4940 9640 4950
rect 80 4930 240 4940
rect 320 4930 400 4940
rect 2200 4930 2240 4940
rect 2320 4930 2360 4940
rect 2480 4930 2640 4940
rect 3320 4930 3360 4940
rect 4440 4930 4480 4940
rect 5560 4930 5640 4940
rect 5800 4930 5840 4940
rect 5920 4930 5960 4940
rect 6120 4930 6320 4940
rect 6400 4930 6440 4940
rect 7320 4930 7360 4940
rect 7680 4930 7720 4940
rect 7800 4930 7840 4940
rect 8480 4930 8520 4940
rect 8680 4930 8760 4940
rect 8840 4930 8880 4940
rect 9040 4930 9120 4940
rect 9280 4930 9320 4940
rect 9440 4930 9480 4940
rect 9680 4930 9720 4940
rect 80 4920 240 4930
rect 320 4920 400 4930
rect 2200 4920 2240 4930
rect 2320 4920 2360 4930
rect 2480 4920 2640 4930
rect 3320 4920 3360 4930
rect 4440 4920 4480 4930
rect 5560 4920 5640 4930
rect 5800 4920 5840 4930
rect 5920 4920 5960 4930
rect 6120 4920 6320 4930
rect 6400 4920 6440 4930
rect 7320 4920 7360 4930
rect 7680 4920 7720 4930
rect 7800 4920 7840 4930
rect 8480 4920 8520 4930
rect 8680 4920 8760 4930
rect 8840 4920 8880 4930
rect 9040 4920 9120 4930
rect 9280 4920 9320 4930
rect 9440 4920 9480 4930
rect 9680 4920 9720 4930
rect 80 4910 240 4920
rect 320 4910 400 4920
rect 2200 4910 2240 4920
rect 2320 4910 2360 4920
rect 2480 4910 2640 4920
rect 3320 4910 3360 4920
rect 4440 4910 4480 4920
rect 5560 4910 5640 4920
rect 5800 4910 5840 4920
rect 5920 4910 5960 4920
rect 6120 4910 6320 4920
rect 6400 4910 6440 4920
rect 7320 4910 7360 4920
rect 7680 4910 7720 4920
rect 7800 4910 7840 4920
rect 8480 4910 8520 4920
rect 8680 4910 8760 4920
rect 8840 4910 8880 4920
rect 9040 4910 9120 4920
rect 9280 4910 9320 4920
rect 9440 4910 9480 4920
rect 9680 4910 9720 4920
rect 80 4900 240 4910
rect 320 4900 400 4910
rect 2200 4900 2240 4910
rect 2320 4900 2360 4910
rect 2480 4900 2640 4910
rect 3320 4900 3360 4910
rect 4440 4900 4480 4910
rect 5560 4900 5640 4910
rect 5800 4900 5840 4910
rect 5920 4900 5960 4910
rect 6120 4900 6320 4910
rect 6400 4900 6440 4910
rect 7320 4900 7360 4910
rect 7680 4900 7720 4910
rect 7800 4900 7840 4910
rect 8480 4900 8520 4910
rect 8680 4900 8760 4910
rect 8840 4900 8880 4910
rect 9040 4900 9120 4910
rect 9280 4900 9320 4910
rect 9440 4900 9480 4910
rect 9680 4900 9720 4910
rect 0 4890 80 4900
rect 2560 4890 2680 4900
rect 3880 4890 4080 4900
rect 4760 4890 4840 4900
rect 5520 4890 5600 4900
rect 5680 4890 5720 4900
rect 5800 4890 5840 4900
rect 5960 4890 6040 4900
rect 6080 4890 6120 4900
rect 6440 4890 6480 4900
rect 7320 4890 7360 4900
rect 7880 4890 7920 4900
rect 8080 4890 8160 4900
rect 8440 4890 8480 4900
rect 8840 4890 8880 4900
rect 9000 4890 9040 4900
rect 9360 4890 9400 4900
rect 9600 4890 9640 4900
rect 9680 4890 9720 4900
rect 0 4880 80 4890
rect 2560 4880 2680 4890
rect 3880 4880 4080 4890
rect 4760 4880 4840 4890
rect 5520 4880 5600 4890
rect 5680 4880 5720 4890
rect 5800 4880 5840 4890
rect 5960 4880 6040 4890
rect 6080 4880 6120 4890
rect 6440 4880 6480 4890
rect 7320 4880 7360 4890
rect 7880 4880 7920 4890
rect 8080 4880 8160 4890
rect 8440 4880 8480 4890
rect 8840 4880 8880 4890
rect 9000 4880 9040 4890
rect 9360 4880 9400 4890
rect 9600 4880 9640 4890
rect 9680 4880 9720 4890
rect 0 4870 80 4880
rect 2560 4870 2680 4880
rect 3880 4870 4080 4880
rect 4760 4870 4840 4880
rect 5520 4870 5600 4880
rect 5680 4870 5720 4880
rect 5800 4870 5840 4880
rect 5960 4870 6040 4880
rect 6080 4870 6120 4880
rect 6440 4870 6480 4880
rect 7320 4870 7360 4880
rect 7880 4870 7920 4880
rect 8080 4870 8160 4880
rect 8440 4870 8480 4880
rect 8840 4870 8880 4880
rect 9000 4870 9040 4880
rect 9360 4870 9400 4880
rect 9600 4870 9640 4880
rect 9680 4870 9720 4880
rect 0 4860 80 4870
rect 2560 4860 2680 4870
rect 3880 4860 4080 4870
rect 4760 4860 4840 4870
rect 5520 4860 5600 4870
rect 5680 4860 5720 4870
rect 5800 4860 5840 4870
rect 5960 4860 6040 4870
rect 6080 4860 6120 4870
rect 6440 4860 6480 4870
rect 7320 4860 7360 4870
rect 7880 4860 7920 4870
rect 8080 4860 8160 4870
rect 8440 4860 8480 4870
rect 8840 4860 8880 4870
rect 9000 4860 9040 4870
rect 9360 4860 9400 4870
rect 9600 4860 9640 4870
rect 9680 4860 9720 4870
rect 0 4850 160 4860
rect 2360 4850 2400 4860
rect 2640 4850 2680 4860
rect 3720 4850 3840 4860
rect 3960 4850 4000 4860
rect 4920 4850 4960 4860
rect 5480 4850 5560 4860
rect 5680 4850 5720 4860
rect 5840 4850 6000 4860
rect 6480 4850 6520 4860
rect 8200 4850 8280 4860
rect 8360 4850 8400 4860
rect 8560 4850 8640 4860
rect 8720 4850 8760 4860
rect 8840 4850 8880 4860
rect 9040 4850 9080 4860
rect 9320 4850 9360 4860
rect 9440 4850 9480 4860
rect 0 4840 160 4850
rect 2360 4840 2400 4850
rect 2640 4840 2680 4850
rect 3720 4840 3840 4850
rect 3960 4840 4000 4850
rect 4920 4840 4960 4850
rect 5480 4840 5560 4850
rect 5680 4840 5720 4850
rect 5840 4840 6000 4850
rect 6480 4840 6520 4850
rect 8200 4840 8280 4850
rect 8360 4840 8400 4850
rect 8560 4840 8640 4850
rect 8720 4840 8760 4850
rect 8840 4840 8880 4850
rect 9040 4840 9080 4850
rect 9320 4840 9360 4850
rect 9440 4840 9480 4850
rect 0 4830 160 4840
rect 2360 4830 2400 4840
rect 2640 4830 2680 4840
rect 3720 4830 3840 4840
rect 3960 4830 4000 4840
rect 4920 4830 4960 4840
rect 5480 4830 5560 4840
rect 5680 4830 5720 4840
rect 5840 4830 6000 4840
rect 6480 4830 6520 4840
rect 8200 4830 8280 4840
rect 8360 4830 8400 4840
rect 8560 4830 8640 4840
rect 8720 4830 8760 4840
rect 8840 4830 8880 4840
rect 9040 4830 9080 4840
rect 9320 4830 9360 4840
rect 9440 4830 9480 4840
rect 0 4820 160 4830
rect 2360 4820 2400 4830
rect 2640 4820 2680 4830
rect 3720 4820 3840 4830
rect 3960 4820 4000 4830
rect 4920 4820 4960 4830
rect 5480 4820 5560 4830
rect 5680 4820 5720 4830
rect 5840 4820 6000 4830
rect 6480 4820 6520 4830
rect 8200 4820 8280 4830
rect 8360 4820 8400 4830
rect 8560 4820 8640 4830
rect 8720 4820 8760 4830
rect 8840 4820 8880 4830
rect 9040 4820 9080 4830
rect 9320 4820 9360 4830
rect 9440 4820 9480 4830
rect 0 4810 200 4820
rect 2360 4810 2400 4820
rect 2680 4810 2760 4820
rect 5000 4810 5040 4820
rect 5440 4810 5520 4820
rect 5640 4810 5680 4820
rect 5960 4810 6000 4820
rect 6240 4810 6360 4820
rect 6520 4810 6560 4820
rect 7680 4810 7720 4820
rect 7760 4810 7840 4820
rect 8000 4810 8080 4820
rect 8160 4810 8200 4820
rect 8240 4810 8280 4820
rect 8360 4810 8400 4820
rect 8520 4810 8560 4820
rect 8600 4810 8640 4820
rect 9600 4810 9680 4820
rect 0 4800 200 4810
rect 2360 4800 2400 4810
rect 2680 4800 2760 4810
rect 5000 4800 5040 4810
rect 5440 4800 5520 4810
rect 5640 4800 5680 4810
rect 5960 4800 6000 4810
rect 6240 4800 6360 4810
rect 6520 4800 6560 4810
rect 7680 4800 7720 4810
rect 7760 4800 7840 4810
rect 8000 4800 8080 4810
rect 8160 4800 8200 4810
rect 8240 4800 8280 4810
rect 8360 4800 8400 4810
rect 8520 4800 8560 4810
rect 8600 4800 8640 4810
rect 9600 4800 9680 4810
rect 0 4790 200 4800
rect 2360 4790 2400 4800
rect 2680 4790 2760 4800
rect 5000 4790 5040 4800
rect 5440 4790 5520 4800
rect 5640 4790 5680 4800
rect 5960 4790 6000 4800
rect 6240 4790 6360 4800
rect 6520 4790 6560 4800
rect 7680 4790 7720 4800
rect 7760 4790 7840 4800
rect 8000 4790 8080 4800
rect 8160 4790 8200 4800
rect 8240 4790 8280 4800
rect 8360 4790 8400 4800
rect 8520 4790 8560 4800
rect 8600 4790 8640 4800
rect 9600 4790 9680 4800
rect 0 4780 200 4790
rect 2360 4780 2400 4790
rect 2680 4780 2760 4790
rect 5000 4780 5040 4790
rect 5440 4780 5520 4790
rect 5640 4780 5680 4790
rect 5960 4780 6000 4790
rect 6240 4780 6360 4790
rect 6520 4780 6560 4790
rect 7680 4780 7720 4790
rect 7760 4780 7840 4790
rect 8000 4780 8080 4790
rect 8160 4780 8200 4790
rect 8240 4780 8280 4790
rect 8360 4780 8400 4790
rect 8520 4780 8560 4790
rect 8600 4780 8640 4790
rect 9600 4780 9680 4790
rect 0 4770 160 4780
rect 2440 4770 2480 4780
rect 2720 4770 2840 4780
rect 3320 4770 3360 4780
rect 5040 4770 5080 4780
rect 5400 4770 5480 4780
rect 5600 4770 5640 4780
rect 6000 4770 6400 4780
rect 6560 4770 6640 4780
rect 7880 4770 8000 4780
rect 8240 4770 8360 4780
rect 8480 4770 8560 4780
rect 8960 4770 9000 4780
rect 9400 4770 9520 4780
rect 9880 4770 9990 4780
rect 0 4760 160 4770
rect 2440 4760 2480 4770
rect 2720 4760 2840 4770
rect 3320 4760 3360 4770
rect 5040 4760 5080 4770
rect 5400 4760 5480 4770
rect 5600 4760 5640 4770
rect 6000 4760 6400 4770
rect 6560 4760 6640 4770
rect 7880 4760 8000 4770
rect 8240 4760 8360 4770
rect 8480 4760 8560 4770
rect 8960 4760 9000 4770
rect 9400 4760 9520 4770
rect 9880 4760 9990 4770
rect 0 4750 160 4760
rect 2440 4750 2480 4760
rect 2720 4750 2840 4760
rect 3320 4750 3360 4760
rect 5040 4750 5080 4760
rect 5400 4750 5480 4760
rect 5600 4750 5640 4760
rect 6000 4750 6400 4760
rect 6560 4750 6640 4760
rect 7880 4750 8000 4760
rect 8240 4750 8360 4760
rect 8480 4750 8560 4760
rect 8960 4750 9000 4760
rect 9400 4750 9520 4760
rect 9880 4750 9990 4760
rect 0 4740 160 4750
rect 2440 4740 2480 4750
rect 2720 4740 2840 4750
rect 3320 4740 3360 4750
rect 5040 4740 5080 4750
rect 5400 4740 5480 4750
rect 5600 4740 5640 4750
rect 6000 4740 6400 4750
rect 6560 4740 6640 4750
rect 7880 4740 8000 4750
rect 8240 4740 8360 4750
rect 8480 4740 8560 4750
rect 8960 4740 9000 4750
rect 9400 4740 9520 4750
rect 9880 4740 9990 4750
rect 0 4730 160 4740
rect 2520 4730 2560 4740
rect 2720 4730 2840 4740
rect 2960 4730 3000 4740
rect 3240 4730 3320 4740
rect 3520 4730 3560 4740
rect 5400 4730 5480 4740
rect 5600 4730 5640 4740
rect 6040 4730 6240 4740
rect 6320 4730 6440 4740
rect 6560 4730 6640 4740
rect 7720 4730 7760 4740
rect 7800 4730 7840 4740
rect 7960 4730 8000 4740
rect 8360 4730 8400 4740
rect 8600 4730 8680 4740
rect 8760 4730 8800 4740
rect 8880 4730 8920 4740
rect 9280 4730 9360 4740
rect 0 4720 160 4730
rect 2520 4720 2560 4730
rect 2720 4720 2840 4730
rect 2960 4720 3000 4730
rect 3240 4720 3320 4730
rect 3520 4720 3560 4730
rect 5400 4720 5480 4730
rect 5600 4720 5640 4730
rect 6040 4720 6240 4730
rect 6320 4720 6440 4730
rect 6560 4720 6640 4730
rect 7720 4720 7760 4730
rect 7800 4720 7840 4730
rect 7960 4720 8000 4730
rect 8360 4720 8400 4730
rect 8600 4720 8680 4730
rect 8760 4720 8800 4730
rect 8880 4720 8920 4730
rect 9280 4720 9360 4730
rect 0 4710 160 4720
rect 2520 4710 2560 4720
rect 2720 4710 2840 4720
rect 2960 4710 3000 4720
rect 3240 4710 3320 4720
rect 3520 4710 3560 4720
rect 5400 4710 5480 4720
rect 5600 4710 5640 4720
rect 6040 4710 6240 4720
rect 6320 4710 6440 4720
rect 6560 4710 6640 4720
rect 7720 4710 7760 4720
rect 7800 4710 7840 4720
rect 7960 4710 8000 4720
rect 8360 4710 8400 4720
rect 8600 4710 8680 4720
rect 8760 4710 8800 4720
rect 8880 4710 8920 4720
rect 9280 4710 9360 4720
rect 0 4700 160 4710
rect 2520 4700 2560 4710
rect 2720 4700 2840 4710
rect 2960 4700 3000 4710
rect 3240 4700 3320 4710
rect 3520 4700 3560 4710
rect 5400 4700 5480 4710
rect 5600 4700 5640 4710
rect 6040 4700 6240 4710
rect 6320 4700 6440 4710
rect 6560 4700 6640 4710
rect 7720 4700 7760 4710
rect 7800 4700 7840 4710
rect 7960 4700 8000 4710
rect 8360 4700 8400 4710
rect 8600 4700 8680 4710
rect 8760 4700 8800 4710
rect 8880 4700 8920 4710
rect 9280 4700 9360 4710
rect 0 4690 120 4700
rect 2560 4690 2600 4700
rect 2960 4690 3000 4700
rect 3120 4690 3160 4700
rect 3240 4690 3320 4700
rect 3480 4690 3520 4700
rect 5120 4690 5160 4700
rect 5400 4690 5480 4700
rect 5640 4690 5760 4700
rect 6320 4690 6440 4700
rect 6560 4690 6640 4700
rect 7680 4690 7720 4700
rect 7960 4690 8000 4700
rect 8120 4690 8160 4700
rect 8240 4690 8280 4700
rect 8480 4690 8560 4700
rect 8640 4690 8680 4700
rect 8760 4690 8800 4700
rect 8840 4690 8880 4700
rect 0 4680 120 4690
rect 2560 4680 2600 4690
rect 2960 4680 3000 4690
rect 3120 4680 3160 4690
rect 3240 4680 3320 4690
rect 3480 4680 3520 4690
rect 5120 4680 5160 4690
rect 5400 4680 5480 4690
rect 5640 4680 5760 4690
rect 6320 4680 6440 4690
rect 6560 4680 6640 4690
rect 7680 4680 7720 4690
rect 7960 4680 8000 4690
rect 8120 4680 8160 4690
rect 8240 4680 8280 4690
rect 8480 4680 8560 4690
rect 8640 4680 8680 4690
rect 8760 4680 8800 4690
rect 8840 4680 8880 4690
rect 0 4670 120 4680
rect 2560 4670 2600 4680
rect 2960 4670 3000 4680
rect 3120 4670 3160 4680
rect 3240 4670 3320 4680
rect 3480 4670 3520 4680
rect 5120 4670 5160 4680
rect 5400 4670 5480 4680
rect 5640 4670 5760 4680
rect 6320 4670 6440 4680
rect 6560 4670 6640 4680
rect 7680 4670 7720 4680
rect 7960 4670 8000 4680
rect 8120 4670 8160 4680
rect 8240 4670 8280 4680
rect 8480 4670 8560 4680
rect 8640 4670 8680 4680
rect 8760 4670 8800 4680
rect 8840 4670 8880 4680
rect 0 4660 120 4670
rect 2560 4660 2600 4670
rect 2960 4660 3000 4670
rect 3120 4660 3160 4670
rect 3240 4660 3320 4670
rect 3480 4660 3520 4670
rect 5120 4660 5160 4670
rect 5400 4660 5480 4670
rect 5640 4660 5760 4670
rect 6320 4660 6440 4670
rect 6560 4660 6640 4670
rect 7680 4660 7720 4670
rect 7960 4660 8000 4670
rect 8120 4660 8160 4670
rect 8240 4660 8280 4670
rect 8480 4660 8560 4670
rect 8640 4660 8680 4670
rect 8760 4660 8800 4670
rect 8840 4660 8880 4670
rect 5400 4650 5520 4660
rect 5800 4650 6080 4660
rect 6200 4650 6400 4660
rect 6560 4650 6640 4660
rect 7680 4650 7720 4660
rect 7880 4650 7920 4660
rect 8080 4650 8120 4660
rect 8280 4650 8320 4660
rect 8640 4650 8680 4660
rect 8920 4650 8960 4660
rect 5400 4640 5520 4650
rect 5800 4640 6080 4650
rect 6200 4640 6400 4650
rect 6560 4640 6640 4650
rect 7680 4640 7720 4650
rect 7880 4640 7920 4650
rect 8080 4640 8120 4650
rect 8280 4640 8320 4650
rect 8640 4640 8680 4650
rect 8920 4640 8960 4650
rect 5400 4630 5520 4640
rect 5800 4630 6080 4640
rect 6200 4630 6400 4640
rect 6560 4630 6640 4640
rect 7680 4630 7720 4640
rect 7880 4630 7920 4640
rect 8080 4630 8120 4640
rect 8280 4630 8320 4640
rect 8640 4630 8680 4640
rect 8920 4630 8960 4640
rect 5400 4620 5520 4630
rect 5800 4620 6080 4630
rect 6200 4620 6400 4630
rect 6560 4620 6640 4630
rect 7680 4620 7720 4630
rect 7880 4620 7920 4630
rect 8080 4620 8120 4630
rect 8280 4620 8320 4630
rect 8640 4620 8680 4630
rect 8920 4620 8960 4630
rect 3440 4610 3480 4620
rect 5200 4610 5240 4620
rect 5400 4610 5520 4620
rect 5600 4610 5640 4620
rect 5760 4610 5920 4620
rect 6000 4610 6120 4620
rect 6560 4610 6600 4620
rect 7680 4610 7720 4620
rect 8240 4610 8280 4620
rect 8800 4610 8880 4620
rect 3440 4600 3480 4610
rect 5200 4600 5240 4610
rect 5400 4600 5520 4610
rect 5600 4600 5640 4610
rect 5760 4600 5920 4610
rect 6000 4600 6120 4610
rect 6560 4600 6600 4610
rect 7680 4600 7720 4610
rect 8240 4600 8280 4610
rect 8800 4600 8880 4610
rect 3440 4590 3480 4600
rect 5200 4590 5240 4600
rect 5400 4590 5520 4600
rect 5600 4590 5640 4600
rect 5760 4590 5920 4600
rect 6000 4590 6120 4600
rect 6560 4590 6600 4600
rect 7680 4590 7720 4600
rect 8240 4590 8280 4600
rect 8800 4590 8880 4600
rect 3440 4580 3480 4590
rect 5200 4580 5240 4590
rect 5400 4580 5520 4590
rect 5600 4580 5640 4590
rect 5760 4580 5920 4590
rect 6000 4580 6120 4590
rect 6560 4580 6600 4590
rect 7680 4580 7720 4590
rect 8240 4580 8280 4590
rect 8800 4580 8880 4590
rect 5440 4570 5560 4580
rect 5640 4570 5680 4580
rect 6160 4570 6280 4580
rect 6520 4570 6560 4580
rect 7360 4570 7400 4580
rect 7760 4570 7800 4580
rect 8000 4570 8040 4580
rect 8120 4570 8160 4580
rect 8200 4570 8240 4580
rect 8640 4570 8680 4580
rect 5440 4560 5560 4570
rect 5640 4560 5680 4570
rect 6160 4560 6280 4570
rect 6520 4560 6560 4570
rect 7360 4560 7400 4570
rect 7760 4560 7800 4570
rect 8000 4560 8040 4570
rect 8120 4560 8160 4570
rect 8200 4560 8240 4570
rect 8640 4560 8680 4570
rect 5440 4550 5560 4560
rect 5640 4550 5680 4560
rect 6160 4550 6280 4560
rect 6520 4550 6560 4560
rect 7360 4550 7400 4560
rect 7760 4550 7800 4560
rect 8000 4550 8040 4560
rect 8120 4550 8160 4560
rect 8200 4550 8240 4560
rect 8640 4550 8680 4560
rect 5440 4540 5560 4550
rect 5640 4540 5680 4550
rect 6160 4540 6280 4550
rect 6520 4540 6560 4550
rect 7360 4540 7400 4550
rect 7760 4540 7800 4550
rect 8000 4540 8040 4550
rect 8120 4540 8160 4550
rect 8200 4540 8240 4550
rect 8640 4540 8680 4550
rect 3000 4530 3040 4540
rect 5240 4530 5280 4540
rect 5480 4530 5600 4540
rect 5680 4530 5720 4540
rect 5800 4530 5840 4540
rect 6240 4530 6280 4540
rect 7640 4530 7680 4540
rect 7800 4530 7840 4540
rect 8240 4530 8280 4540
rect 9960 4530 9990 4540
rect 3000 4520 3040 4530
rect 5240 4520 5280 4530
rect 5480 4520 5600 4530
rect 5680 4520 5720 4530
rect 5800 4520 5840 4530
rect 6240 4520 6280 4530
rect 7640 4520 7680 4530
rect 7800 4520 7840 4530
rect 8240 4520 8280 4530
rect 9960 4520 9990 4530
rect 3000 4510 3040 4520
rect 5240 4510 5280 4520
rect 5480 4510 5600 4520
rect 5680 4510 5720 4520
rect 5800 4510 5840 4520
rect 6240 4510 6280 4520
rect 7640 4510 7680 4520
rect 7800 4510 7840 4520
rect 8240 4510 8280 4520
rect 9960 4510 9990 4520
rect 3000 4500 3040 4510
rect 5240 4500 5280 4510
rect 5480 4500 5600 4510
rect 5680 4500 5720 4510
rect 5800 4500 5840 4510
rect 6240 4500 6280 4510
rect 7640 4500 7680 4510
rect 7800 4500 7840 4510
rect 8240 4500 8280 4510
rect 9960 4500 9990 4510
rect 3080 4490 3120 4500
rect 3240 4490 3280 4500
rect 5320 4490 5360 4500
rect 5480 4490 5600 4500
rect 5720 4490 5760 4500
rect 6200 4490 6240 4500
rect 7840 4490 7880 4500
rect 7920 4490 7960 4500
rect 8000 4490 8040 4500
rect 8280 4490 8400 4500
rect 9920 4490 9960 4500
rect 3080 4480 3120 4490
rect 3240 4480 3280 4490
rect 5320 4480 5360 4490
rect 5480 4480 5600 4490
rect 5720 4480 5760 4490
rect 6200 4480 6240 4490
rect 7840 4480 7880 4490
rect 7920 4480 7960 4490
rect 8000 4480 8040 4490
rect 8280 4480 8400 4490
rect 9920 4480 9960 4490
rect 3080 4470 3120 4480
rect 3240 4470 3280 4480
rect 5320 4470 5360 4480
rect 5480 4470 5600 4480
rect 5720 4470 5760 4480
rect 6200 4470 6240 4480
rect 7840 4470 7880 4480
rect 7920 4470 7960 4480
rect 8000 4470 8040 4480
rect 8280 4470 8400 4480
rect 9920 4470 9960 4480
rect 3080 4460 3120 4470
rect 3240 4460 3280 4470
rect 5320 4460 5360 4470
rect 5480 4460 5600 4470
rect 5720 4460 5760 4470
rect 6200 4460 6240 4470
rect 7840 4460 7880 4470
rect 7920 4460 7960 4470
rect 8000 4460 8040 4470
rect 8280 4460 8400 4470
rect 9920 4460 9960 4470
rect 3040 4450 3120 4460
rect 3240 4450 3280 4460
rect 5280 4450 5320 4460
rect 5520 4450 5600 4460
rect 5760 4450 5800 4460
rect 6120 4450 6200 4460
rect 6360 4450 6440 4460
rect 6480 4450 6520 4460
rect 7400 4450 7440 4460
rect 7920 4450 7960 4460
rect 8000 4450 8040 4460
rect 8160 4450 8200 4460
rect 8240 4450 8280 4460
rect 8840 4450 8880 4460
rect 9200 4450 9240 4460
rect 9880 4450 9920 4460
rect 3040 4440 3120 4450
rect 3240 4440 3280 4450
rect 5280 4440 5320 4450
rect 5520 4440 5600 4450
rect 5760 4440 5800 4450
rect 6120 4440 6200 4450
rect 6360 4440 6440 4450
rect 6480 4440 6520 4450
rect 7400 4440 7440 4450
rect 7920 4440 7960 4450
rect 8000 4440 8040 4450
rect 8160 4440 8200 4450
rect 8240 4440 8280 4450
rect 8840 4440 8880 4450
rect 9200 4440 9240 4450
rect 9880 4440 9920 4450
rect 3040 4430 3120 4440
rect 3240 4430 3280 4440
rect 5280 4430 5320 4440
rect 5520 4430 5600 4440
rect 5760 4430 5800 4440
rect 6120 4430 6200 4440
rect 6360 4430 6440 4440
rect 6480 4430 6520 4440
rect 7400 4430 7440 4440
rect 7920 4430 7960 4440
rect 8000 4430 8040 4440
rect 8160 4430 8200 4440
rect 8240 4430 8280 4440
rect 8840 4430 8880 4440
rect 9200 4430 9240 4440
rect 9880 4430 9920 4440
rect 3040 4420 3120 4430
rect 3240 4420 3280 4430
rect 5280 4420 5320 4430
rect 5520 4420 5600 4430
rect 5760 4420 5800 4430
rect 6120 4420 6200 4430
rect 6360 4420 6440 4430
rect 6480 4420 6520 4430
rect 7400 4420 7440 4430
rect 7920 4420 7960 4430
rect 8000 4420 8040 4430
rect 8160 4420 8200 4430
rect 8240 4420 8280 4430
rect 8840 4420 8880 4430
rect 9200 4420 9240 4430
rect 9880 4420 9920 4430
rect 3040 4410 3080 4420
rect 3280 4410 3320 4420
rect 4600 4410 4720 4420
rect 5400 4410 5440 4420
rect 5520 4410 5560 4420
rect 6000 4410 6200 4420
rect 6320 4410 6520 4420
rect 7840 4410 7920 4420
rect 8040 4410 8080 4420
rect 8680 4410 8720 4420
rect 9840 4410 9880 4420
rect 3040 4400 3080 4410
rect 3280 4400 3320 4410
rect 4600 4400 4720 4410
rect 5400 4400 5440 4410
rect 5520 4400 5560 4410
rect 6000 4400 6200 4410
rect 6320 4400 6520 4410
rect 7840 4400 7920 4410
rect 8040 4400 8080 4410
rect 8680 4400 8720 4410
rect 9840 4400 9880 4410
rect 3040 4390 3080 4400
rect 3280 4390 3320 4400
rect 4600 4390 4720 4400
rect 5400 4390 5440 4400
rect 5520 4390 5560 4400
rect 6000 4390 6200 4400
rect 6320 4390 6520 4400
rect 7840 4390 7920 4400
rect 8040 4390 8080 4400
rect 8680 4390 8720 4400
rect 9840 4390 9880 4400
rect 3040 4380 3080 4390
rect 3280 4380 3320 4390
rect 4600 4380 4720 4390
rect 5400 4380 5440 4390
rect 5520 4380 5560 4390
rect 6000 4380 6200 4390
rect 6320 4380 6520 4390
rect 7840 4380 7920 4390
rect 8040 4380 8080 4390
rect 8680 4380 8720 4390
rect 9840 4380 9880 4390
rect 2920 4370 2960 4380
rect 3040 4370 3080 4380
rect 3240 4370 3320 4380
rect 4560 4370 4600 4380
rect 4760 4370 4880 4380
rect 5400 4370 5480 4380
rect 5960 4370 6480 4380
rect 7400 4370 7440 4380
rect 7800 4370 7880 4380
rect 8520 4370 8680 4380
rect 9840 4370 9880 4380
rect 9920 4370 9990 4380
rect 2920 4360 2960 4370
rect 3040 4360 3080 4370
rect 3240 4360 3320 4370
rect 4560 4360 4600 4370
rect 4760 4360 4880 4370
rect 5400 4360 5480 4370
rect 5960 4360 6480 4370
rect 7400 4360 7440 4370
rect 7800 4360 7880 4370
rect 8520 4360 8680 4370
rect 9840 4360 9880 4370
rect 9920 4360 9990 4370
rect 2920 4350 2960 4360
rect 3040 4350 3080 4360
rect 3240 4350 3320 4360
rect 4560 4350 4600 4360
rect 4760 4350 4880 4360
rect 5400 4350 5480 4360
rect 5960 4350 6480 4360
rect 7400 4350 7440 4360
rect 7800 4350 7880 4360
rect 8520 4350 8680 4360
rect 9840 4350 9880 4360
rect 9920 4350 9990 4360
rect 2920 4340 2960 4350
rect 3040 4340 3080 4350
rect 3240 4340 3320 4350
rect 4560 4340 4600 4350
rect 4760 4340 4880 4350
rect 5400 4340 5480 4350
rect 5960 4340 6480 4350
rect 7400 4340 7440 4350
rect 7800 4340 7880 4350
rect 8520 4340 8680 4350
rect 9840 4340 9880 4350
rect 9920 4340 9990 4350
rect 3000 4330 3040 4340
rect 3160 4330 3240 4340
rect 3280 4330 3320 4340
rect 4560 4330 4600 4340
rect 4880 4330 4920 4340
rect 5320 4330 5360 4340
rect 5440 4330 5480 4340
rect 6120 4330 6480 4340
rect 8600 4330 8680 4340
rect 8840 4330 8880 4340
rect 3000 4320 3040 4330
rect 3160 4320 3240 4330
rect 3280 4320 3320 4330
rect 4560 4320 4600 4330
rect 4880 4320 4920 4330
rect 5320 4320 5360 4330
rect 5440 4320 5480 4330
rect 6120 4320 6480 4330
rect 8600 4320 8680 4330
rect 8840 4320 8880 4330
rect 3000 4310 3040 4320
rect 3160 4310 3240 4320
rect 3280 4310 3320 4320
rect 4560 4310 4600 4320
rect 4880 4310 4920 4320
rect 5320 4310 5360 4320
rect 5440 4310 5480 4320
rect 6120 4310 6480 4320
rect 8600 4310 8680 4320
rect 8840 4310 8880 4320
rect 3000 4300 3040 4310
rect 3160 4300 3240 4310
rect 3280 4300 3320 4310
rect 4560 4300 4600 4310
rect 4880 4300 4920 4310
rect 5320 4300 5360 4310
rect 5440 4300 5480 4310
rect 6120 4300 6480 4310
rect 8600 4300 8680 4310
rect 8840 4300 8880 4310
rect 2920 4290 3000 4300
rect 3040 4290 3080 4300
rect 3120 4290 3200 4300
rect 4160 4290 4320 4300
rect 4520 4290 4560 4300
rect 4920 4290 4960 4300
rect 5440 4290 5520 4300
rect 5960 4290 6440 4300
rect 8520 4290 8640 4300
rect 8680 4290 8720 4300
rect 9760 4290 9800 4300
rect 2920 4280 3000 4290
rect 3040 4280 3080 4290
rect 3120 4280 3200 4290
rect 4160 4280 4320 4290
rect 4520 4280 4560 4290
rect 4920 4280 4960 4290
rect 5440 4280 5520 4290
rect 5960 4280 6440 4290
rect 8520 4280 8640 4290
rect 8680 4280 8720 4290
rect 9760 4280 9800 4290
rect 2920 4270 3000 4280
rect 3040 4270 3080 4280
rect 3120 4270 3200 4280
rect 4160 4270 4320 4280
rect 4520 4270 4560 4280
rect 4920 4270 4960 4280
rect 5440 4270 5520 4280
rect 5960 4270 6440 4280
rect 8520 4270 8640 4280
rect 8680 4270 8720 4280
rect 9760 4270 9800 4280
rect 2920 4260 3000 4270
rect 3040 4260 3080 4270
rect 3120 4260 3200 4270
rect 4160 4260 4320 4270
rect 4520 4260 4560 4270
rect 4920 4260 4960 4270
rect 5440 4260 5520 4270
rect 5960 4260 6440 4270
rect 8520 4260 8640 4270
rect 8680 4260 8720 4270
rect 9760 4260 9800 4270
rect 2880 4250 2960 4260
rect 3040 4250 3240 4260
rect 4320 4250 4360 4260
rect 4920 4250 5000 4260
rect 5480 4250 5520 4260
rect 6000 4250 6280 4260
rect 6320 4250 6360 4260
rect 6520 4250 6560 4260
rect 7120 4250 7160 4260
rect 7240 4250 7440 4260
rect 8440 4250 8520 4260
rect 9360 4250 9400 4260
rect 9720 4250 9760 4260
rect 9800 4250 9840 4260
rect 2880 4240 2960 4250
rect 3040 4240 3240 4250
rect 4320 4240 4360 4250
rect 4920 4240 5000 4250
rect 5480 4240 5520 4250
rect 6000 4240 6280 4250
rect 6320 4240 6360 4250
rect 6520 4240 6560 4250
rect 7120 4240 7160 4250
rect 7240 4240 7440 4250
rect 8440 4240 8520 4250
rect 9360 4240 9400 4250
rect 9720 4240 9760 4250
rect 9800 4240 9840 4250
rect 2880 4230 2960 4240
rect 3040 4230 3240 4240
rect 4320 4230 4360 4240
rect 4920 4230 5000 4240
rect 5480 4230 5520 4240
rect 6000 4230 6280 4240
rect 6320 4230 6360 4240
rect 6520 4230 6560 4240
rect 7120 4230 7160 4240
rect 7240 4230 7440 4240
rect 8440 4230 8520 4240
rect 9360 4230 9400 4240
rect 9720 4230 9760 4240
rect 9800 4230 9840 4240
rect 2880 4220 2960 4230
rect 3040 4220 3240 4230
rect 4320 4220 4360 4230
rect 4920 4220 5000 4230
rect 5480 4220 5520 4230
rect 6000 4220 6280 4230
rect 6320 4220 6360 4230
rect 6520 4220 6560 4230
rect 7120 4220 7160 4230
rect 7240 4220 7440 4230
rect 8440 4220 8520 4230
rect 9360 4220 9400 4230
rect 9720 4220 9760 4230
rect 9800 4220 9840 4230
rect 3040 4210 3240 4220
rect 4120 4210 4160 4220
rect 4360 4210 4400 4220
rect 4440 4210 4480 4220
rect 4960 4210 5000 4220
rect 5480 4210 5560 4220
rect 6480 4210 6560 4220
rect 7240 4210 7280 4220
rect 8800 4210 8840 4220
rect 9760 4210 9840 4220
rect 3040 4200 3240 4210
rect 4120 4200 4160 4210
rect 4360 4200 4400 4210
rect 4440 4200 4480 4210
rect 4960 4200 5000 4210
rect 5480 4200 5560 4210
rect 6480 4200 6560 4210
rect 7240 4200 7280 4210
rect 8800 4200 8840 4210
rect 9760 4200 9840 4210
rect 3040 4190 3240 4200
rect 4120 4190 4160 4200
rect 4360 4190 4400 4200
rect 4440 4190 4480 4200
rect 4960 4190 5000 4200
rect 5480 4190 5560 4200
rect 6480 4190 6560 4200
rect 7240 4190 7280 4200
rect 8800 4190 8840 4200
rect 9760 4190 9840 4200
rect 3040 4180 3240 4190
rect 4120 4180 4160 4190
rect 4360 4180 4400 4190
rect 4440 4180 4480 4190
rect 4960 4180 5000 4190
rect 5480 4180 5560 4190
rect 6480 4180 6560 4190
rect 7240 4180 7280 4190
rect 8800 4180 8840 4190
rect 9760 4180 9840 4190
rect 2880 4170 2960 4180
rect 3000 4170 3120 4180
rect 3160 4170 3200 4180
rect 4080 4170 4120 4180
rect 4640 4170 4720 4180
rect 5000 4170 5040 4180
rect 5400 4170 5440 4180
rect 5480 4170 5520 4180
rect 5560 4170 5600 4180
rect 6440 4170 6520 4180
rect 7240 4170 7280 4180
rect 7320 4170 7360 4180
rect 9280 4170 9320 4180
rect 9840 4170 9880 4180
rect 2880 4160 2960 4170
rect 3000 4160 3120 4170
rect 3160 4160 3200 4170
rect 4080 4160 4120 4170
rect 4640 4160 4720 4170
rect 5000 4160 5040 4170
rect 5400 4160 5440 4170
rect 5480 4160 5520 4170
rect 5560 4160 5600 4170
rect 6440 4160 6520 4170
rect 7240 4160 7280 4170
rect 7320 4160 7360 4170
rect 9280 4160 9320 4170
rect 9840 4160 9880 4170
rect 2880 4150 2960 4160
rect 3000 4150 3120 4160
rect 3160 4150 3200 4160
rect 4080 4150 4120 4160
rect 4640 4150 4720 4160
rect 5000 4150 5040 4160
rect 5400 4150 5440 4160
rect 5480 4150 5520 4160
rect 5560 4150 5600 4160
rect 6440 4150 6520 4160
rect 7240 4150 7280 4160
rect 7320 4150 7360 4160
rect 9280 4150 9320 4160
rect 9840 4150 9880 4160
rect 2880 4140 2960 4150
rect 3000 4140 3120 4150
rect 3160 4140 3200 4150
rect 4080 4140 4120 4150
rect 4640 4140 4720 4150
rect 5000 4140 5040 4150
rect 5400 4140 5440 4150
rect 5480 4140 5520 4150
rect 5560 4140 5600 4150
rect 6440 4140 6520 4150
rect 7240 4140 7280 4150
rect 7320 4140 7360 4150
rect 9280 4140 9320 4150
rect 9840 4140 9880 4150
rect 2960 4130 3000 4140
rect 3040 4130 3080 4140
rect 3120 4130 3240 4140
rect 4560 4130 4720 4140
rect 4920 4130 5080 4140
rect 5600 4130 5640 4140
rect 6400 4130 6480 4140
rect 9880 4130 9920 4140
rect 9960 4130 9990 4140
rect 2960 4120 3000 4130
rect 3040 4120 3080 4130
rect 3120 4120 3240 4130
rect 4560 4120 4720 4130
rect 4920 4120 5080 4130
rect 5600 4120 5640 4130
rect 6400 4120 6480 4130
rect 9880 4120 9920 4130
rect 9960 4120 9990 4130
rect 2960 4110 3000 4120
rect 3040 4110 3080 4120
rect 3120 4110 3240 4120
rect 4560 4110 4720 4120
rect 4920 4110 5080 4120
rect 5600 4110 5640 4120
rect 6400 4110 6480 4120
rect 9880 4110 9920 4120
rect 9960 4110 9990 4120
rect 2960 4100 3000 4110
rect 3040 4100 3080 4110
rect 3120 4100 3240 4110
rect 4560 4100 4720 4110
rect 4920 4100 5080 4110
rect 5600 4100 5640 4110
rect 6400 4100 6480 4110
rect 9880 4100 9920 4110
rect 9960 4100 9990 4110
rect 3080 4090 3160 4100
rect 4040 4090 4080 4100
rect 4560 4090 4640 4100
rect 4800 4090 4840 4100
rect 5080 4090 5120 4100
rect 6360 4090 6440 4100
rect 7600 4090 7640 4100
rect 9920 4090 9990 4100
rect 3080 4080 3160 4090
rect 4040 4080 4080 4090
rect 4560 4080 4640 4090
rect 4800 4080 4840 4090
rect 5080 4080 5120 4090
rect 6360 4080 6440 4090
rect 7600 4080 7640 4090
rect 9920 4080 9990 4090
rect 3080 4070 3160 4080
rect 4040 4070 4080 4080
rect 4560 4070 4640 4080
rect 4800 4070 4840 4080
rect 5080 4070 5120 4080
rect 6360 4070 6440 4080
rect 7600 4070 7640 4080
rect 9920 4070 9990 4080
rect 3080 4060 3160 4070
rect 4040 4060 4080 4070
rect 4560 4060 4640 4070
rect 4800 4060 4840 4070
rect 5080 4060 5120 4070
rect 6360 4060 6440 4070
rect 7600 4060 7640 4070
rect 9920 4060 9990 4070
rect 2960 4050 3000 4060
rect 3040 4050 3080 4060
rect 4560 4050 4640 4060
rect 5080 4050 5120 4060
rect 5720 4050 5760 4060
rect 6280 4050 6400 4060
rect 8520 4050 8680 4060
rect 2960 4040 3000 4050
rect 3040 4040 3080 4050
rect 4560 4040 4640 4050
rect 5080 4040 5120 4050
rect 5720 4040 5760 4050
rect 6280 4040 6400 4050
rect 8520 4040 8680 4050
rect 2960 4030 3000 4040
rect 3040 4030 3080 4040
rect 4560 4030 4640 4040
rect 5080 4030 5120 4040
rect 5720 4030 5760 4040
rect 6280 4030 6400 4040
rect 8520 4030 8680 4040
rect 2960 4020 3000 4030
rect 3040 4020 3080 4030
rect 4560 4020 4640 4030
rect 5080 4020 5120 4030
rect 5720 4020 5760 4030
rect 6280 4020 6400 4030
rect 8520 4020 8680 4030
rect 3080 4010 3120 4020
rect 4000 4010 4040 4020
rect 4560 4010 4640 4020
rect 4680 4010 4720 4020
rect 5120 4010 5160 4020
rect 5480 4010 5520 4020
rect 5760 4010 6000 4020
rect 6200 4010 6400 4020
rect 7160 4010 7200 4020
rect 8320 4010 8360 4020
rect 8480 4010 8560 4020
rect 8640 4010 8760 4020
rect 3080 4000 3120 4010
rect 4000 4000 4040 4010
rect 4560 4000 4640 4010
rect 4680 4000 4720 4010
rect 5120 4000 5160 4010
rect 5480 4000 5520 4010
rect 5760 4000 6000 4010
rect 6200 4000 6400 4010
rect 7160 4000 7200 4010
rect 8320 4000 8360 4010
rect 8480 4000 8560 4010
rect 8640 4000 8760 4010
rect 3080 3990 3120 4000
rect 4000 3990 4040 4000
rect 4560 3990 4640 4000
rect 4680 3990 4720 4000
rect 5120 3990 5160 4000
rect 5480 3990 5520 4000
rect 5760 3990 6000 4000
rect 6200 3990 6400 4000
rect 7160 3990 7200 4000
rect 8320 3990 8360 4000
rect 8480 3990 8560 4000
rect 8640 3990 8760 4000
rect 3080 3980 3120 3990
rect 4000 3980 4040 3990
rect 4560 3980 4640 3990
rect 4680 3980 4720 3990
rect 5120 3980 5160 3990
rect 5480 3980 5520 3990
rect 5760 3980 6000 3990
rect 6200 3980 6400 3990
rect 7160 3980 7200 3990
rect 8320 3980 8360 3990
rect 8480 3980 8560 3990
rect 8640 3980 8760 3990
rect 3120 3970 3200 3980
rect 3240 3970 3280 3980
rect 3960 3970 4000 3980
rect 4160 3970 4280 3980
rect 4720 3970 4800 3980
rect 5120 3970 5160 3980
rect 5400 3970 5440 3980
rect 6000 3970 6240 3980
rect 6320 3970 6400 3980
rect 7840 3970 7880 3980
rect 8160 3970 8240 3980
rect 8280 3970 8320 3980
rect 8400 3970 8440 3980
rect 3120 3960 3200 3970
rect 3240 3960 3280 3970
rect 3960 3960 4000 3970
rect 4160 3960 4280 3970
rect 4720 3960 4800 3970
rect 5120 3960 5160 3970
rect 5400 3960 5440 3970
rect 6000 3960 6240 3970
rect 6320 3960 6400 3970
rect 7840 3960 7880 3970
rect 8160 3960 8240 3970
rect 8280 3960 8320 3970
rect 8400 3960 8440 3970
rect 3120 3950 3200 3960
rect 3240 3950 3280 3960
rect 3960 3950 4000 3960
rect 4160 3950 4280 3960
rect 4720 3950 4800 3960
rect 5120 3950 5160 3960
rect 5400 3950 5440 3960
rect 6000 3950 6240 3960
rect 6320 3950 6400 3960
rect 7840 3950 7880 3960
rect 8160 3950 8240 3960
rect 8280 3950 8320 3960
rect 8400 3950 8440 3960
rect 3120 3940 3200 3950
rect 3240 3940 3280 3950
rect 3960 3940 4000 3950
rect 4160 3940 4280 3950
rect 4720 3940 4800 3950
rect 5120 3940 5160 3950
rect 5400 3940 5440 3950
rect 6000 3940 6240 3950
rect 6320 3940 6400 3950
rect 7840 3940 7880 3950
rect 8160 3940 8240 3950
rect 8280 3940 8320 3950
rect 8400 3940 8440 3950
rect 2920 3930 2960 3940
rect 3040 3930 3200 3940
rect 3920 3930 3960 3940
rect 4120 3930 4200 3940
rect 4280 3930 4320 3940
rect 5160 3930 5200 3940
rect 6320 3930 6400 3940
rect 7960 3930 8000 3940
rect 8040 3930 8080 3940
rect 8120 3930 8200 3940
rect 8280 3930 8320 3940
rect 8560 3930 8640 3940
rect 9640 3930 9720 3940
rect 2920 3920 2960 3930
rect 3040 3920 3200 3930
rect 3920 3920 3960 3930
rect 4120 3920 4200 3930
rect 4280 3920 4320 3930
rect 5160 3920 5200 3930
rect 6320 3920 6400 3930
rect 7960 3920 8000 3930
rect 8040 3920 8080 3930
rect 8120 3920 8200 3930
rect 8280 3920 8320 3930
rect 8560 3920 8640 3930
rect 9640 3920 9720 3930
rect 2920 3910 2960 3920
rect 3040 3910 3200 3920
rect 3920 3910 3960 3920
rect 4120 3910 4200 3920
rect 4280 3910 4320 3920
rect 5160 3910 5200 3920
rect 6320 3910 6400 3920
rect 7960 3910 8000 3920
rect 8040 3910 8080 3920
rect 8120 3910 8200 3920
rect 8280 3910 8320 3920
rect 8560 3910 8640 3920
rect 9640 3910 9720 3920
rect 2920 3900 2960 3910
rect 3040 3900 3200 3910
rect 3920 3900 3960 3910
rect 4120 3900 4200 3910
rect 4280 3900 4320 3910
rect 5160 3900 5200 3910
rect 6320 3900 6400 3910
rect 7960 3900 8000 3910
rect 8040 3900 8080 3910
rect 8120 3900 8200 3910
rect 8280 3900 8320 3910
rect 8560 3900 8640 3910
rect 9640 3900 9720 3910
rect 2880 3890 3160 3900
rect 3880 3890 3920 3900
rect 4080 3890 4120 3900
rect 4280 3890 4320 3900
rect 5200 3890 5240 3900
rect 6320 3890 6440 3900
rect 7120 3890 7160 3900
rect 8040 3890 8080 3900
rect 8280 3890 8320 3900
rect 8520 3890 8600 3900
rect 9480 3890 9600 3900
rect 9680 3890 9720 3900
rect 2880 3880 3160 3890
rect 3880 3880 3920 3890
rect 4080 3880 4120 3890
rect 4280 3880 4320 3890
rect 5200 3880 5240 3890
rect 6320 3880 6440 3890
rect 7120 3880 7160 3890
rect 8040 3880 8080 3890
rect 8280 3880 8320 3890
rect 8520 3880 8600 3890
rect 9480 3880 9600 3890
rect 9680 3880 9720 3890
rect 2880 3870 3160 3880
rect 3880 3870 3920 3880
rect 4080 3870 4120 3880
rect 4280 3870 4320 3880
rect 5200 3870 5240 3880
rect 6320 3870 6440 3880
rect 7120 3870 7160 3880
rect 8040 3870 8080 3880
rect 8280 3870 8320 3880
rect 8520 3870 8600 3880
rect 9480 3870 9600 3880
rect 9680 3870 9720 3880
rect 2880 3860 3160 3870
rect 3880 3860 3920 3870
rect 4080 3860 4120 3870
rect 4280 3860 4320 3870
rect 5200 3860 5240 3870
rect 6320 3860 6440 3870
rect 7120 3860 7160 3870
rect 8040 3860 8080 3870
rect 8280 3860 8320 3870
rect 8520 3860 8600 3870
rect 9480 3860 9600 3870
rect 9680 3860 9720 3870
rect 2880 3850 3160 3860
rect 4080 3850 4120 3860
rect 4280 3850 4320 3860
rect 5200 3850 5240 3860
rect 6320 3850 6520 3860
rect 2880 3840 3160 3850
rect 4080 3840 4120 3850
rect 4280 3840 4320 3850
rect 5200 3840 5240 3850
rect 6320 3840 6520 3850
rect 2880 3830 3160 3840
rect 4080 3830 4120 3840
rect 4280 3830 4320 3840
rect 5200 3830 5240 3840
rect 6320 3830 6520 3840
rect 2880 3820 3160 3830
rect 4080 3820 4120 3830
rect 4280 3820 4320 3830
rect 5200 3820 5240 3830
rect 6320 3820 6520 3830
rect 2920 3810 3000 3820
rect 3080 3810 3200 3820
rect 4040 3810 4080 3820
rect 5240 3810 5280 3820
rect 6280 3810 6520 3820
rect 8120 3810 8160 3820
rect 8200 3810 8280 3820
rect 9600 3810 9640 3820
rect 9720 3810 9840 3820
rect 2920 3800 3000 3810
rect 3080 3800 3200 3810
rect 4040 3800 4080 3810
rect 5240 3800 5280 3810
rect 6280 3800 6520 3810
rect 8120 3800 8160 3810
rect 8200 3800 8280 3810
rect 9600 3800 9640 3810
rect 9720 3800 9840 3810
rect 2920 3790 3000 3800
rect 3080 3790 3200 3800
rect 4040 3790 4080 3800
rect 5240 3790 5280 3800
rect 6280 3790 6520 3800
rect 8120 3790 8160 3800
rect 8200 3790 8280 3800
rect 9600 3790 9640 3800
rect 9720 3790 9840 3800
rect 2920 3780 3000 3790
rect 3080 3780 3200 3790
rect 4040 3780 4080 3790
rect 5240 3780 5280 3790
rect 6280 3780 6520 3790
rect 8120 3780 8160 3790
rect 8200 3780 8280 3790
rect 9600 3780 9640 3790
rect 9720 3780 9840 3790
rect 2920 3770 2960 3780
rect 3080 3770 3200 3780
rect 3880 3770 3920 3780
rect 4120 3770 4160 3780
rect 5240 3770 5280 3780
rect 6320 3770 6520 3780
rect 7040 3770 7080 3780
rect 8160 3770 8320 3780
rect 9720 3770 9840 3780
rect 2920 3760 2960 3770
rect 3080 3760 3200 3770
rect 3880 3760 3920 3770
rect 4120 3760 4160 3770
rect 5240 3760 5280 3770
rect 6320 3760 6520 3770
rect 7040 3760 7080 3770
rect 8160 3760 8320 3770
rect 9720 3760 9840 3770
rect 2920 3750 2960 3760
rect 3080 3750 3200 3760
rect 3880 3750 3920 3760
rect 4120 3750 4160 3760
rect 5240 3750 5280 3760
rect 6320 3750 6520 3760
rect 7040 3750 7080 3760
rect 8160 3750 8320 3760
rect 9720 3750 9840 3760
rect 2920 3740 2960 3750
rect 3080 3740 3200 3750
rect 3880 3740 3920 3750
rect 4120 3740 4160 3750
rect 5240 3740 5280 3750
rect 6320 3740 6520 3750
rect 7040 3740 7080 3750
rect 8160 3740 8320 3750
rect 9720 3740 9840 3750
rect 2880 3730 3000 3740
rect 3120 3730 3160 3740
rect 3280 3730 3320 3740
rect 3880 3730 3920 3740
rect 4200 3730 4240 3740
rect 4840 3730 4880 3740
rect 6440 3730 6520 3740
rect 8160 3730 8440 3740
rect 8560 3730 8600 3740
rect 2880 3720 3000 3730
rect 3120 3720 3160 3730
rect 3280 3720 3320 3730
rect 3880 3720 3920 3730
rect 4200 3720 4240 3730
rect 4840 3720 4880 3730
rect 6440 3720 6520 3730
rect 8160 3720 8440 3730
rect 8560 3720 8600 3730
rect 2880 3710 3000 3720
rect 3120 3710 3160 3720
rect 3280 3710 3320 3720
rect 3880 3710 3920 3720
rect 4200 3710 4240 3720
rect 4840 3710 4880 3720
rect 6440 3710 6520 3720
rect 8160 3710 8440 3720
rect 8560 3710 8600 3720
rect 2880 3700 3000 3710
rect 3120 3700 3160 3710
rect 3280 3700 3320 3710
rect 3880 3700 3920 3710
rect 4200 3700 4240 3710
rect 4840 3700 4880 3710
rect 6440 3700 6520 3710
rect 8160 3700 8440 3710
rect 8560 3700 8600 3710
rect 3040 3690 3080 3700
rect 3280 3690 3320 3700
rect 3880 3690 4000 3700
rect 4120 3690 4160 3700
rect 4880 3690 5000 3700
rect 5280 3690 5320 3700
rect 6480 3690 6560 3700
rect 8560 3690 8600 3700
rect 3040 3680 3080 3690
rect 3280 3680 3320 3690
rect 3880 3680 4000 3690
rect 4120 3680 4160 3690
rect 4880 3680 5000 3690
rect 5280 3680 5320 3690
rect 6480 3680 6560 3690
rect 8560 3680 8600 3690
rect 3040 3670 3080 3680
rect 3280 3670 3320 3680
rect 3880 3670 4000 3680
rect 4120 3670 4160 3680
rect 4880 3670 5000 3680
rect 5280 3670 5320 3680
rect 6480 3670 6560 3680
rect 8560 3670 8600 3680
rect 3040 3660 3080 3670
rect 3280 3660 3320 3670
rect 3880 3660 4000 3670
rect 4120 3660 4160 3670
rect 4880 3660 5000 3670
rect 5280 3660 5320 3670
rect 6480 3660 6560 3670
rect 8560 3660 8600 3670
rect 3120 3650 3240 3660
rect 3280 3650 3320 3660
rect 4960 3650 5120 3660
rect 5280 3650 5320 3660
rect 6440 3650 6520 3660
rect 8200 3650 8240 3660
rect 8360 3650 8400 3660
rect 8520 3650 8560 3660
rect 9560 3650 9640 3660
rect 3120 3640 3240 3650
rect 3280 3640 3320 3650
rect 4960 3640 5120 3650
rect 5280 3640 5320 3650
rect 6440 3640 6520 3650
rect 8200 3640 8240 3650
rect 8360 3640 8400 3650
rect 8520 3640 8560 3650
rect 9560 3640 9640 3650
rect 3120 3630 3240 3640
rect 3280 3630 3320 3640
rect 4960 3630 5120 3640
rect 5280 3630 5320 3640
rect 6440 3630 6520 3640
rect 8200 3630 8240 3640
rect 8360 3630 8400 3640
rect 8520 3630 8560 3640
rect 9560 3630 9640 3640
rect 3120 3620 3240 3630
rect 3280 3620 3320 3630
rect 4960 3620 5120 3630
rect 5280 3620 5320 3630
rect 6440 3620 6520 3630
rect 8200 3620 8240 3630
rect 8360 3620 8400 3630
rect 8520 3620 8560 3630
rect 9560 3620 9640 3630
rect 3240 3610 3360 3620
rect 5040 3610 5120 3620
rect 6440 3610 6520 3620
rect 6920 3610 6960 3620
rect 8240 3610 8280 3620
rect 8360 3610 8400 3620
rect 8480 3610 8520 3620
rect 9480 3610 9560 3620
rect 3240 3600 3360 3610
rect 5040 3600 5120 3610
rect 6440 3600 6520 3610
rect 6920 3600 6960 3610
rect 8240 3600 8280 3610
rect 8360 3600 8400 3610
rect 8480 3600 8520 3610
rect 9480 3600 9560 3610
rect 3240 3590 3360 3600
rect 5040 3590 5120 3600
rect 6440 3590 6520 3600
rect 6920 3590 6960 3600
rect 8240 3590 8280 3600
rect 8360 3590 8400 3600
rect 8480 3590 8520 3600
rect 9480 3590 9560 3600
rect 3240 3580 3360 3590
rect 5040 3580 5120 3590
rect 6440 3580 6520 3590
rect 6920 3580 6960 3590
rect 8240 3580 8280 3590
rect 8360 3580 8400 3590
rect 8480 3580 8520 3590
rect 9480 3580 9560 3590
rect 3240 3570 3280 3580
rect 3360 3570 3400 3580
rect 3920 3570 3960 3580
rect 4720 3570 4800 3580
rect 5080 3570 5120 3580
rect 6360 3570 6520 3580
rect 8400 3570 8440 3580
rect 9400 3570 9440 3580
rect 9480 3570 9520 3580
rect 3240 3560 3280 3570
rect 3360 3560 3400 3570
rect 3920 3560 3960 3570
rect 4720 3560 4800 3570
rect 5080 3560 5120 3570
rect 6360 3560 6520 3570
rect 8400 3560 8440 3570
rect 9400 3560 9440 3570
rect 9480 3560 9520 3570
rect 3240 3550 3280 3560
rect 3360 3550 3400 3560
rect 3920 3550 3960 3560
rect 4720 3550 4800 3560
rect 5080 3550 5120 3560
rect 6360 3550 6520 3560
rect 8400 3550 8440 3560
rect 9400 3550 9440 3560
rect 9480 3550 9520 3560
rect 3240 3540 3280 3550
rect 3360 3540 3400 3550
rect 3920 3540 3960 3550
rect 4720 3540 4800 3550
rect 5080 3540 5120 3550
rect 6360 3540 6520 3550
rect 8400 3540 8440 3550
rect 9400 3540 9440 3550
rect 9480 3540 9520 3550
rect 3280 3530 3320 3540
rect 3920 3530 4000 3540
rect 4680 3530 4760 3540
rect 5000 3530 5080 3540
rect 6360 3530 6480 3540
rect 8320 3530 8360 3540
rect 8400 3530 8440 3540
rect 9240 3530 9440 3540
rect 3280 3520 3320 3530
rect 3920 3520 4000 3530
rect 4680 3520 4760 3530
rect 5000 3520 5080 3530
rect 6360 3520 6480 3530
rect 8320 3520 8360 3530
rect 8400 3520 8440 3530
rect 9240 3520 9440 3530
rect 3280 3510 3320 3520
rect 3920 3510 4000 3520
rect 4680 3510 4760 3520
rect 5000 3510 5080 3520
rect 6360 3510 6480 3520
rect 8320 3510 8360 3520
rect 8400 3510 8440 3520
rect 9240 3510 9440 3520
rect 3280 3500 3320 3510
rect 3920 3500 4000 3510
rect 4680 3500 4760 3510
rect 5000 3500 5080 3510
rect 6360 3500 6480 3510
rect 8320 3500 8360 3510
rect 8400 3500 8440 3510
rect 9240 3500 9440 3510
rect 2680 3490 2760 3500
rect 3400 3490 3440 3500
rect 3960 3490 4000 3500
rect 4280 3490 4400 3500
rect 4480 3490 4760 3500
rect 6320 3490 6480 3500
rect 8400 3490 8480 3500
rect 9200 3490 9240 3500
rect 9320 3490 9360 3500
rect 9560 3490 9600 3500
rect 2680 3480 2760 3490
rect 3400 3480 3440 3490
rect 3960 3480 4000 3490
rect 4280 3480 4400 3490
rect 4480 3480 4760 3490
rect 6320 3480 6480 3490
rect 8400 3480 8480 3490
rect 9200 3480 9240 3490
rect 9320 3480 9360 3490
rect 9560 3480 9600 3490
rect 2680 3470 2760 3480
rect 3400 3470 3440 3480
rect 3960 3470 4000 3480
rect 4280 3470 4400 3480
rect 4480 3470 4760 3480
rect 6320 3470 6480 3480
rect 8400 3470 8480 3480
rect 9200 3470 9240 3480
rect 9320 3470 9360 3480
rect 9560 3470 9600 3480
rect 2680 3460 2760 3470
rect 3400 3460 3440 3470
rect 3960 3460 4000 3470
rect 4280 3460 4400 3470
rect 4480 3460 4760 3470
rect 6320 3460 6480 3470
rect 8400 3460 8480 3470
rect 9200 3460 9240 3470
rect 9320 3460 9360 3470
rect 9560 3460 9600 3470
rect 2880 3450 2920 3460
rect 3960 3450 4000 3460
rect 4280 3450 4440 3460
rect 4680 3450 4760 3460
rect 4880 3450 4920 3460
rect 5000 3450 5040 3460
rect 6280 3450 6440 3460
rect 8520 3450 8560 3460
rect 9160 3450 9200 3460
rect 9520 3450 9600 3460
rect 2880 3440 2920 3450
rect 3960 3440 4000 3450
rect 4280 3440 4440 3450
rect 4680 3440 4760 3450
rect 4880 3440 4920 3450
rect 5000 3440 5040 3450
rect 6280 3440 6440 3450
rect 8520 3440 8560 3450
rect 9160 3440 9200 3450
rect 9520 3440 9600 3450
rect 2880 3430 2920 3440
rect 3960 3430 4000 3440
rect 4280 3430 4440 3440
rect 4680 3430 4760 3440
rect 4880 3430 4920 3440
rect 5000 3430 5040 3440
rect 6280 3430 6440 3440
rect 8520 3430 8560 3440
rect 9160 3430 9200 3440
rect 9520 3430 9600 3440
rect 2880 3420 2920 3430
rect 3960 3420 4000 3430
rect 4280 3420 4440 3430
rect 4680 3420 4760 3430
rect 4880 3420 4920 3430
rect 5000 3420 5040 3430
rect 6280 3420 6440 3430
rect 8520 3420 8560 3430
rect 9160 3420 9200 3430
rect 9520 3420 9600 3430
rect 2200 3410 2240 3420
rect 2960 3410 3000 3420
rect 3960 3410 4000 3420
rect 4240 3410 4280 3420
rect 4320 3410 4360 3420
rect 4400 3410 4480 3420
rect 4560 3410 4840 3420
rect 4920 3410 5000 3420
rect 6200 3410 6400 3420
rect 9080 3410 9120 3420
rect 9160 3410 9200 3420
rect 9440 3410 9560 3420
rect 2200 3400 2240 3410
rect 2960 3400 3000 3410
rect 3960 3400 4000 3410
rect 4240 3400 4280 3410
rect 4320 3400 4360 3410
rect 4400 3400 4480 3410
rect 4560 3400 4840 3410
rect 4920 3400 5000 3410
rect 6200 3400 6400 3410
rect 9080 3400 9120 3410
rect 9160 3400 9200 3410
rect 9440 3400 9560 3410
rect 2200 3390 2240 3400
rect 2960 3390 3000 3400
rect 3960 3390 4000 3400
rect 4240 3390 4280 3400
rect 4320 3390 4360 3400
rect 4400 3390 4480 3400
rect 4560 3390 4840 3400
rect 4920 3390 5000 3400
rect 6200 3390 6400 3400
rect 9080 3390 9120 3400
rect 9160 3390 9200 3400
rect 9440 3390 9560 3400
rect 2200 3380 2240 3390
rect 2960 3380 3000 3390
rect 3960 3380 4000 3390
rect 4240 3380 4280 3390
rect 4320 3380 4360 3390
rect 4400 3380 4480 3390
rect 4560 3380 4840 3390
rect 4920 3380 5000 3390
rect 6200 3380 6400 3390
rect 9080 3380 9120 3390
rect 9160 3380 9200 3390
rect 9440 3380 9560 3390
rect 2160 3370 2200 3380
rect 3040 3370 3080 3380
rect 4000 3370 4040 3380
rect 4240 3370 4280 3380
rect 4320 3370 4360 3380
rect 4600 3370 4720 3380
rect 5280 3370 5320 3380
rect 6160 3370 6360 3380
rect 9440 3370 9520 3380
rect 9720 3370 9760 3380
rect 2160 3360 2200 3370
rect 3040 3360 3080 3370
rect 4000 3360 4040 3370
rect 4240 3360 4280 3370
rect 4320 3360 4360 3370
rect 4600 3360 4720 3370
rect 5280 3360 5320 3370
rect 6160 3360 6360 3370
rect 9440 3360 9520 3370
rect 9720 3360 9760 3370
rect 2160 3350 2200 3360
rect 3040 3350 3080 3360
rect 4000 3350 4040 3360
rect 4240 3350 4280 3360
rect 4320 3350 4360 3360
rect 4600 3350 4720 3360
rect 5280 3350 5320 3360
rect 6160 3350 6360 3360
rect 9440 3350 9520 3360
rect 9720 3350 9760 3360
rect 2160 3340 2200 3350
rect 3040 3340 3080 3350
rect 4000 3340 4040 3350
rect 4240 3340 4280 3350
rect 4320 3340 4360 3350
rect 4600 3340 4720 3350
rect 5280 3340 5320 3350
rect 6160 3340 6360 3350
rect 9440 3340 9520 3350
rect 9720 3340 9760 3350
rect 2120 3330 2160 3340
rect 3080 3330 3120 3340
rect 4040 3330 4240 3340
rect 4320 3330 4360 3340
rect 4560 3330 4600 3340
rect 4800 3330 4840 3340
rect 5280 3330 5320 3340
rect 6160 3330 6320 3340
rect 9040 3330 9080 3340
rect 9400 3330 9480 3340
rect 9680 3330 9760 3340
rect 2120 3320 2160 3330
rect 3080 3320 3120 3330
rect 4040 3320 4240 3330
rect 4320 3320 4360 3330
rect 4560 3320 4600 3330
rect 4800 3320 4840 3330
rect 5280 3320 5320 3330
rect 6160 3320 6320 3330
rect 9040 3320 9080 3330
rect 9400 3320 9480 3330
rect 9680 3320 9760 3330
rect 2120 3310 2160 3320
rect 3080 3310 3120 3320
rect 4040 3310 4240 3320
rect 4320 3310 4360 3320
rect 4560 3310 4600 3320
rect 4800 3310 4840 3320
rect 5280 3310 5320 3320
rect 6160 3310 6320 3320
rect 9040 3310 9080 3320
rect 9400 3310 9480 3320
rect 9680 3310 9760 3320
rect 2120 3300 2160 3310
rect 3080 3300 3120 3310
rect 4040 3300 4240 3310
rect 4320 3300 4360 3310
rect 4560 3300 4600 3310
rect 4800 3300 4840 3310
rect 5280 3300 5320 3310
rect 6160 3300 6320 3310
rect 9040 3300 9080 3310
rect 9400 3300 9480 3310
rect 9680 3300 9760 3310
rect 2080 3290 2120 3300
rect 4080 3290 4240 3300
rect 4320 3290 4360 3300
rect 4480 3290 4520 3300
rect 4720 3290 4760 3300
rect 4960 3290 5000 3300
rect 5280 3290 5320 3300
rect 6160 3290 6240 3300
rect 6640 3290 6680 3300
rect 8440 3290 8480 3300
rect 9040 3290 9120 3300
rect 9360 3290 9440 3300
rect 9600 3290 9640 3300
rect 9680 3290 9720 3300
rect 2080 3280 2120 3290
rect 4080 3280 4240 3290
rect 4320 3280 4360 3290
rect 4480 3280 4520 3290
rect 4720 3280 4760 3290
rect 4960 3280 5000 3290
rect 5280 3280 5320 3290
rect 6160 3280 6240 3290
rect 6640 3280 6680 3290
rect 8440 3280 8480 3290
rect 9040 3280 9120 3290
rect 9360 3280 9440 3290
rect 9600 3280 9640 3290
rect 9680 3280 9720 3290
rect 2080 3270 2120 3280
rect 4080 3270 4240 3280
rect 4320 3270 4360 3280
rect 4480 3270 4520 3280
rect 4720 3270 4760 3280
rect 4960 3270 5000 3280
rect 5280 3270 5320 3280
rect 6160 3270 6240 3280
rect 6640 3270 6680 3280
rect 8440 3270 8480 3280
rect 9040 3270 9120 3280
rect 9360 3270 9440 3280
rect 9600 3270 9640 3280
rect 9680 3270 9720 3280
rect 2080 3260 2120 3270
rect 4080 3260 4240 3270
rect 4320 3260 4360 3270
rect 4480 3260 4520 3270
rect 4720 3260 4760 3270
rect 4960 3260 5000 3270
rect 5280 3260 5320 3270
rect 6160 3260 6240 3270
rect 6640 3260 6680 3270
rect 8440 3260 8480 3270
rect 9040 3260 9120 3270
rect 9360 3260 9440 3270
rect 9600 3260 9640 3270
rect 9680 3260 9720 3270
rect 2080 3250 2120 3260
rect 3560 3250 3600 3260
rect 4120 3250 4280 3260
rect 4360 3250 4400 3260
rect 4640 3250 4680 3260
rect 4920 3250 5000 3260
rect 6200 3250 6240 3260
rect 6480 3250 6520 3260
rect 6600 3250 6640 3260
rect 9080 3250 9120 3260
rect 9400 3250 9440 3260
rect 9520 3250 9680 3260
rect 2080 3240 2120 3250
rect 3560 3240 3600 3250
rect 4120 3240 4280 3250
rect 4360 3240 4400 3250
rect 4640 3240 4680 3250
rect 4920 3240 5000 3250
rect 6200 3240 6240 3250
rect 6480 3240 6520 3250
rect 6600 3240 6640 3250
rect 9080 3240 9120 3250
rect 9400 3240 9440 3250
rect 9520 3240 9680 3250
rect 2080 3230 2120 3240
rect 3560 3230 3600 3240
rect 4120 3230 4280 3240
rect 4360 3230 4400 3240
rect 4640 3230 4680 3240
rect 4920 3230 5000 3240
rect 6200 3230 6240 3240
rect 6480 3230 6520 3240
rect 6600 3230 6640 3240
rect 9080 3230 9120 3240
rect 9400 3230 9440 3240
rect 9520 3230 9680 3240
rect 2080 3220 2120 3230
rect 3560 3220 3600 3230
rect 4120 3220 4280 3230
rect 4360 3220 4400 3230
rect 4640 3220 4680 3230
rect 4920 3220 5000 3230
rect 6200 3220 6240 3230
rect 6480 3220 6520 3230
rect 6600 3220 6640 3230
rect 9080 3220 9120 3230
rect 9400 3220 9440 3230
rect 9520 3220 9680 3230
rect 4160 3210 4280 3220
rect 4520 3210 4600 3220
rect 4880 3210 4920 3220
rect 6200 3210 6280 3220
rect 6400 3210 6440 3220
rect 6600 3210 6640 3220
rect 8400 3210 8440 3220
rect 9040 3210 9080 3220
rect 9160 3210 9280 3220
rect 9320 3210 9400 3220
rect 9480 3210 9520 3220
rect 4160 3200 4280 3210
rect 4520 3200 4600 3210
rect 4880 3200 4920 3210
rect 6200 3200 6280 3210
rect 6400 3200 6440 3210
rect 6600 3200 6640 3210
rect 8400 3200 8440 3210
rect 9040 3200 9080 3210
rect 9160 3200 9280 3210
rect 9320 3200 9400 3210
rect 9480 3200 9520 3210
rect 4160 3190 4280 3200
rect 4520 3190 4600 3200
rect 4880 3190 4920 3200
rect 6200 3190 6280 3200
rect 6400 3190 6440 3200
rect 6600 3190 6640 3200
rect 8400 3190 8440 3200
rect 9040 3190 9080 3200
rect 9160 3190 9280 3200
rect 9320 3190 9400 3200
rect 9480 3190 9520 3200
rect 4160 3180 4280 3190
rect 4520 3180 4600 3190
rect 4880 3180 4920 3190
rect 6200 3180 6280 3190
rect 6400 3180 6440 3190
rect 6600 3180 6640 3190
rect 8400 3180 8440 3190
rect 9040 3180 9080 3190
rect 9160 3180 9280 3190
rect 9320 3180 9400 3190
rect 9480 3180 9520 3190
rect 2040 3170 2080 3180
rect 3160 3170 3200 3180
rect 4160 3170 4240 3180
rect 4320 3170 4400 3180
rect 4480 3170 4600 3180
rect 4920 3170 4960 3180
rect 5240 3170 5280 3180
rect 6240 3170 6320 3180
rect 6600 3170 6640 3180
rect 9000 3170 9080 3180
rect 9280 3170 9400 3180
rect 9440 3170 9480 3180
rect 9520 3170 9560 3180
rect 9920 3170 9960 3180
rect 2040 3160 2080 3170
rect 3160 3160 3200 3170
rect 4160 3160 4240 3170
rect 4320 3160 4400 3170
rect 4480 3160 4600 3170
rect 4920 3160 4960 3170
rect 5240 3160 5280 3170
rect 6240 3160 6320 3170
rect 6600 3160 6640 3170
rect 9000 3160 9080 3170
rect 9280 3160 9400 3170
rect 9440 3160 9480 3170
rect 9520 3160 9560 3170
rect 9920 3160 9960 3170
rect 2040 3150 2080 3160
rect 3160 3150 3200 3160
rect 4160 3150 4240 3160
rect 4320 3150 4400 3160
rect 4480 3150 4600 3160
rect 4920 3150 4960 3160
rect 5240 3150 5280 3160
rect 6240 3150 6320 3160
rect 6600 3150 6640 3160
rect 9000 3150 9080 3160
rect 9280 3150 9400 3160
rect 9440 3150 9480 3160
rect 9520 3150 9560 3160
rect 9920 3150 9960 3160
rect 2040 3140 2080 3150
rect 3160 3140 3200 3150
rect 4160 3140 4240 3150
rect 4320 3140 4400 3150
rect 4480 3140 4600 3150
rect 4920 3140 4960 3150
rect 5240 3140 5280 3150
rect 6240 3140 6320 3150
rect 6600 3140 6640 3150
rect 9000 3140 9080 3150
rect 9280 3140 9400 3150
rect 9440 3140 9480 3150
rect 9520 3140 9560 3150
rect 9920 3140 9960 3150
rect 2040 3130 2080 3140
rect 3160 3130 3200 3140
rect 4200 3130 4240 3140
rect 4520 3130 4600 3140
rect 4800 3130 4840 3140
rect 5240 3130 5280 3140
rect 6560 3130 6600 3140
rect 8360 3130 8400 3140
rect 8920 3130 8960 3140
rect 9040 3130 9080 3140
rect 9240 3130 9440 3140
rect 9520 3130 9560 3140
rect 9920 3130 9990 3140
rect 2040 3120 2080 3130
rect 3160 3120 3200 3130
rect 4200 3120 4240 3130
rect 4520 3120 4600 3130
rect 4800 3120 4840 3130
rect 5240 3120 5280 3130
rect 6560 3120 6600 3130
rect 8360 3120 8400 3130
rect 8920 3120 8960 3130
rect 9040 3120 9080 3130
rect 9240 3120 9440 3130
rect 9520 3120 9560 3130
rect 9920 3120 9990 3130
rect 2040 3110 2080 3120
rect 3160 3110 3200 3120
rect 4200 3110 4240 3120
rect 4520 3110 4600 3120
rect 4800 3110 4840 3120
rect 5240 3110 5280 3120
rect 6560 3110 6600 3120
rect 8360 3110 8400 3120
rect 8920 3110 8960 3120
rect 9040 3110 9080 3120
rect 9240 3110 9440 3120
rect 9520 3110 9560 3120
rect 9920 3110 9990 3120
rect 2040 3100 2080 3110
rect 3160 3100 3200 3110
rect 4200 3100 4240 3110
rect 4520 3100 4600 3110
rect 4800 3100 4840 3110
rect 5240 3100 5280 3110
rect 6560 3100 6600 3110
rect 8360 3100 8400 3110
rect 8920 3100 8960 3110
rect 9040 3100 9080 3110
rect 9240 3100 9440 3110
rect 9520 3100 9560 3110
rect 9920 3100 9990 3110
rect 2040 3090 2080 3100
rect 3160 3090 3200 3100
rect 4240 3090 4280 3100
rect 4600 3090 4760 3100
rect 4880 3090 4920 3100
rect 6560 3090 6600 3100
rect 8400 3090 8440 3100
rect 9000 3090 9040 3100
rect 9240 3090 9360 3100
rect 9480 3090 9520 3100
rect 9800 3090 9880 3100
rect 2040 3080 2080 3090
rect 3160 3080 3200 3090
rect 4240 3080 4280 3090
rect 4600 3080 4760 3090
rect 4880 3080 4920 3090
rect 6560 3080 6600 3090
rect 8400 3080 8440 3090
rect 9000 3080 9040 3090
rect 9240 3080 9360 3090
rect 9480 3080 9520 3090
rect 9800 3080 9880 3090
rect 2040 3070 2080 3080
rect 3160 3070 3200 3080
rect 4240 3070 4280 3080
rect 4600 3070 4760 3080
rect 4880 3070 4920 3080
rect 6560 3070 6600 3080
rect 8400 3070 8440 3080
rect 9000 3070 9040 3080
rect 9240 3070 9360 3080
rect 9480 3070 9520 3080
rect 9800 3070 9880 3080
rect 2040 3060 2080 3070
rect 3160 3060 3200 3070
rect 4240 3060 4280 3070
rect 4600 3060 4760 3070
rect 4880 3060 4920 3070
rect 6560 3060 6600 3070
rect 8400 3060 8440 3070
rect 9000 3060 9040 3070
rect 9240 3060 9360 3070
rect 9480 3060 9520 3070
rect 9800 3060 9880 3070
rect 2000 3050 2040 3060
rect 3760 3050 3880 3060
rect 4160 3050 4200 3060
rect 4280 3050 4320 3060
rect 4520 3050 4560 3060
rect 4840 3050 4880 3060
rect 5200 3050 5240 3060
rect 6560 3050 6600 3060
rect 8920 3050 9040 3060
rect 9800 3050 9880 3060
rect 2000 3040 2040 3050
rect 3760 3040 3880 3050
rect 4160 3040 4200 3050
rect 4280 3040 4320 3050
rect 4520 3040 4560 3050
rect 4840 3040 4880 3050
rect 5200 3040 5240 3050
rect 6560 3040 6600 3050
rect 8920 3040 9040 3050
rect 9800 3040 9880 3050
rect 2000 3030 2040 3040
rect 3760 3030 3880 3040
rect 4160 3030 4200 3040
rect 4280 3030 4320 3040
rect 4520 3030 4560 3040
rect 4840 3030 4880 3040
rect 5200 3030 5240 3040
rect 6560 3030 6600 3040
rect 8920 3030 9040 3040
rect 9800 3030 9880 3040
rect 2000 3020 2040 3030
rect 3760 3020 3880 3030
rect 4160 3020 4200 3030
rect 4280 3020 4320 3030
rect 4520 3020 4560 3030
rect 4840 3020 4880 3030
rect 5200 3020 5240 3030
rect 6560 3020 6600 3030
rect 8920 3020 9040 3030
rect 9800 3020 9880 3030
rect 2000 3010 2040 3020
rect 4320 3010 4360 3020
rect 4480 3010 4680 3020
rect 4760 3010 4880 3020
rect 6560 3010 6600 3020
rect 8720 3010 8760 3020
rect 8920 3010 9040 3020
rect 9400 3010 9480 3020
rect 9800 3010 9880 3020
rect 2000 3000 2040 3010
rect 4320 3000 4360 3010
rect 4480 3000 4680 3010
rect 4760 3000 4880 3010
rect 6560 3000 6600 3010
rect 8720 3000 8760 3010
rect 8920 3000 9040 3010
rect 9400 3000 9480 3010
rect 9800 3000 9880 3010
rect 2000 2990 2040 3000
rect 4320 2990 4360 3000
rect 4480 2990 4680 3000
rect 4760 2990 4880 3000
rect 6560 2990 6600 3000
rect 8720 2990 8760 3000
rect 8920 2990 9040 3000
rect 9400 2990 9480 3000
rect 9800 2990 9880 3000
rect 2000 2980 2040 2990
rect 4320 2980 4360 2990
rect 4480 2980 4680 2990
rect 4760 2980 4880 2990
rect 6560 2980 6600 2990
rect 8720 2980 8760 2990
rect 8920 2980 9040 2990
rect 9400 2980 9480 2990
rect 9800 2980 9880 2990
rect 2000 2970 2040 2980
rect 4000 2970 4040 2980
rect 4160 2970 4200 2980
rect 4360 2970 4400 2980
rect 4480 2970 4920 2980
rect 5160 2970 5200 2980
rect 8280 2970 8320 2980
rect 8800 2970 8840 2980
rect 8920 2970 8960 2980
rect 9120 2970 9200 2980
rect 9280 2970 9440 2980
rect 2000 2960 2040 2970
rect 4000 2960 4040 2970
rect 4160 2960 4200 2970
rect 4360 2960 4400 2970
rect 4480 2960 4920 2970
rect 5160 2960 5200 2970
rect 8280 2960 8320 2970
rect 8800 2960 8840 2970
rect 8920 2960 8960 2970
rect 9120 2960 9200 2970
rect 9280 2960 9440 2970
rect 2000 2950 2040 2960
rect 4000 2950 4040 2960
rect 4160 2950 4200 2960
rect 4360 2950 4400 2960
rect 4480 2950 4920 2960
rect 5160 2950 5200 2960
rect 8280 2950 8320 2960
rect 8800 2950 8840 2960
rect 8920 2950 8960 2960
rect 9120 2950 9200 2960
rect 9280 2950 9440 2960
rect 2000 2940 2040 2950
rect 4000 2940 4040 2950
rect 4160 2940 4200 2950
rect 4360 2940 4400 2950
rect 4480 2940 4920 2950
rect 5160 2940 5200 2950
rect 8280 2940 8320 2950
rect 8800 2940 8840 2950
rect 8920 2940 8960 2950
rect 9120 2940 9200 2950
rect 9280 2940 9440 2950
rect 2000 2930 2040 2940
rect 3120 2930 3160 2940
rect 3880 2930 3960 2940
rect 4000 2930 4040 2940
rect 4200 2930 4240 2940
rect 4400 2930 4440 2940
rect 4520 2930 4920 2940
rect 8680 2930 8960 2940
rect 9120 2930 9200 2940
rect 9240 2930 9360 2940
rect 2000 2920 2040 2930
rect 3120 2920 3160 2930
rect 3880 2920 3960 2930
rect 4000 2920 4040 2930
rect 4200 2920 4240 2930
rect 4400 2920 4440 2930
rect 4520 2920 4920 2930
rect 8680 2920 8960 2930
rect 9120 2920 9200 2930
rect 9240 2920 9360 2930
rect 2000 2910 2040 2920
rect 3120 2910 3160 2920
rect 3880 2910 3960 2920
rect 4000 2910 4040 2920
rect 4200 2910 4240 2920
rect 4400 2910 4440 2920
rect 4520 2910 4920 2920
rect 8680 2910 8960 2920
rect 9120 2910 9200 2920
rect 9240 2910 9360 2920
rect 2000 2900 2040 2910
rect 3120 2900 3160 2910
rect 3880 2900 3960 2910
rect 4000 2900 4040 2910
rect 4200 2900 4240 2910
rect 4400 2900 4440 2910
rect 4520 2900 4920 2910
rect 8680 2900 8960 2910
rect 9120 2900 9200 2910
rect 9240 2900 9360 2910
rect 3120 2890 3160 2900
rect 4440 2890 5160 2900
rect 7400 2890 7480 2900
rect 8640 2890 8720 2900
rect 8800 2890 9000 2900
rect 9080 2890 9120 2900
rect 9200 2890 9360 2900
rect 3120 2880 3160 2890
rect 4440 2880 5160 2890
rect 7400 2880 7480 2890
rect 8640 2880 8720 2890
rect 8800 2880 9000 2890
rect 9080 2880 9120 2890
rect 9200 2880 9360 2890
rect 3120 2870 3160 2880
rect 4440 2870 5160 2880
rect 7400 2870 7480 2880
rect 8640 2870 8720 2880
rect 8800 2870 9000 2880
rect 9080 2870 9120 2880
rect 9200 2870 9360 2880
rect 3120 2860 3160 2870
rect 4440 2860 5160 2870
rect 7400 2860 7480 2870
rect 8640 2860 8720 2870
rect 8800 2860 9000 2870
rect 9080 2860 9120 2870
rect 9200 2860 9360 2870
rect 3960 2850 4000 2860
rect 4240 2850 4280 2860
rect 4520 2850 4640 2860
rect 4680 2850 5120 2860
rect 7200 2850 7240 2860
rect 7520 2850 7560 2860
rect 8200 2850 8240 2860
rect 8640 2850 8840 2860
rect 8880 2850 8960 2860
rect 9040 2850 9080 2860
rect 9200 2850 9360 2860
rect 3960 2840 4000 2850
rect 4240 2840 4280 2850
rect 4520 2840 4640 2850
rect 4680 2840 5120 2850
rect 7200 2840 7240 2850
rect 7520 2840 7560 2850
rect 8200 2840 8240 2850
rect 8640 2840 8840 2850
rect 8880 2840 8960 2850
rect 9040 2840 9080 2850
rect 9200 2840 9360 2850
rect 3960 2830 4000 2840
rect 4240 2830 4280 2840
rect 4520 2830 4640 2840
rect 4680 2830 5120 2840
rect 7200 2830 7240 2840
rect 7520 2830 7560 2840
rect 8200 2830 8240 2840
rect 8640 2830 8840 2840
rect 8880 2830 8960 2840
rect 9040 2830 9080 2840
rect 9200 2830 9360 2840
rect 3960 2820 4000 2830
rect 4240 2820 4280 2830
rect 4520 2820 4640 2830
rect 4680 2820 5120 2830
rect 7200 2820 7240 2830
rect 7520 2820 7560 2830
rect 8200 2820 8240 2830
rect 8640 2820 8840 2830
rect 8880 2820 8960 2830
rect 9040 2820 9080 2830
rect 9200 2820 9360 2830
rect 3120 2810 3160 2820
rect 4760 2810 5080 2820
rect 7560 2810 7600 2820
rect 8640 2810 8720 2820
rect 8800 2810 8880 2820
rect 9000 2810 9040 2820
rect 9160 2810 9200 2820
rect 9280 2810 9320 2820
rect 9400 2810 9440 2820
rect 3120 2800 3160 2810
rect 4760 2800 5080 2810
rect 7560 2800 7600 2810
rect 8640 2800 8720 2810
rect 8800 2800 8880 2810
rect 9000 2800 9040 2810
rect 9160 2800 9200 2810
rect 9280 2800 9320 2810
rect 9400 2800 9440 2810
rect 3120 2790 3160 2800
rect 4760 2790 5080 2800
rect 7560 2790 7600 2800
rect 8640 2790 8720 2800
rect 8800 2790 8880 2800
rect 9000 2790 9040 2800
rect 9160 2790 9200 2800
rect 9280 2790 9320 2800
rect 9400 2790 9440 2800
rect 3120 2780 3160 2790
rect 4760 2780 5080 2790
rect 7560 2780 7600 2790
rect 8640 2780 8720 2790
rect 8800 2780 8880 2790
rect 9000 2780 9040 2790
rect 9160 2780 9200 2790
rect 9280 2780 9320 2790
rect 9400 2780 9440 2790
rect 2000 2770 2040 2780
rect 3120 2770 3160 2780
rect 4840 2770 4920 2780
rect 5040 2770 5120 2780
rect 6040 2770 6120 2780
rect 8640 2770 8720 2780
rect 8920 2770 9200 2780
rect 9280 2770 9320 2780
rect 9480 2770 9520 2780
rect 9640 2770 9680 2780
rect 9920 2770 9990 2780
rect 2000 2760 2040 2770
rect 3120 2760 3160 2770
rect 4840 2760 4920 2770
rect 5040 2760 5120 2770
rect 6040 2760 6120 2770
rect 8640 2760 8720 2770
rect 8920 2760 9200 2770
rect 9280 2760 9320 2770
rect 9480 2760 9520 2770
rect 9640 2760 9680 2770
rect 9920 2760 9990 2770
rect 2000 2750 2040 2760
rect 3120 2750 3160 2760
rect 4840 2750 4920 2760
rect 5040 2750 5120 2760
rect 6040 2750 6120 2760
rect 8640 2750 8720 2760
rect 8920 2750 9200 2760
rect 9280 2750 9320 2760
rect 9480 2750 9520 2760
rect 9640 2750 9680 2760
rect 9920 2750 9990 2760
rect 2000 2740 2040 2750
rect 3120 2740 3160 2750
rect 4840 2740 4920 2750
rect 5040 2740 5120 2750
rect 6040 2740 6120 2750
rect 8640 2740 8720 2750
rect 8920 2740 9200 2750
rect 9280 2740 9320 2750
rect 9480 2740 9520 2750
rect 9640 2740 9680 2750
rect 9920 2740 9990 2750
rect 2000 2730 2040 2740
rect 5000 2730 5120 2740
rect 5960 2730 6160 2740
rect 7640 2730 7680 2740
rect 8640 2730 8680 2740
rect 8840 2730 8880 2740
rect 8920 2730 9280 2740
rect 9640 2730 9680 2740
rect 9920 2730 9960 2740
rect 2000 2720 2040 2730
rect 5000 2720 5120 2730
rect 5960 2720 6160 2730
rect 7640 2720 7680 2730
rect 8640 2720 8680 2730
rect 8840 2720 8880 2730
rect 8920 2720 9280 2730
rect 9640 2720 9680 2730
rect 9920 2720 9960 2730
rect 2000 2710 2040 2720
rect 5000 2710 5120 2720
rect 5960 2710 6160 2720
rect 7640 2710 7680 2720
rect 8640 2710 8680 2720
rect 8840 2710 8880 2720
rect 8920 2710 9280 2720
rect 9640 2710 9680 2720
rect 9920 2710 9960 2720
rect 2000 2700 2040 2710
rect 5000 2700 5120 2710
rect 5960 2700 6160 2710
rect 7640 2700 7680 2710
rect 8640 2700 8680 2710
rect 8840 2700 8880 2710
rect 8920 2700 9280 2710
rect 9640 2700 9680 2710
rect 9920 2700 9960 2710
rect 2280 2690 2320 2700
rect 2800 2690 2840 2700
rect 2920 2690 2960 2700
rect 3120 2690 3160 2700
rect 3880 2690 3920 2700
rect 5000 2690 5120 2700
rect 5880 2690 6200 2700
rect 6920 2690 6960 2700
rect 8640 2690 9000 2700
rect 9080 2690 9160 2700
rect 9640 2690 9680 2700
rect 9960 2690 9990 2700
rect 2280 2680 2320 2690
rect 2800 2680 2840 2690
rect 2920 2680 2960 2690
rect 3120 2680 3160 2690
rect 3880 2680 3920 2690
rect 5000 2680 5120 2690
rect 5880 2680 6200 2690
rect 6920 2680 6960 2690
rect 8640 2680 9000 2690
rect 9080 2680 9160 2690
rect 9640 2680 9680 2690
rect 9960 2680 9990 2690
rect 2280 2670 2320 2680
rect 2800 2670 2840 2680
rect 2920 2670 2960 2680
rect 3120 2670 3160 2680
rect 3880 2670 3920 2680
rect 5000 2670 5120 2680
rect 5880 2670 6200 2680
rect 6920 2670 6960 2680
rect 8640 2670 9000 2680
rect 9080 2670 9160 2680
rect 9640 2670 9680 2680
rect 9960 2670 9990 2680
rect 2280 2660 2320 2670
rect 2800 2660 2840 2670
rect 2920 2660 2960 2670
rect 3120 2660 3160 2670
rect 3880 2660 3920 2670
rect 5000 2660 5120 2670
rect 5880 2660 6200 2670
rect 6920 2660 6960 2670
rect 8640 2660 9000 2670
rect 9080 2660 9160 2670
rect 9640 2660 9680 2670
rect 9960 2660 9990 2670
rect 1960 2650 2000 2660
rect 2120 2650 2280 2660
rect 2400 2650 2440 2660
rect 2760 2650 2880 2660
rect 2920 2650 2960 2660
rect 3040 2650 3080 2660
rect 3880 2650 3920 2660
rect 4200 2650 4240 2660
rect 4960 2650 5080 2660
rect 5840 2650 6200 2660
rect 6880 2650 6920 2660
rect 8880 2650 9040 2660
rect 9720 2650 9760 2660
rect 9960 2650 9990 2660
rect 1960 2640 2000 2650
rect 2120 2640 2280 2650
rect 2400 2640 2440 2650
rect 2760 2640 2880 2650
rect 2920 2640 2960 2650
rect 3040 2640 3080 2650
rect 3880 2640 3920 2650
rect 4200 2640 4240 2650
rect 4960 2640 5080 2650
rect 5840 2640 6200 2650
rect 6880 2640 6920 2650
rect 8880 2640 9040 2650
rect 9720 2640 9760 2650
rect 9960 2640 9990 2650
rect 1960 2630 2000 2640
rect 2120 2630 2280 2640
rect 2400 2630 2440 2640
rect 2760 2630 2880 2640
rect 2920 2630 2960 2640
rect 3040 2630 3080 2640
rect 3880 2630 3920 2640
rect 4200 2630 4240 2640
rect 4960 2630 5080 2640
rect 5840 2630 6200 2640
rect 6880 2630 6920 2640
rect 8880 2630 9040 2640
rect 9720 2630 9760 2640
rect 9960 2630 9990 2640
rect 1960 2620 2000 2630
rect 2120 2620 2280 2630
rect 2400 2620 2440 2630
rect 2760 2620 2880 2630
rect 2920 2620 2960 2630
rect 3040 2620 3080 2630
rect 3880 2620 3920 2630
rect 4200 2620 4240 2630
rect 4960 2620 5080 2630
rect 5840 2620 6200 2630
rect 6880 2620 6920 2630
rect 8880 2620 9040 2630
rect 9720 2620 9760 2630
rect 9960 2620 9990 2630
rect 2040 2610 2080 2620
rect 2400 2610 2440 2620
rect 2760 2610 2840 2620
rect 4200 2610 4240 2620
rect 5800 2610 6240 2620
rect 6840 2610 6880 2620
rect 7720 2610 7760 2620
rect 8880 2610 9040 2620
rect 9160 2610 9200 2620
rect 9800 2610 9920 2620
rect 2040 2600 2080 2610
rect 2400 2600 2440 2610
rect 2760 2600 2840 2610
rect 4200 2600 4240 2610
rect 5800 2600 6240 2610
rect 6840 2600 6880 2610
rect 7720 2600 7760 2610
rect 8880 2600 9040 2610
rect 9160 2600 9200 2610
rect 9800 2600 9920 2610
rect 2040 2590 2080 2600
rect 2400 2590 2440 2600
rect 2760 2590 2840 2600
rect 4200 2590 4240 2600
rect 5800 2590 6240 2600
rect 6840 2590 6880 2600
rect 7720 2590 7760 2600
rect 8880 2590 9040 2600
rect 9160 2590 9200 2600
rect 9800 2590 9920 2600
rect 2040 2580 2080 2590
rect 2400 2580 2440 2590
rect 2760 2580 2840 2590
rect 4200 2580 4240 2590
rect 5800 2580 6240 2590
rect 6840 2580 6880 2590
rect 7720 2580 7760 2590
rect 8880 2580 9040 2590
rect 9160 2580 9200 2590
rect 9800 2580 9920 2590
rect 1920 2570 1960 2580
rect 2000 2570 2040 2580
rect 3920 2570 3960 2580
rect 4160 2570 4240 2580
rect 5760 2570 6280 2580
rect 6800 2570 6840 2580
rect 7240 2570 7280 2580
rect 7760 2570 7800 2580
rect 8880 2570 8920 2580
rect 9000 2570 9040 2580
rect 9880 2570 9990 2580
rect 1920 2560 1960 2570
rect 2000 2560 2040 2570
rect 3920 2560 3960 2570
rect 4160 2560 4240 2570
rect 5760 2560 6280 2570
rect 6800 2560 6840 2570
rect 7240 2560 7280 2570
rect 7760 2560 7800 2570
rect 8880 2560 8920 2570
rect 9000 2560 9040 2570
rect 9880 2560 9990 2570
rect 1920 2550 1960 2560
rect 2000 2550 2040 2560
rect 3920 2550 3960 2560
rect 4160 2550 4240 2560
rect 5760 2550 6280 2560
rect 6800 2550 6840 2560
rect 7240 2550 7280 2560
rect 7760 2550 7800 2560
rect 8880 2550 8920 2560
rect 9000 2550 9040 2560
rect 9880 2550 9990 2560
rect 1920 2540 1960 2550
rect 2000 2540 2040 2550
rect 3920 2540 3960 2550
rect 4160 2540 4240 2550
rect 5760 2540 6280 2550
rect 6800 2540 6840 2550
rect 7240 2540 7280 2550
rect 7760 2540 7800 2550
rect 8880 2540 8920 2550
rect 9000 2540 9040 2550
rect 9880 2540 9990 2550
rect 1920 2530 2120 2540
rect 2160 2530 2360 2540
rect 3160 2530 3200 2540
rect 3960 2530 4000 2540
rect 4080 2530 4160 2540
rect 5760 2530 6280 2540
rect 7240 2530 7320 2540
rect 7880 2530 7920 2540
rect 9000 2530 9080 2540
rect 9120 2530 9160 2540
rect 9360 2530 9600 2540
rect 9960 2530 9990 2540
rect 1920 2520 2120 2530
rect 2160 2520 2360 2530
rect 3160 2520 3200 2530
rect 3960 2520 4000 2530
rect 4080 2520 4160 2530
rect 5760 2520 6280 2530
rect 7240 2520 7320 2530
rect 7880 2520 7920 2530
rect 9000 2520 9080 2530
rect 9120 2520 9160 2530
rect 9360 2520 9600 2530
rect 9960 2520 9990 2530
rect 1920 2510 2120 2520
rect 2160 2510 2360 2520
rect 3160 2510 3200 2520
rect 3960 2510 4000 2520
rect 4080 2510 4160 2520
rect 5760 2510 6280 2520
rect 7240 2510 7320 2520
rect 7880 2510 7920 2520
rect 9000 2510 9080 2520
rect 9120 2510 9160 2520
rect 9360 2510 9600 2520
rect 9960 2510 9990 2520
rect 1920 2500 2120 2510
rect 2160 2500 2360 2510
rect 3160 2500 3200 2510
rect 3960 2500 4000 2510
rect 4080 2500 4160 2510
rect 5760 2500 6280 2510
rect 7240 2500 7320 2510
rect 7880 2500 7920 2510
rect 9000 2500 9080 2510
rect 9120 2500 9160 2510
rect 9360 2500 9600 2510
rect 9960 2500 9990 2510
rect 1920 2490 1960 2500
rect 3200 2490 3240 2500
rect 5600 2490 5640 2500
rect 5760 2490 6320 2500
rect 7320 2490 7360 2500
rect 8960 2490 9120 2500
rect 9280 2490 9320 2500
rect 9600 2490 9680 2500
rect 1920 2480 1960 2490
rect 3200 2480 3240 2490
rect 5600 2480 5640 2490
rect 5760 2480 6320 2490
rect 7320 2480 7360 2490
rect 8960 2480 9120 2490
rect 9280 2480 9320 2490
rect 9600 2480 9680 2490
rect 1920 2470 1960 2480
rect 3200 2470 3240 2480
rect 5600 2470 5640 2480
rect 5760 2470 6320 2480
rect 7320 2470 7360 2480
rect 8960 2470 9120 2480
rect 9280 2470 9320 2480
rect 9600 2470 9680 2480
rect 1920 2460 1960 2470
rect 3200 2460 3240 2470
rect 5600 2460 5640 2470
rect 5760 2460 6320 2470
rect 7320 2460 7360 2470
rect 8960 2460 9120 2470
rect 9280 2460 9320 2470
rect 9600 2460 9680 2470
rect 5560 2450 5640 2460
rect 5720 2450 6360 2460
rect 6760 2450 6800 2460
rect 7360 2450 7400 2460
rect 9280 2450 9400 2460
rect 9480 2450 9560 2460
rect 9640 2450 9760 2460
rect 5560 2440 5640 2450
rect 5720 2440 6360 2450
rect 6760 2440 6800 2450
rect 7360 2440 7400 2450
rect 9280 2440 9400 2450
rect 9480 2440 9560 2450
rect 9640 2440 9760 2450
rect 5560 2430 5640 2440
rect 5720 2430 6360 2440
rect 6760 2430 6800 2440
rect 7360 2430 7400 2440
rect 9280 2430 9400 2440
rect 9480 2430 9560 2440
rect 9640 2430 9760 2440
rect 5560 2420 5640 2430
rect 5720 2420 6360 2430
rect 6760 2420 6800 2430
rect 7360 2420 7400 2430
rect 9280 2420 9400 2430
rect 9480 2420 9560 2430
rect 9640 2420 9760 2430
rect 1880 2410 1920 2420
rect 3240 2410 3280 2420
rect 5560 2410 5600 2420
rect 5680 2410 6360 2420
rect 6760 2410 6880 2420
rect 7360 2410 7440 2420
rect 9280 2410 9480 2420
rect 9560 2410 9800 2420
rect 1880 2400 1920 2410
rect 3240 2400 3280 2410
rect 5560 2400 5600 2410
rect 5680 2400 6360 2410
rect 6760 2400 6880 2410
rect 7360 2400 7440 2410
rect 9280 2400 9480 2410
rect 9560 2400 9800 2410
rect 1880 2390 1920 2400
rect 3240 2390 3280 2400
rect 5560 2390 5600 2400
rect 5680 2390 6360 2400
rect 6760 2390 6880 2400
rect 7360 2390 7440 2400
rect 9280 2390 9480 2400
rect 9560 2390 9800 2400
rect 1880 2380 1920 2390
rect 3240 2380 3280 2390
rect 5560 2380 5600 2390
rect 5680 2380 6360 2390
rect 6760 2380 6880 2390
rect 7360 2380 7440 2390
rect 9280 2380 9480 2390
rect 9560 2380 9800 2390
rect 1880 2370 1920 2380
rect 3240 2370 3280 2380
rect 5680 2370 6400 2380
rect 6720 2370 6920 2380
rect 7440 2370 7480 2380
rect 8400 2370 8440 2380
rect 9280 2370 9480 2380
rect 9560 2370 9680 2380
rect 9760 2370 9800 2380
rect 1880 2360 1920 2370
rect 3240 2360 3280 2370
rect 5680 2360 6400 2370
rect 6720 2360 6920 2370
rect 7440 2360 7480 2370
rect 8400 2360 8440 2370
rect 9280 2360 9480 2370
rect 9560 2360 9680 2370
rect 9760 2360 9800 2370
rect 1880 2350 1920 2360
rect 3240 2350 3280 2360
rect 5680 2350 6400 2360
rect 6720 2350 6920 2360
rect 7440 2350 7480 2360
rect 8400 2350 8440 2360
rect 9280 2350 9480 2360
rect 9560 2350 9680 2360
rect 9760 2350 9800 2360
rect 1880 2340 1920 2350
rect 3240 2340 3280 2350
rect 5680 2340 6400 2350
rect 6720 2340 6920 2350
rect 7440 2340 7480 2350
rect 8400 2340 8440 2350
rect 9280 2340 9480 2350
rect 9560 2340 9680 2350
rect 9760 2340 9800 2350
rect 5640 2330 6400 2340
rect 6720 2330 6840 2340
rect 6920 2330 7040 2340
rect 7480 2330 7520 2340
rect 8520 2330 8560 2340
rect 9200 2330 9240 2340
rect 9280 2330 9320 2340
rect 9400 2330 9480 2340
rect 9560 2330 9600 2340
rect 9760 2330 9800 2340
rect 5640 2320 6400 2330
rect 6720 2320 6840 2330
rect 6920 2320 7040 2330
rect 7480 2320 7520 2330
rect 8520 2320 8560 2330
rect 9200 2320 9240 2330
rect 9280 2320 9320 2330
rect 9400 2320 9480 2330
rect 9560 2320 9600 2330
rect 9760 2320 9800 2330
rect 5640 2310 6400 2320
rect 6720 2310 6840 2320
rect 6920 2310 7040 2320
rect 7480 2310 7520 2320
rect 8520 2310 8560 2320
rect 9200 2310 9240 2320
rect 9280 2310 9320 2320
rect 9400 2310 9480 2320
rect 9560 2310 9600 2320
rect 9760 2310 9800 2320
rect 5640 2300 6400 2310
rect 6720 2300 6840 2310
rect 6920 2300 7040 2310
rect 7480 2300 7520 2310
rect 8520 2300 8560 2310
rect 9200 2300 9240 2310
rect 9280 2300 9320 2310
rect 9400 2300 9480 2310
rect 9560 2300 9600 2310
rect 9760 2300 9800 2310
rect 3280 2290 3320 2300
rect 5440 2290 5520 2300
rect 5640 2290 6440 2300
rect 6720 2290 6840 2300
rect 6960 2290 7080 2300
rect 7120 2290 7240 2300
rect 7560 2290 7600 2300
rect 8560 2290 8600 2300
rect 9120 2290 9160 2300
rect 9480 2290 9600 2300
rect 9760 2290 9800 2300
rect 3280 2280 3320 2290
rect 5440 2280 5520 2290
rect 5640 2280 6440 2290
rect 6720 2280 6840 2290
rect 6960 2280 7080 2290
rect 7120 2280 7240 2290
rect 7560 2280 7600 2290
rect 8560 2280 8600 2290
rect 9120 2280 9160 2290
rect 9480 2280 9600 2290
rect 9760 2280 9800 2290
rect 3280 2270 3320 2280
rect 5440 2270 5520 2280
rect 5640 2270 6440 2280
rect 6720 2270 6840 2280
rect 6960 2270 7080 2280
rect 7120 2270 7240 2280
rect 7560 2270 7600 2280
rect 8560 2270 8600 2280
rect 9120 2270 9160 2280
rect 9480 2270 9600 2280
rect 9760 2270 9800 2280
rect 3280 2260 3320 2270
rect 5440 2260 5520 2270
rect 5640 2260 6440 2270
rect 6720 2260 6840 2270
rect 6960 2260 7080 2270
rect 7120 2260 7240 2270
rect 7560 2260 7600 2270
rect 8560 2260 8600 2270
rect 9120 2260 9160 2270
rect 9480 2260 9600 2270
rect 9760 2260 9800 2270
rect 1840 2250 1880 2260
rect 3280 2250 3320 2260
rect 5400 2250 5520 2260
rect 5600 2250 6400 2260
rect 6440 2250 6480 2260
rect 6800 2250 6840 2260
rect 7280 2250 7400 2260
rect 7600 2250 7640 2260
rect 8640 2250 8680 2260
rect 8720 2250 8800 2260
rect 9080 2250 9120 2260
rect 9320 2250 9360 2260
rect 9760 2250 9800 2260
rect 1840 2240 1880 2250
rect 3280 2240 3320 2250
rect 5400 2240 5520 2250
rect 5600 2240 6400 2250
rect 6440 2240 6480 2250
rect 6800 2240 6840 2250
rect 7280 2240 7400 2250
rect 7600 2240 7640 2250
rect 8640 2240 8680 2250
rect 8720 2240 8800 2250
rect 9080 2240 9120 2250
rect 9320 2240 9360 2250
rect 9760 2240 9800 2250
rect 1840 2230 1880 2240
rect 3280 2230 3320 2240
rect 5400 2230 5520 2240
rect 5600 2230 6400 2240
rect 6440 2230 6480 2240
rect 6800 2230 6840 2240
rect 7280 2230 7400 2240
rect 7600 2230 7640 2240
rect 8640 2230 8680 2240
rect 8720 2230 8800 2240
rect 9080 2230 9120 2240
rect 9320 2230 9360 2240
rect 9760 2230 9800 2240
rect 1840 2220 1880 2230
rect 3280 2220 3320 2230
rect 5400 2220 5520 2230
rect 5600 2220 6400 2230
rect 6440 2220 6480 2230
rect 6800 2220 6840 2230
rect 7280 2220 7400 2230
rect 7600 2220 7640 2230
rect 8640 2220 8680 2230
rect 8720 2220 8800 2230
rect 9080 2220 9120 2230
rect 9320 2220 9360 2230
rect 9760 2220 9800 2230
rect 1840 2210 1880 2220
rect 2600 2210 2720 2220
rect 3280 2210 3320 2220
rect 5360 2210 6400 2220
rect 6440 2210 6480 2220
rect 6800 2210 6920 2220
rect 7360 2210 7400 2220
rect 7640 2210 7680 2220
rect 8840 2210 9000 2220
rect 9400 2210 9480 2220
rect 9760 2210 9800 2220
rect 1840 2200 1880 2210
rect 2600 2200 2720 2210
rect 3280 2200 3320 2210
rect 5360 2200 6400 2210
rect 6440 2200 6480 2210
rect 6800 2200 6920 2210
rect 7360 2200 7400 2210
rect 7640 2200 7680 2210
rect 8840 2200 9000 2210
rect 9400 2200 9480 2210
rect 9760 2200 9800 2210
rect 1840 2190 1880 2200
rect 2600 2190 2720 2200
rect 3280 2190 3320 2200
rect 5360 2190 6400 2200
rect 6440 2190 6480 2200
rect 6800 2190 6920 2200
rect 7360 2190 7400 2200
rect 7640 2190 7680 2200
rect 8840 2190 9000 2200
rect 9400 2190 9480 2200
rect 9760 2190 9800 2200
rect 1840 2180 1880 2190
rect 2600 2180 2720 2190
rect 3280 2180 3320 2190
rect 5360 2180 6400 2190
rect 6440 2180 6480 2190
rect 6800 2180 6920 2190
rect 7360 2180 7400 2190
rect 7640 2180 7680 2190
rect 8840 2180 9000 2190
rect 9400 2180 9480 2190
rect 9760 2180 9800 2190
rect 1840 2170 1880 2180
rect 2400 2170 2440 2180
rect 2520 2170 2640 2180
rect 2720 2170 2800 2180
rect 3280 2170 3320 2180
rect 5320 2170 6400 2180
rect 6840 2170 6960 2180
rect 7400 2170 7480 2180
rect 7720 2170 7760 2180
rect 8360 2170 8400 2180
rect 9480 2170 9600 2180
rect 9680 2170 9760 2180
rect 1840 2160 1880 2170
rect 2400 2160 2440 2170
rect 2520 2160 2640 2170
rect 2720 2160 2800 2170
rect 3280 2160 3320 2170
rect 5320 2160 6400 2170
rect 6840 2160 6960 2170
rect 7400 2160 7480 2170
rect 7720 2160 7760 2170
rect 8360 2160 8400 2170
rect 9480 2160 9600 2170
rect 9680 2160 9760 2170
rect 1840 2150 1880 2160
rect 2400 2150 2440 2160
rect 2520 2150 2640 2160
rect 2720 2150 2800 2160
rect 3280 2150 3320 2160
rect 5320 2150 6400 2160
rect 6840 2150 6960 2160
rect 7400 2150 7480 2160
rect 7720 2150 7760 2160
rect 8360 2150 8400 2160
rect 9480 2150 9600 2160
rect 9680 2150 9760 2160
rect 1840 2140 1880 2150
rect 2400 2140 2440 2150
rect 2520 2140 2640 2150
rect 2720 2140 2800 2150
rect 3280 2140 3320 2150
rect 5320 2140 6400 2150
rect 6840 2140 6960 2150
rect 7400 2140 7480 2150
rect 7720 2140 7760 2150
rect 8360 2140 8400 2150
rect 9480 2140 9600 2150
rect 9680 2140 9760 2150
rect 1840 2130 1880 2140
rect 2560 2130 2640 2140
rect 3280 2130 3320 2140
rect 5280 2130 6360 2140
rect 6480 2130 6520 2140
rect 6760 2130 6800 2140
rect 6880 2130 7000 2140
rect 7280 2130 7320 2140
rect 9240 2130 9320 2140
rect 9640 2130 9680 2140
rect 1840 2120 1880 2130
rect 2560 2120 2640 2130
rect 3280 2120 3320 2130
rect 5280 2120 6360 2130
rect 6480 2120 6520 2130
rect 6760 2120 6800 2130
rect 6880 2120 7000 2130
rect 7280 2120 7320 2130
rect 9240 2120 9320 2130
rect 9640 2120 9680 2130
rect 1840 2110 1880 2120
rect 2560 2110 2640 2120
rect 3280 2110 3320 2120
rect 5280 2110 6360 2120
rect 6480 2110 6520 2120
rect 6760 2110 6800 2120
rect 6880 2110 7000 2120
rect 7280 2110 7320 2120
rect 9240 2110 9320 2120
rect 9640 2110 9680 2120
rect 1840 2100 1880 2110
rect 2560 2100 2640 2110
rect 3280 2100 3320 2110
rect 5280 2100 6360 2110
rect 6480 2100 6520 2110
rect 6760 2100 6800 2110
rect 6880 2100 7000 2110
rect 7280 2100 7320 2110
rect 9240 2100 9320 2110
rect 9640 2100 9680 2110
rect 1840 2090 1880 2100
rect 3280 2090 3320 2100
rect 5280 2090 6400 2100
rect 6480 2090 6520 2100
rect 6760 2090 6800 2100
rect 6920 2090 7080 2100
rect 7240 2090 7280 2100
rect 8400 2090 8440 2100
rect 9200 2090 9240 2100
rect 9280 2090 9320 2100
rect 9480 2090 9520 2100
rect 1840 2080 1880 2090
rect 3280 2080 3320 2090
rect 5280 2080 6400 2090
rect 6480 2080 6520 2090
rect 6760 2080 6800 2090
rect 6920 2080 7080 2090
rect 7240 2080 7280 2090
rect 8400 2080 8440 2090
rect 9200 2080 9240 2090
rect 9280 2080 9320 2090
rect 9480 2080 9520 2090
rect 1840 2070 1880 2080
rect 3280 2070 3320 2080
rect 5280 2070 6400 2080
rect 6480 2070 6520 2080
rect 6760 2070 6800 2080
rect 6920 2070 7080 2080
rect 7240 2070 7280 2080
rect 8400 2070 8440 2080
rect 9200 2070 9240 2080
rect 9280 2070 9320 2080
rect 9480 2070 9520 2080
rect 1840 2060 1880 2070
rect 3280 2060 3320 2070
rect 5280 2060 6400 2070
rect 6480 2060 6520 2070
rect 6760 2060 6800 2070
rect 6920 2060 7080 2070
rect 7240 2060 7280 2070
rect 8400 2060 8440 2070
rect 9200 2060 9240 2070
rect 9280 2060 9320 2070
rect 9480 2060 9520 2070
rect 1840 2050 1880 2060
rect 3240 2050 3320 2060
rect 5120 2050 5160 2060
rect 5240 2050 6360 2060
rect 6480 2050 6520 2060
rect 6760 2050 6800 2060
rect 6960 2050 7280 2060
rect 7880 2050 8000 2060
rect 8400 2050 8520 2060
rect 9120 2050 9240 2060
rect 9320 2050 9360 2060
rect 1840 2040 1880 2050
rect 3240 2040 3320 2050
rect 5120 2040 5160 2050
rect 5240 2040 6360 2050
rect 6480 2040 6520 2050
rect 6760 2040 6800 2050
rect 6960 2040 7280 2050
rect 7880 2040 8000 2050
rect 8400 2040 8520 2050
rect 9120 2040 9240 2050
rect 9320 2040 9360 2050
rect 1840 2030 1880 2040
rect 3240 2030 3320 2040
rect 5120 2030 5160 2040
rect 5240 2030 6360 2040
rect 6480 2030 6520 2040
rect 6760 2030 6800 2040
rect 6960 2030 7280 2040
rect 7880 2030 8000 2040
rect 8400 2030 8520 2040
rect 9120 2030 9240 2040
rect 9320 2030 9360 2040
rect 1840 2020 1880 2030
rect 3240 2020 3320 2030
rect 5120 2020 5160 2030
rect 5240 2020 6360 2030
rect 6480 2020 6520 2030
rect 6760 2020 6800 2030
rect 6960 2020 7280 2030
rect 7880 2020 8000 2030
rect 8400 2020 8520 2030
rect 9120 2020 9240 2030
rect 9320 2020 9360 2030
rect 1840 2010 1880 2020
rect 3240 2010 3320 2020
rect 5120 2010 6360 2020
rect 6480 2010 6520 2020
rect 6800 2010 6840 2020
rect 7040 2010 7280 2020
rect 7320 2010 7360 2020
rect 8400 2010 8440 2020
rect 8520 2010 8600 2020
rect 9040 2010 9080 2020
rect 1840 2000 1880 2010
rect 3240 2000 3320 2010
rect 5120 2000 6360 2010
rect 6480 2000 6520 2010
rect 6800 2000 6840 2010
rect 7040 2000 7280 2010
rect 7320 2000 7360 2010
rect 8400 2000 8440 2010
rect 8520 2000 8600 2010
rect 9040 2000 9080 2010
rect 1840 1990 1880 2000
rect 3240 1990 3320 2000
rect 5120 1990 6360 2000
rect 6480 1990 6520 2000
rect 6800 1990 6840 2000
rect 7040 1990 7280 2000
rect 7320 1990 7360 2000
rect 8400 1990 8440 2000
rect 8520 1990 8600 2000
rect 9040 1990 9080 2000
rect 1840 1980 1880 1990
rect 3240 1980 3320 1990
rect 5120 1980 6360 1990
rect 6480 1980 6520 1990
rect 6800 1980 6840 1990
rect 7040 1980 7280 1990
rect 7320 1980 7360 1990
rect 8400 1980 8440 1990
rect 8520 1980 8600 1990
rect 9040 1980 9080 1990
rect 1840 1970 1880 1980
rect 3240 1970 3320 1980
rect 5040 1970 6200 1980
rect 6280 1970 6360 1980
rect 6480 1970 6520 1980
rect 6800 1970 6840 1980
rect 7120 1970 7240 1980
rect 7320 1970 7360 1980
rect 7760 1970 7880 1980
rect 8400 1970 8440 1980
rect 8640 1970 8760 1980
rect 8800 1970 9040 1980
rect 1840 1960 1880 1970
rect 3240 1960 3320 1970
rect 5040 1960 6200 1970
rect 6280 1960 6360 1970
rect 6480 1960 6520 1970
rect 6800 1960 6840 1970
rect 7120 1960 7240 1970
rect 7320 1960 7360 1970
rect 7760 1960 7880 1970
rect 8400 1960 8440 1970
rect 8640 1960 8760 1970
rect 8800 1960 9040 1970
rect 1840 1950 1880 1960
rect 3240 1950 3320 1960
rect 5040 1950 6200 1960
rect 6280 1950 6360 1960
rect 6480 1950 6520 1960
rect 6800 1950 6840 1960
rect 7120 1950 7240 1960
rect 7320 1950 7360 1960
rect 7760 1950 7880 1960
rect 8400 1950 8440 1960
rect 8640 1950 8760 1960
rect 8800 1950 9040 1960
rect 1840 1940 1880 1950
rect 3240 1940 3320 1950
rect 5040 1940 6200 1950
rect 6280 1940 6360 1950
rect 6480 1940 6520 1950
rect 6800 1940 6840 1950
rect 7120 1940 7240 1950
rect 7320 1940 7360 1950
rect 7760 1940 7880 1950
rect 8400 1940 8440 1950
rect 8640 1940 8760 1950
rect 8800 1940 9040 1950
rect 1840 1930 1880 1940
rect 3240 1930 3320 1940
rect 4520 1930 4640 1940
rect 4760 1930 4800 1940
rect 4840 1930 4880 1940
rect 4960 1930 6200 1940
rect 6320 1930 6400 1940
rect 6480 1930 6520 1940
rect 6800 1930 6840 1940
rect 7320 1930 7360 1940
rect 7760 1930 7840 1940
rect 8400 1930 8440 1940
rect 1840 1920 1880 1930
rect 3240 1920 3320 1930
rect 4520 1920 4640 1930
rect 4760 1920 4800 1930
rect 4840 1920 4880 1930
rect 4960 1920 6200 1930
rect 6320 1920 6400 1930
rect 6480 1920 6520 1930
rect 6800 1920 6840 1930
rect 7320 1920 7360 1930
rect 7760 1920 7840 1930
rect 8400 1920 8440 1930
rect 1840 1910 1880 1920
rect 3240 1910 3320 1920
rect 4520 1910 4640 1920
rect 4760 1910 4800 1920
rect 4840 1910 4880 1920
rect 4960 1910 6200 1920
rect 6320 1910 6400 1920
rect 6480 1910 6520 1920
rect 6800 1910 6840 1920
rect 7320 1910 7360 1920
rect 7760 1910 7840 1920
rect 8400 1910 8440 1920
rect 1840 1900 1880 1910
rect 3240 1900 3320 1910
rect 4520 1900 4640 1910
rect 4760 1900 4800 1910
rect 4840 1900 4880 1910
rect 4960 1900 6200 1910
rect 6320 1900 6400 1910
rect 6480 1900 6520 1910
rect 6800 1900 6840 1910
rect 7320 1900 7360 1910
rect 7760 1900 7840 1910
rect 8400 1900 8440 1910
rect 1840 1890 1880 1900
rect 2440 1890 2480 1900
rect 2720 1890 2800 1900
rect 3280 1890 3320 1900
rect 4400 1890 4440 1900
rect 4520 1890 4600 1900
rect 4640 1890 4680 1900
rect 4760 1890 4800 1900
rect 4840 1890 4920 1900
rect 4960 1890 5000 1900
rect 5040 1890 5080 1900
rect 5160 1890 6160 1900
rect 6360 1890 6480 1900
rect 6800 1890 6840 1900
rect 7320 1890 7360 1900
rect 7800 1890 7840 1900
rect 8400 1890 8440 1900
rect 1840 1880 1880 1890
rect 2440 1880 2480 1890
rect 2720 1880 2800 1890
rect 3280 1880 3320 1890
rect 4400 1880 4440 1890
rect 4520 1880 4600 1890
rect 4640 1880 4680 1890
rect 4760 1880 4800 1890
rect 4840 1880 4920 1890
rect 4960 1880 5000 1890
rect 5040 1880 5080 1890
rect 5160 1880 6160 1890
rect 6360 1880 6480 1890
rect 6800 1880 6840 1890
rect 7320 1880 7360 1890
rect 7800 1880 7840 1890
rect 8400 1880 8440 1890
rect 1840 1870 1880 1880
rect 2440 1870 2480 1880
rect 2720 1870 2800 1880
rect 3280 1870 3320 1880
rect 4400 1870 4440 1880
rect 4520 1870 4600 1880
rect 4640 1870 4680 1880
rect 4760 1870 4800 1880
rect 4840 1870 4920 1880
rect 4960 1870 5000 1880
rect 5040 1870 5080 1880
rect 5160 1870 6160 1880
rect 6360 1870 6480 1880
rect 6800 1870 6840 1880
rect 7320 1870 7360 1880
rect 7800 1870 7840 1880
rect 8400 1870 8440 1880
rect 1840 1860 1880 1870
rect 2440 1860 2480 1870
rect 2720 1860 2800 1870
rect 3280 1860 3320 1870
rect 4400 1860 4440 1870
rect 4520 1860 4600 1870
rect 4640 1860 4680 1870
rect 4760 1860 4800 1870
rect 4840 1860 4920 1870
rect 4960 1860 5000 1870
rect 5040 1860 5080 1870
rect 5160 1860 6160 1870
rect 6360 1860 6480 1870
rect 6800 1860 6840 1870
rect 7320 1860 7360 1870
rect 7800 1860 7840 1870
rect 8400 1860 8440 1870
rect 1840 1850 1880 1860
rect 2360 1850 2400 1860
rect 2840 1850 2880 1860
rect 3280 1850 3320 1860
rect 4520 1850 4600 1860
rect 4640 1850 4680 1860
rect 4720 1850 4800 1860
rect 4840 1850 5000 1860
rect 5040 1850 5160 1860
rect 5200 1850 5240 1860
rect 5320 1850 6120 1860
rect 6280 1850 6480 1860
rect 6800 1850 6840 1860
rect 7320 1850 7360 1860
rect 7800 1850 7840 1860
rect 8360 1850 8440 1860
rect 9120 1850 9200 1860
rect 9720 1850 9760 1860
rect 9960 1850 9990 1860
rect 1840 1840 1880 1850
rect 2360 1840 2400 1850
rect 2840 1840 2880 1850
rect 3280 1840 3320 1850
rect 4520 1840 4600 1850
rect 4640 1840 4680 1850
rect 4720 1840 4800 1850
rect 4840 1840 5000 1850
rect 5040 1840 5160 1850
rect 5200 1840 5240 1850
rect 5320 1840 6120 1850
rect 6280 1840 6480 1850
rect 6800 1840 6840 1850
rect 7320 1840 7360 1850
rect 7800 1840 7840 1850
rect 8360 1840 8440 1850
rect 9120 1840 9200 1850
rect 9720 1840 9760 1850
rect 9960 1840 9990 1850
rect 1840 1830 1880 1840
rect 2360 1830 2400 1840
rect 2840 1830 2880 1840
rect 3280 1830 3320 1840
rect 4520 1830 4600 1840
rect 4640 1830 4680 1840
rect 4720 1830 4800 1840
rect 4840 1830 5000 1840
rect 5040 1830 5160 1840
rect 5200 1830 5240 1840
rect 5320 1830 6120 1840
rect 6280 1830 6480 1840
rect 6800 1830 6840 1840
rect 7320 1830 7360 1840
rect 7800 1830 7840 1840
rect 8360 1830 8440 1840
rect 9120 1830 9200 1840
rect 9720 1830 9760 1840
rect 9960 1830 9990 1840
rect 1840 1820 1880 1830
rect 2360 1820 2400 1830
rect 2840 1820 2880 1830
rect 3280 1820 3320 1830
rect 4520 1820 4600 1830
rect 4640 1820 4680 1830
rect 4720 1820 4800 1830
rect 4840 1820 5000 1830
rect 5040 1820 5160 1830
rect 5200 1820 5240 1830
rect 5320 1820 6120 1830
rect 6280 1820 6480 1830
rect 6800 1820 6840 1830
rect 7320 1820 7360 1830
rect 7800 1820 7840 1830
rect 8360 1820 8440 1830
rect 9120 1820 9200 1830
rect 9720 1820 9760 1830
rect 9960 1820 9990 1830
rect 1840 1810 1880 1820
rect 2280 1810 2320 1820
rect 2760 1810 2800 1820
rect 3280 1810 3320 1820
rect 4080 1810 4120 1820
rect 4360 1810 4400 1820
rect 4560 1810 4640 1820
rect 4720 1810 4800 1820
rect 4880 1810 5000 1820
rect 5080 1810 5160 1820
rect 5200 1810 5320 1820
rect 5360 1810 6080 1820
rect 6280 1810 6360 1820
rect 6440 1810 6520 1820
rect 6800 1810 6840 1820
rect 7320 1810 7360 1820
rect 7800 1810 7840 1820
rect 8360 1810 8440 1820
rect 9720 1810 9760 1820
rect 1840 1800 1880 1810
rect 2280 1800 2320 1810
rect 2760 1800 2800 1810
rect 3280 1800 3320 1810
rect 4080 1800 4120 1810
rect 4360 1800 4400 1810
rect 4560 1800 4640 1810
rect 4720 1800 4800 1810
rect 4880 1800 5000 1810
rect 5080 1800 5160 1810
rect 5200 1800 5320 1810
rect 5360 1800 6080 1810
rect 6280 1800 6360 1810
rect 6440 1800 6520 1810
rect 6800 1800 6840 1810
rect 7320 1800 7360 1810
rect 7800 1800 7840 1810
rect 8360 1800 8440 1810
rect 9720 1800 9760 1810
rect 1840 1790 1880 1800
rect 2280 1790 2320 1800
rect 2760 1790 2800 1800
rect 3280 1790 3320 1800
rect 4080 1790 4120 1800
rect 4360 1790 4400 1800
rect 4560 1790 4640 1800
rect 4720 1790 4800 1800
rect 4880 1790 5000 1800
rect 5080 1790 5160 1800
rect 5200 1790 5320 1800
rect 5360 1790 6080 1800
rect 6280 1790 6360 1800
rect 6440 1790 6520 1800
rect 6800 1790 6840 1800
rect 7320 1790 7360 1800
rect 7800 1790 7840 1800
rect 8360 1790 8440 1800
rect 9720 1790 9760 1800
rect 1840 1780 1880 1790
rect 2280 1780 2320 1790
rect 2760 1780 2800 1790
rect 3280 1780 3320 1790
rect 4080 1780 4120 1790
rect 4360 1780 4400 1790
rect 4560 1780 4640 1790
rect 4720 1780 4800 1790
rect 4880 1780 5000 1790
rect 5080 1780 5160 1790
rect 5200 1780 5320 1790
rect 5360 1780 6080 1790
rect 6280 1780 6360 1790
rect 6440 1780 6520 1790
rect 6800 1780 6840 1790
rect 7320 1780 7360 1790
rect 7800 1780 7840 1790
rect 8360 1780 8440 1790
rect 9720 1780 9760 1790
rect 2440 1770 2520 1780
rect 3240 1770 3280 1780
rect 4360 1770 4400 1780
rect 4520 1770 4560 1780
rect 4600 1770 4640 1780
rect 4760 1770 4840 1780
rect 4880 1770 4960 1780
rect 5080 1770 5120 1780
rect 5160 1770 5200 1780
rect 5320 1770 5400 1780
rect 5480 1770 6040 1780
rect 6320 1770 6360 1780
rect 6400 1770 6560 1780
rect 6800 1770 6840 1780
rect 7800 1770 7840 1780
rect 8400 1770 8480 1780
rect 9720 1770 9760 1780
rect 9920 1770 9960 1780
rect 2440 1760 2520 1770
rect 3240 1760 3280 1770
rect 4360 1760 4400 1770
rect 4520 1760 4560 1770
rect 4600 1760 4640 1770
rect 4760 1760 4840 1770
rect 4880 1760 4960 1770
rect 5080 1760 5120 1770
rect 5160 1760 5200 1770
rect 5320 1760 5400 1770
rect 5480 1760 6040 1770
rect 6320 1760 6360 1770
rect 6400 1760 6560 1770
rect 6800 1760 6840 1770
rect 7800 1760 7840 1770
rect 8400 1760 8480 1770
rect 9720 1760 9760 1770
rect 9920 1760 9960 1770
rect 2440 1750 2520 1760
rect 3240 1750 3280 1760
rect 4360 1750 4400 1760
rect 4520 1750 4560 1760
rect 4600 1750 4640 1760
rect 4760 1750 4840 1760
rect 4880 1750 4960 1760
rect 5080 1750 5120 1760
rect 5160 1750 5200 1760
rect 5320 1750 5400 1760
rect 5480 1750 6040 1760
rect 6320 1750 6360 1760
rect 6400 1750 6560 1760
rect 6800 1750 6840 1760
rect 7800 1750 7840 1760
rect 8400 1750 8480 1760
rect 9720 1750 9760 1760
rect 9920 1750 9960 1760
rect 2440 1740 2520 1750
rect 3240 1740 3280 1750
rect 4360 1740 4400 1750
rect 4520 1740 4560 1750
rect 4600 1740 4640 1750
rect 4760 1740 4840 1750
rect 4880 1740 4960 1750
rect 5080 1740 5120 1750
rect 5160 1740 5200 1750
rect 5320 1740 5400 1750
rect 5480 1740 6040 1750
rect 6320 1740 6360 1750
rect 6400 1740 6560 1750
rect 6800 1740 6840 1750
rect 7800 1740 7840 1750
rect 8400 1740 8480 1750
rect 9720 1740 9760 1750
rect 9920 1740 9960 1750
rect 1880 1730 1920 1740
rect 3240 1730 3280 1740
rect 4040 1730 4080 1740
rect 4520 1730 4760 1740
rect 4800 1730 4840 1740
rect 4880 1730 4960 1740
rect 5000 1730 5120 1740
rect 5160 1730 5240 1740
rect 5320 1730 5360 1740
rect 5400 1730 5480 1740
rect 5560 1730 6040 1740
rect 6320 1730 6560 1740
rect 6800 1730 6840 1740
rect 7800 1730 7840 1740
rect 8360 1730 8520 1740
rect 9160 1730 9200 1740
rect 9720 1730 9760 1740
rect 1880 1720 1920 1730
rect 3240 1720 3280 1730
rect 4040 1720 4080 1730
rect 4520 1720 4760 1730
rect 4800 1720 4840 1730
rect 4880 1720 4960 1730
rect 5000 1720 5120 1730
rect 5160 1720 5240 1730
rect 5320 1720 5360 1730
rect 5400 1720 5480 1730
rect 5560 1720 6040 1730
rect 6320 1720 6560 1730
rect 6800 1720 6840 1730
rect 7800 1720 7840 1730
rect 8360 1720 8520 1730
rect 9160 1720 9200 1730
rect 9720 1720 9760 1730
rect 1880 1710 1920 1720
rect 3240 1710 3280 1720
rect 4040 1710 4080 1720
rect 4520 1710 4760 1720
rect 4800 1710 4840 1720
rect 4880 1710 4960 1720
rect 5000 1710 5120 1720
rect 5160 1710 5240 1720
rect 5320 1710 5360 1720
rect 5400 1710 5480 1720
rect 5560 1710 6040 1720
rect 6320 1710 6560 1720
rect 6800 1710 6840 1720
rect 7800 1710 7840 1720
rect 8360 1710 8520 1720
rect 9160 1710 9200 1720
rect 9720 1710 9760 1720
rect 1880 1700 1920 1710
rect 3240 1700 3280 1710
rect 4040 1700 4080 1710
rect 4520 1700 4760 1710
rect 4800 1700 4840 1710
rect 4880 1700 4960 1710
rect 5000 1700 5120 1710
rect 5160 1700 5240 1710
rect 5320 1700 5360 1710
rect 5400 1700 5480 1710
rect 5560 1700 6040 1710
rect 6320 1700 6560 1710
rect 6800 1700 6840 1710
rect 7800 1700 7840 1710
rect 8360 1700 8520 1710
rect 9160 1700 9200 1710
rect 9720 1700 9760 1710
rect 1880 1690 1920 1700
rect 3200 1690 3240 1700
rect 4240 1690 4280 1700
rect 4400 1690 4440 1700
rect 4480 1690 4520 1700
rect 4560 1690 4840 1700
rect 4880 1690 4960 1700
rect 5000 1690 5080 1700
rect 5120 1690 5200 1700
rect 5280 1690 5320 1700
rect 5480 1690 5520 1700
rect 5560 1690 6000 1700
rect 6320 1690 6520 1700
rect 6800 1690 6840 1700
rect 7800 1690 7880 1700
rect 8400 1690 8520 1700
rect 9120 1690 9200 1700
rect 9880 1690 9920 1700
rect 1880 1680 1920 1690
rect 3200 1680 3240 1690
rect 4240 1680 4280 1690
rect 4400 1680 4440 1690
rect 4480 1680 4520 1690
rect 4560 1680 4840 1690
rect 4880 1680 4960 1690
rect 5000 1680 5080 1690
rect 5120 1680 5200 1690
rect 5280 1680 5320 1690
rect 5480 1680 5520 1690
rect 5560 1680 6000 1690
rect 6320 1680 6520 1690
rect 6800 1680 6840 1690
rect 7800 1680 7880 1690
rect 8400 1680 8520 1690
rect 9120 1680 9200 1690
rect 9880 1680 9920 1690
rect 1880 1670 1920 1680
rect 3200 1670 3240 1680
rect 4240 1670 4280 1680
rect 4400 1670 4440 1680
rect 4480 1670 4520 1680
rect 4560 1670 4840 1680
rect 4880 1670 4960 1680
rect 5000 1670 5080 1680
rect 5120 1670 5200 1680
rect 5280 1670 5320 1680
rect 5480 1670 5520 1680
rect 5560 1670 6000 1680
rect 6320 1670 6520 1680
rect 6800 1670 6840 1680
rect 7800 1670 7880 1680
rect 8400 1670 8520 1680
rect 9120 1670 9200 1680
rect 9880 1670 9920 1680
rect 1880 1660 1920 1670
rect 3200 1660 3240 1670
rect 4240 1660 4280 1670
rect 4400 1660 4440 1670
rect 4480 1660 4520 1670
rect 4560 1660 4840 1670
rect 4880 1660 4960 1670
rect 5000 1660 5080 1670
rect 5120 1660 5200 1670
rect 5280 1660 5320 1670
rect 5480 1660 5520 1670
rect 5560 1660 6000 1670
rect 6320 1660 6520 1670
rect 6800 1660 6840 1670
rect 7800 1660 7880 1670
rect 8400 1660 8520 1670
rect 9120 1660 9200 1670
rect 9880 1660 9920 1670
rect 3200 1650 3240 1660
rect 4080 1650 4200 1660
rect 4400 1650 4480 1660
rect 4520 1650 4560 1660
rect 4600 1650 4640 1660
rect 4720 1650 4760 1660
rect 4800 1650 4960 1660
rect 5000 1650 5080 1660
rect 5120 1650 5200 1660
rect 5360 1650 5400 1660
rect 5560 1650 6000 1660
rect 6320 1650 6520 1660
rect 6800 1650 6840 1660
rect 7800 1650 7880 1660
rect 8320 1650 8480 1660
rect 9120 1650 9200 1660
rect 3200 1640 3240 1650
rect 4080 1640 4200 1650
rect 4400 1640 4480 1650
rect 4520 1640 4560 1650
rect 4600 1640 4640 1650
rect 4720 1640 4760 1650
rect 4800 1640 4960 1650
rect 5000 1640 5080 1650
rect 5120 1640 5200 1650
rect 5360 1640 5400 1650
rect 5560 1640 6000 1650
rect 6320 1640 6520 1650
rect 6800 1640 6840 1650
rect 7800 1640 7880 1650
rect 8320 1640 8480 1650
rect 9120 1640 9200 1650
rect 3200 1630 3240 1640
rect 4080 1630 4200 1640
rect 4400 1630 4480 1640
rect 4520 1630 4560 1640
rect 4600 1630 4640 1640
rect 4720 1630 4760 1640
rect 4800 1630 4960 1640
rect 5000 1630 5080 1640
rect 5120 1630 5200 1640
rect 5360 1630 5400 1640
rect 5560 1630 6000 1640
rect 6320 1630 6520 1640
rect 6800 1630 6840 1640
rect 7800 1630 7880 1640
rect 8320 1630 8480 1640
rect 9120 1630 9200 1640
rect 3200 1620 3240 1630
rect 4080 1620 4200 1630
rect 4400 1620 4480 1630
rect 4520 1620 4560 1630
rect 4600 1620 4640 1630
rect 4720 1620 4760 1630
rect 4800 1620 4960 1630
rect 5000 1620 5080 1630
rect 5120 1620 5200 1630
rect 5360 1620 5400 1630
rect 5560 1620 6000 1630
rect 6320 1620 6520 1630
rect 6800 1620 6840 1630
rect 7800 1620 7880 1630
rect 8320 1620 8480 1630
rect 9120 1620 9200 1630
rect 1920 1610 1960 1620
rect 3160 1610 3200 1620
rect 4120 1610 4200 1620
rect 4280 1610 4320 1620
rect 4840 1610 5160 1620
rect 5240 1610 5280 1620
rect 5320 1610 5360 1620
rect 5520 1610 5560 1620
rect 5680 1610 5960 1620
rect 6320 1610 6440 1620
rect 6800 1610 6840 1620
rect 7800 1610 7880 1620
rect 8360 1610 8440 1620
rect 9840 1610 9880 1620
rect 1920 1600 1960 1610
rect 3160 1600 3200 1610
rect 4120 1600 4200 1610
rect 4280 1600 4320 1610
rect 4840 1600 5160 1610
rect 5240 1600 5280 1610
rect 5320 1600 5360 1610
rect 5520 1600 5560 1610
rect 5680 1600 5960 1610
rect 6320 1600 6440 1610
rect 6800 1600 6840 1610
rect 7800 1600 7880 1610
rect 8360 1600 8440 1610
rect 9840 1600 9880 1610
rect 1920 1590 1960 1600
rect 3160 1590 3200 1600
rect 4120 1590 4200 1600
rect 4280 1590 4320 1600
rect 4840 1590 5160 1600
rect 5240 1590 5280 1600
rect 5320 1590 5360 1600
rect 5520 1590 5560 1600
rect 5680 1590 5960 1600
rect 6320 1590 6440 1600
rect 6800 1590 6840 1600
rect 7800 1590 7880 1600
rect 8360 1590 8440 1600
rect 9840 1590 9880 1600
rect 1920 1580 1960 1590
rect 3160 1580 3200 1590
rect 4120 1580 4200 1590
rect 4280 1580 4320 1590
rect 4840 1580 5160 1590
rect 5240 1580 5280 1590
rect 5320 1580 5360 1590
rect 5520 1580 5560 1590
rect 5680 1580 5960 1590
rect 6320 1580 6440 1590
rect 6800 1580 6840 1590
rect 7800 1580 7880 1590
rect 8360 1580 8440 1590
rect 9840 1580 9880 1590
rect 1960 1570 2000 1580
rect 3120 1570 3200 1580
rect 4120 1570 4240 1580
rect 4800 1570 5240 1580
rect 5320 1570 5560 1580
rect 5600 1570 5640 1580
rect 5720 1570 5960 1580
rect 6320 1570 6400 1580
rect 6800 1570 6840 1580
rect 7840 1570 7880 1580
rect 8400 1570 8440 1580
rect 9760 1570 9840 1580
rect 9960 1570 9990 1580
rect 1960 1560 2000 1570
rect 3120 1560 3200 1570
rect 4120 1560 4240 1570
rect 4800 1560 5240 1570
rect 5320 1560 5560 1570
rect 5600 1560 5640 1570
rect 5720 1560 5960 1570
rect 6320 1560 6400 1570
rect 6800 1560 6840 1570
rect 7840 1560 7880 1570
rect 8400 1560 8440 1570
rect 9760 1560 9840 1570
rect 9960 1560 9990 1570
rect 1960 1550 2000 1560
rect 3120 1550 3200 1560
rect 4120 1550 4240 1560
rect 4800 1550 5240 1560
rect 5320 1550 5560 1560
rect 5600 1550 5640 1560
rect 5720 1550 5960 1560
rect 6320 1550 6400 1560
rect 6800 1550 6840 1560
rect 7840 1550 7880 1560
rect 8400 1550 8440 1560
rect 9760 1550 9840 1560
rect 9960 1550 9990 1560
rect 1960 1540 2000 1550
rect 3120 1540 3200 1550
rect 4120 1540 4240 1550
rect 4800 1540 5240 1550
rect 5320 1540 5560 1550
rect 5600 1540 5640 1550
rect 5720 1540 5960 1550
rect 6320 1540 6400 1550
rect 6800 1540 6840 1550
rect 7840 1540 7880 1550
rect 8400 1540 8440 1550
rect 9760 1540 9840 1550
rect 9960 1540 9990 1550
rect 3080 1530 3160 1540
rect 4120 1530 4240 1540
rect 4920 1530 5280 1540
rect 5320 1530 5560 1540
rect 5640 1530 5680 1540
rect 5720 1530 5960 1540
rect 6320 1530 6400 1540
rect 6800 1530 6840 1540
rect 7360 1530 7400 1540
rect 7840 1530 7880 1540
rect 8360 1530 8440 1540
rect 9720 1530 9760 1540
rect 9800 1530 9840 1540
rect 3080 1520 3160 1530
rect 4120 1520 4240 1530
rect 4920 1520 5280 1530
rect 5320 1520 5560 1530
rect 5640 1520 5680 1530
rect 5720 1520 5960 1530
rect 6320 1520 6400 1530
rect 6800 1520 6840 1530
rect 7360 1520 7400 1530
rect 7840 1520 7880 1530
rect 8360 1520 8440 1530
rect 9720 1520 9760 1530
rect 9800 1520 9840 1530
rect 3080 1510 3160 1520
rect 4120 1510 4240 1520
rect 4920 1510 5280 1520
rect 5320 1510 5560 1520
rect 5640 1510 5680 1520
rect 5720 1510 5960 1520
rect 6320 1510 6400 1520
rect 6800 1510 6840 1520
rect 7360 1510 7400 1520
rect 7840 1510 7880 1520
rect 8360 1510 8440 1520
rect 9720 1510 9760 1520
rect 9800 1510 9840 1520
rect 3080 1500 3160 1510
rect 4120 1500 4240 1510
rect 4920 1500 5280 1510
rect 5320 1500 5560 1510
rect 5640 1500 5680 1510
rect 5720 1500 5960 1510
rect 6320 1500 6400 1510
rect 6800 1500 6840 1510
rect 7360 1500 7400 1510
rect 7840 1500 7880 1510
rect 8360 1500 8440 1510
rect 9720 1500 9760 1510
rect 9800 1500 9840 1510
rect 2000 1490 2040 1500
rect 2960 1490 3000 1500
rect 3040 1490 3120 1500
rect 4120 1490 4160 1500
rect 5000 1490 5440 1500
rect 5520 1490 5560 1500
rect 5640 1490 5680 1500
rect 5720 1490 5880 1500
rect 6320 1490 6360 1500
rect 7360 1490 7400 1500
rect 7840 1490 7880 1500
rect 8280 1490 8320 1500
rect 8360 1490 8440 1500
rect 2000 1480 2040 1490
rect 2960 1480 3000 1490
rect 3040 1480 3120 1490
rect 4120 1480 4160 1490
rect 5000 1480 5440 1490
rect 5520 1480 5560 1490
rect 5640 1480 5680 1490
rect 5720 1480 5880 1490
rect 6320 1480 6360 1490
rect 7360 1480 7400 1490
rect 7840 1480 7880 1490
rect 8280 1480 8320 1490
rect 8360 1480 8440 1490
rect 2000 1470 2040 1480
rect 2960 1470 3000 1480
rect 3040 1470 3120 1480
rect 4120 1470 4160 1480
rect 5000 1470 5440 1480
rect 5520 1470 5560 1480
rect 5640 1470 5680 1480
rect 5720 1470 5880 1480
rect 6320 1470 6360 1480
rect 7360 1470 7400 1480
rect 7840 1470 7880 1480
rect 8280 1470 8320 1480
rect 8360 1470 8440 1480
rect 2000 1460 2040 1470
rect 2960 1460 3000 1470
rect 3040 1460 3120 1470
rect 4120 1460 4160 1470
rect 5000 1460 5440 1470
rect 5520 1460 5560 1470
rect 5640 1460 5680 1470
rect 5720 1460 5880 1470
rect 6320 1460 6360 1470
rect 7360 1460 7400 1470
rect 7840 1460 7880 1470
rect 8280 1460 8320 1470
rect 8360 1460 8440 1470
rect 880 1450 1000 1460
rect 2040 1450 2080 1460
rect 2920 1450 3040 1460
rect 4360 1450 4400 1460
rect 5040 1450 5440 1460
rect 5560 1450 5600 1460
rect 5640 1450 5880 1460
rect 7360 1450 7400 1460
rect 7840 1450 7880 1460
rect 8280 1450 8320 1460
rect 8360 1450 8440 1460
rect 880 1440 1000 1450
rect 2040 1440 2080 1450
rect 2920 1440 3040 1450
rect 4360 1440 4400 1450
rect 5040 1440 5440 1450
rect 5560 1440 5600 1450
rect 5640 1440 5880 1450
rect 7360 1440 7400 1450
rect 7840 1440 7880 1450
rect 8280 1440 8320 1450
rect 8360 1440 8440 1450
rect 880 1430 1000 1440
rect 2040 1430 2080 1440
rect 2920 1430 3040 1440
rect 4360 1430 4400 1440
rect 5040 1430 5440 1440
rect 5560 1430 5600 1440
rect 5640 1430 5880 1440
rect 7360 1430 7400 1440
rect 7840 1430 7880 1440
rect 8280 1430 8320 1440
rect 8360 1430 8440 1440
rect 880 1420 1000 1430
rect 2040 1420 2080 1430
rect 2920 1420 3040 1430
rect 4360 1420 4400 1430
rect 5040 1420 5440 1430
rect 5560 1420 5600 1430
rect 5640 1420 5880 1430
rect 7360 1420 7400 1430
rect 7840 1420 7880 1430
rect 8280 1420 8320 1430
rect 8360 1420 8440 1430
rect 840 1410 1000 1420
rect 2080 1410 2120 1420
rect 2880 1410 3000 1420
rect 5120 1410 5440 1420
rect 5520 1410 5560 1420
rect 5600 1410 5920 1420
rect 7360 1410 7400 1420
rect 7840 1410 7920 1420
rect 8360 1410 8440 1420
rect 9680 1410 9720 1420
rect 840 1400 1000 1410
rect 2080 1400 2120 1410
rect 2880 1400 3000 1410
rect 5120 1400 5440 1410
rect 5520 1400 5560 1410
rect 5600 1400 5920 1410
rect 7360 1400 7400 1410
rect 7840 1400 7920 1410
rect 8360 1400 8440 1410
rect 9680 1400 9720 1410
rect 840 1390 1000 1400
rect 2080 1390 2120 1400
rect 2880 1390 3000 1400
rect 5120 1390 5440 1400
rect 5520 1390 5560 1400
rect 5600 1390 5920 1400
rect 7360 1390 7400 1400
rect 7840 1390 7920 1400
rect 8360 1390 8440 1400
rect 9680 1390 9720 1400
rect 840 1380 1000 1390
rect 2080 1380 2120 1390
rect 2880 1380 3000 1390
rect 5120 1380 5440 1390
rect 5520 1380 5560 1390
rect 5600 1380 5920 1390
rect 7360 1380 7400 1390
rect 7840 1380 7920 1390
rect 8360 1380 8440 1390
rect 9680 1380 9720 1390
rect 840 1370 960 1380
rect 2120 1370 2200 1380
rect 2840 1370 2960 1380
rect 3600 1370 3640 1380
rect 4160 1370 4240 1380
rect 5120 1370 5520 1380
rect 5600 1370 5920 1380
rect 6800 1370 6840 1380
rect 7840 1370 7920 1380
rect 8240 1370 8280 1380
rect 8320 1370 8440 1380
rect 840 1360 960 1370
rect 2120 1360 2200 1370
rect 2840 1360 2960 1370
rect 3600 1360 3640 1370
rect 4160 1360 4240 1370
rect 5120 1360 5520 1370
rect 5600 1360 5920 1370
rect 6800 1360 6840 1370
rect 7840 1360 7920 1370
rect 8240 1360 8280 1370
rect 8320 1360 8440 1370
rect 840 1350 960 1360
rect 2120 1350 2200 1360
rect 2840 1350 2960 1360
rect 3600 1350 3640 1360
rect 4160 1350 4240 1360
rect 5120 1350 5520 1360
rect 5600 1350 5920 1360
rect 6800 1350 6840 1360
rect 7840 1350 7920 1360
rect 8240 1350 8280 1360
rect 8320 1350 8440 1360
rect 840 1340 960 1350
rect 2120 1340 2200 1350
rect 2840 1340 2960 1350
rect 3600 1340 3640 1350
rect 4160 1340 4240 1350
rect 5120 1340 5520 1350
rect 5600 1340 5920 1350
rect 6800 1340 6840 1350
rect 7840 1340 7920 1350
rect 8240 1340 8280 1350
rect 8320 1340 8440 1350
rect 840 1330 920 1340
rect 2160 1330 2240 1340
rect 2760 1330 2800 1340
rect 4400 1330 4440 1340
rect 5040 1330 5200 1340
rect 5240 1330 5440 1340
rect 5480 1330 5920 1340
rect 6800 1330 6840 1340
rect 7840 1330 7920 1340
rect 8200 1330 8440 1340
rect 9160 1330 9240 1340
rect 9680 1330 9720 1340
rect 9800 1330 9840 1340
rect 840 1320 920 1330
rect 2160 1320 2240 1330
rect 2760 1320 2800 1330
rect 4400 1320 4440 1330
rect 5040 1320 5200 1330
rect 5240 1320 5440 1330
rect 5480 1320 5920 1330
rect 6800 1320 6840 1330
rect 7840 1320 7920 1330
rect 8200 1320 8440 1330
rect 9160 1320 9240 1330
rect 9680 1320 9720 1330
rect 9800 1320 9840 1330
rect 840 1310 920 1320
rect 2160 1310 2240 1320
rect 2760 1310 2800 1320
rect 4400 1310 4440 1320
rect 5040 1310 5200 1320
rect 5240 1310 5440 1320
rect 5480 1310 5920 1320
rect 6800 1310 6840 1320
rect 7840 1310 7920 1320
rect 8200 1310 8440 1320
rect 9160 1310 9240 1320
rect 9680 1310 9720 1320
rect 9800 1310 9840 1320
rect 840 1300 920 1310
rect 2160 1300 2240 1310
rect 2760 1300 2800 1310
rect 4400 1300 4440 1310
rect 5040 1300 5200 1310
rect 5240 1300 5440 1310
rect 5480 1300 5920 1310
rect 6800 1300 6840 1310
rect 7840 1300 7920 1310
rect 8200 1300 8440 1310
rect 9160 1300 9240 1310
rect 9680 1300 9720 1310
rect 9800 1300 9840 1310
rect 800 1290 920 1300
rect 2200 1290 2440 1300
rect 2680 1290 2720 1300
rect 3480 1290 3520 1300
rect 4960 1290 5120 1300
rect 5160 1290 5200 1300
rect 5240 1290 5920 1300
rect 6800 1290 6840 1300
rect 7880 1290 7920 1300
rect 8160 1290 8440 1300
rect 9080 1290 9120 1300
rect 9160 1290 9200 1300
rect 9240 1290 9280 1300
rect 9760 1290 9840 1300
rect 800 1280 920 1290
rect 2200 1280 2440 1290
rect 2680 1280 2720 1290
rect 3480 1280 3520 1290
rect 4960 1280 5120 1290
rect 5160 1280 5200 1290
rect 5240 1280 5920 1290
rect 6800 1280 6840 1290
rect 7880 1280 7920 1290
rect 8160 1280 8440 1290
rect 9080 1280 9120 1290
rect 9160 1280 9200 1290
rect 9240 1280 9280 1290
rect 9760 1280 9840 1290
rect 800 1270 920 1280
rect 2200 1270 2440 1280
rect 2680 1270 2720 1280
rect 3480 1270 3520 1280
rect 4960 1270 5120 1280
rect 5160 1270 5200 1280
rect 5240 1270 5920 1280
rect 6800 1270 6840 1280
rect 7880 1270 7920 1280
rect 8160 1270 8440 1280
rect 9080 1270 9120 1280
rect 9160 1270 9200 1280
rect 9240 1270 9280 1280
rect 9760 1270 9840 1280
rect 800 1260 920 1270
rect 2200 1260 2440 1270
rect 2680 1260 2720 1270
rect 3480 1260 3520 1270
rect 4960 1260 5120 1270
rect 5160 1260 5200 1270
rect 5240 1260 5920 1270
rect 6800 1260 6840 1270
rect 7880 1260 7920 1270
rect 8160 1260 8440 1270
rect 9080 1260 9120 1270
rect 9160 1260 9200 1270
rect 9240 1260 9280 1270
rect 9760 1260 9840 1270
rect 800 1250 920 1260
rect 2240 1250 2640 1260
rect 3760 1250 3800 1260
rect 5000 1250 5200 1260
rect 5440 1250 5920 1260
rect 6760 1250 6840 1260
rect 7880 1250 7960 1260
rect 8200 1250 8440 1260
rect 8960 1250 9000 1260
rect 9080 1250 9120 1260
rect 9240 1250 9280 1260
rect 9640 1250 9680 1260
rect 9760 1250 9800 1260
rect 9960 1250 9990 1260
rect 800 1240 920 1250
rect 2240 1240 2640 1250
rect 3760 1240 3800 1250
rect 5000 1240 5200 1250
rect 5440 1240 5920 1250
rect 6760 1240 6840 1250
rect 7880 1240 7960 1250
rect 8200 1240 8440 1250
rect 8960 1240 9000 1250
rect 9080 1240 9120 1250
rect 9240 1240 9280 1250
rect 9640 1240 9680 1250
rect 9760 1240 9800 1250
rect 9960 1240 9990 1250
rect 800 1230 920 1240
rect 2240 1230 2640 1240
rect 3760 1230 3800 1240
rect 5000 1230 5200 1240
rect 5440 1230 5920 1240
rect 6760 1230 6840 1240
rect 7880 1230 7960 1240
rect 8200 1230 8440 1240
rect 8960 1230 9000 1240
rect 9080 1230 9120 1240
rect 9240 1230 9280 1240
rect 9640 1230 9680 1240
rect 9760 1230 9800 1240
rect 9960 1230 9990 1240
rect 800 1220 920 1230
rect 2240 1220 2640 1230
rect 3760 1220 3800 1230
rect 5000 1220 5200 1230
rect 5440 1220 5920 1230
rect 6760 1220 6840 1230
rect 7880 1220 7960 1230
rect 8200 1220 8440 1230
rect 8960 1220 9000 1230
rect 9080 1220 9120 1230
rect 9240 1220 9280 1230
rect 9640 1220 9680 1230
rect 9760 1220 9800 1230
rect 9960 1220 9990 1230
rect 800 1210 880 1220
rect 2120 1210 2240 1220
rect 2320 1210 2600 1220
rect 3520 1210 3680 1220
rect 4440 1210 4480 1220
rect 4720 1210 4920 1220
rect 4960 1210 5000 1220
rect 5080 1210 5120 1220
rect 5160 1210 5200 1220
rect 5240 1210 5320 1220
rect 5360 1210 5920 1220
rect 6680 1210 6720 1220
rect 6800 1210 6840 1220
rect 7880 1210 7960 1220
rect 8200 1210 8400 1220
rect 8840 1210 9000 1220
rect 9040 1210 9120 1220
rect 9160 1210 9200 1220
rect 9240 1210 9280 1220
rect 9600 1210 9640 1220
rect 9720 1210 9760 1220
rect 800 1200 880 1210
rect 2120 1200 2240 1210
rect 2320 1200 2600 1210
rect 3520 1200 3680 1210
rect 4440 1200 4480 1210
rect 4720 1200 4920 1210
rect 4960 1200 5000 1210
rect 5080 1200 5120 1210
rect 5160 1200 5200 1210
rect 5240 1200 5320 1210
rect 5360 1200 5920 1210
rect 6680 1200 6720 1210
rect 6800 1200 6840 1210
rect 7880 1200 7960 1210
rect 8200 1200 8400 1210
rect 8840 1200 9000 1210
rect 9040 1200 9120 1210
rect 9160 1200 9200 1210
rect 9240 1200 9280 1210
rect 9600 1200 9640 1210
rect 9720 1200 9760 1210
rect 800 1190 880 1200
rect 2120 1190 2240 1200
rect 2320 1190 2600 1200
rect 3520 1190 3680 1200
rect 4440 1190 4480 1200
rect 4720 1190 4920 1200
rect 4960 1190 5000 1200
rect 5080 1190 5120 1200
rect 5160 1190 5200 1200
rect 5240 1190 5320 1200
rect 5360 1190 5920 1200
rect 6680 1190 6720 1200
rect 6800 1190 6840 1200
rect 7880 1190 7960 1200
rect 8200 1190 8400 1200
rect 8840 1190 9000 1200
rect 9040 1190 9120 1200
rect 9160 1190 9200 1200
rect 9240 1190 9280 1200
rect 9600 1190 9640 1200
rect 9720 1190 9760 1200
rect 800 1180 880 1190
rect 2120 1180 2240 1190
rect 2320 1180 2600 1190
rect 3520 1180 3680 1190
rect 4440 1180 4480 1190
rect 4720 1180 4920 1190
rect 4960 1180 5000 1190
rect 5080 1180 5120 1190
rect 5160 1180 5200 1190
rect 5240 1180 5320 1190
rect 5360 1180 5920 1190
rect 6680 1180 6720 1190
rect 6800 1180 6840 1190
rect 7880 1180 7960 1190
rect 8200 1180 8400 1190
rect 8840 1180 9000 1190
rect 9040 1180 9120 1190
rect 9160 1180 9200 1190
rect 9240 1180 9280 1190
rect 9600 1180 9640 1190
rect 9720 1180 9760 1190
rect 760 1170 800 1180
rect 840 1170 880 1180
rect 2080 1170 2280 1180
rect 3560 1170 3720 1180
rect 3880 1170 3920 1180
rect 4560 1170 4760 1180
rect 4840 1170 4920 1180
rect 5000 1170 5040 1180
rect 5360 1170 5920 1180
rect 6640 1170 6680 1180
rect 6800 1170 6840 1180
rect 7920 1170 7960 1180
rect 8160 1170 8360 1180
rect 8720 1170 9120 1180
rect 9160 1170 9200 1180
rect 9240 1170 9280 1180
rect 9600 1170 9640 1180
rect 9720 1170 9760 1180
rect 760 1160 800 1170
rect 840 1160 880 1170
rect 2080 1160 2280 1170
rect 3560 1160 3720 1170
rect 3880 1160 3920 1170
rect 4560 1160 4760 1170
rect 4840 1160 4920 1170
rect 5000 1160 5040 1170
rect 5360 1160 5920 1170
rect 6640 1160 6680 1170
rect 6800 1160 6840 1170
rect 7920 1160 7960 1170
rect 8160 1160 8360 1170
rect 8720 1160 9120 1170
rect 9160 1160 9200 1170
rect 9240 1160 9280 1170
rect 9600 1160 9640 1170
rect 9720 1160 9760 1170
rect 760 1150 800 1160
rect 840 1150 880 1160
rect 2080 1150 2280 1160
rect 3560 1150 3720 1160
rect 3880 1150 3920 1160
rect 4560 1150 4760 1160
rect 4840 1150 4920 1160
rect 5000 1150 5040 1160
rect 5360 1150 5920 1160
rect 6640 1150 6680 1160
rect 6800 1150 6840 1160
rect 7920 1150 7960 1160
rect 8160 1150 8360 1160
rect 8720 1150 9120 1160
rect 9160 1150 9200 1160
rect 9240 1150 9280 1160
rect 9600 1150 9640 1160
rect 9720 1150 9760 1160
rect 760 1140 800 1150
rect 840 1140 880 1150
rect 2080 1140 2280 1150
rect 3560 1140 3720 1150
rect 3880 1140 3920 1150
rect 4560 1140 4760 1150
rect 4840 1140 4920 1150
rect 5000 1140 5040 1150
rect 5360 1140 5920 1150
rect 6640 1140 6680 1150
rect 6800 1140 6840 1150
rect 7920 1140 7960 1150
rect 8160 1140 8360 1150
rect 8720 1140 9120 1150
rect 9160 1140 9200 1150
rect 9240 1140 9280 1150
rect 9600 1140 9640 1150
rect 9720 1140 9760 1150
rect 840 1130 880 1140
rect 2040 1130 2360 1140
rect 3600 1130 3720 1140
rect 4200 1130 4240 1140
rect 4560 1130 4760 1140
rect 5400 1130 5680 1140
rect 5720 1130 5920 1140
rect 6560 1130 6600 1140
rect 6800 1130 6840 1140
rect 7920 1130 7960 1140
rect 8160 1130 8360 1140
rect 8680 1130 9120 1140
rect 9160 1130 9280 1140
rect 9560 1130 9600 1140
rect 9720 1130 9760 1140
rect 9800 1130 9840 1140
rect 840 1120 880 1130
rect 2040 1120 2360 1130
rect 3600 1120 3720 1130
rect 4200 1120 4240 1130
rect 4560 1120 4760 1130
rect 5400 1120 5680 1130
rect 5720 1120 5920 1130
rect 6560 1120 6600 1130
rect 6800 1120 6840 1130
rect 7920 1120 7960 1130
rect 8160 1120 8360 1130
rect 8680 1120 9120 1130
rect 9160 1120 9280 1130
rect 9560 1120 9600 1130
rect 9720 1120 9760 1130
rect 9800 1120 9840 1130
rect 840 1110 880 1120
rect 2040 1110 2360 1120
rect 3600 1110 3720 1120
rect 4200 1110 4240 1120
rect 4560 1110 4760 1120
rect 5400 1110 5680 1120
rect 5720 1110 5920 1120
rect 6560 1110 6600 1120
rect 6800 1110 6840 1120
rect 7920 1110 7960 1120
rect 8160 1110 8360 1120
rect 8680 1110 9120 1120
rect 9160 1110 9280 1120
rect 9560 1110 9600 1120
rect 9720 1110 9760 1120
rect 9800 1110 9840 1120
rect 840 1100 880 1110
rect 2040 1100 2360 1110
rect 3600 1100 3720 1110
rect 4200 1100 4240 1110
rect 4560 1100 4760 1110
rect 5400 1100 5680 1110
rect 5720 1100 5920 1110
rect 6560 1100 6600 1110
rect 6800 1100 6840 1110
rect 7920 1100 7960 1110
rect 8160 1100 8360 1110
rect 8680 1100 9120 1110
rect 9160 1100 9280 1110
rect 9560 1100 9600 1110
rect 9720 1100 9760 1110
rect 9800 1100 9840 1110
rect 840 1090 880 1100
rect 2000 1090 2840 1100
rect 3640 1090 3680 1100
rect 4000 1090 4040 1100
rect 4200 1090 4240 1100
rect 5480 1090 5640 1100
rect 5880 1090 5960 1100
rect 6480 1090 6520 1100
rect 6800 1090 6840 1100
rect 7920 1090 7960 1100
rect 8160 1090 8360 1100
rect 8680 1090 9120 1100
rect 9720 1090 9760 1100
rect 9800 1090 9840 1100
rect 840 1080 880 1090
rect 2000 1080 2840 1090
rect 3640 1080 3680 1090
rect 4000 1080 4040 1090
rect 4200 1080 4240 1090
rect 5480 1080 5640 1090
rect 5880 1080 5960 1090
rect 6480 1080 6520 1090
rect 6800 1080 6840 1090
rect 7920 1080 7960 1090
rect 8160 1080 8360 1090
rect 8680 1080 9120 1090
rect 9720 1080 9760 1090
rect 9800 1080 9840 1090
rect 840 1070 880 1080
rect 2000 1070 2840 1080
rect 3640 1070 3680 1080
rect 4000 1070 4040 1080
rect 4200 1070 4240 1080
rect 5480 1070 5640 1080
rect 5880 1070 5960 1080
rect 6480 1070 6520 1080
rect 6800 1070 6840 1080
rect 7920 1070 7960 1080
rect 8160 1070 8360 1080
rect 8680 1070 9120 1080
rect 9720 1070 9760 1080
rect 9800 1070 9840 1080
rect 840 1060 880 1070
rect 2000 1060 2840 1070
rect 3640 1060 3680 1070
rect 4000 1060 4040 1070
rect 4200 1060 4240 1070
rect 5480 1060 5640 1070
rect 5880 1060 5960 1070
rect 6480 1060 6520 1070
rect 6800 1060 6840 1070
rect 7920 1060 7960 1070
rect 8160 1060 8360 1070
rect 8680 1060 9120 1070
rect 9720 1060 9760 1070
rect 9800 1060 9840 1070
rect 720 1050 760 1060
rect 800 1050 840 1060
rect 1520 1050 1640 1060
rect 2000 1050 2080 1060
rect 2200 1050 2840 1060
rect 3680 1050 3720 1060
rect 3760 1050 3840 1060
rect 4600 1050 4640 1060
rect 5480 1050 5520 1060
rect 5840 1050 5880 1060
rect 6440 1050 6480 1060
rect 6800 1050 6840 1060
rect 7400 1050 7440 1060
rect 7920 1050 7960 1060
rect 8160 1050 8360 1060
rect 8560 1050 9120 1060
rect 9520 1050 9560 1060
rect 9800 1050 9840 1060
rect 720 1040 760 1050
rect 800 1040 840 1050
rect 1520 1040 1640 1050
rect 2000 1040 2080 1050
rect 2200 1040 2840 1050
rect 3680 1040 3720 1050
rect 3760 1040 3840 1050
rect 4600 1040 4640 1050
rect 5480 1040 5520 1050
rect 5840 1040 5880 1050
rect 6440 1040 6480 1050
rect 6800 1040 6840 1050
rect 7400 1040 7440 1050
rect 7920 1040 7960 1050
rect 8160 1040 8360 1050
rect 8560 1040 9120 1050
rect 9520 1040 9560 1050
rect 9800 1040 9840 1050
rect 720 1030 760 1040
rect 800 1030 840 1040
rect 1520 1030 1640 1040
rect 2000 1030 2080 1040
rect 2200 1030 2840 1040
rect 3680 1030 3720 1040
rect 3760 1030 3840 1040
rect 4600 1030 4640 1040
rect 5480 1030 5520 1040
rect 5840 1030 5880 1040
rect 6440 1030 6480 1040
rect 6800 1030 6840 1040
rect 7400 1030 7440 1040
rect 7920 1030 7960 1040
rect 8160 1030 8360 1040
rect 8560 1030 9120 1040
rect 9520 1030 9560 1040
rect 9800 1030 9840 1040
rect 720 1020 760 1030
rect 800 1020 840 1030
rect 1520 1020 1640 1030
rect 2000 1020 2080 1030
rect 2200 1020 2840 1030
rect 3680 1020 3720 1030
rect 3760 1020 3840 1030
rect 4600 1020 4640 1030
rect 5480 1020 5520 1030
rect 5840 1020 5880 1030
rect 6440 1020 6480 1030
rect 6800 1020 6840 1030
rect 7400 1020 7440 1030
rect 7920 1020 7960 1030
rect 8160 1020 8360 1030
rect 8560 1020 9120 1030
rect 9520 1020 9560 1030
rect 9800 1020 9840 1030
rect 800 1010 840 1020
rect 1480 1010 1560 1020
rect 2000 1010 2040 1020
rect 2280 1010 2680 1020
rect 2720 1010 2840 1020
rect 3720 1010 3840 1020
rect 4120 1010 4160 1020
rect 5440 1010 5520 1020
rect 5600 1010 5640 1020
rect 6400 1010 6440 1020
rect 6800 1010 6840 1020
rect 7400 1010 7440 1020
rect 7920 1010 7960 1020
rect 8120 1010 8360 1020
rect 8560 1010 9000 1020
rect 9080 1010 9120 1020
rect 9760 1010 9800 1020
rect 800 1000 840 1010
rect 1480 1000 1560 1010
rect 2000 1000 2040 1010
rect 2280 1000 2680 1010
rect 2720 1000 2840 1010
rect 3720 1000 3840 1010
rect 4120 1000 4160 1010
rect 5440 1000 5520 1010
rect 5600 1000 5640 1010
rect 6400 1000 6440 1010
rect 6800 1000 6840 1010
rect 7400 1000 7440 1010
rect 7920 1000 7960 1010
rect 8120 1000 8360 1010
rect 8560 1000 9000 1010
rect 9080 1000 9120 1010
rect 9760 1000 9800 1010
rect 800 990 840 1000
rect 1480 990 1560 1000
rect 2000 990 2040 1000
rect 2280 990 2680 1000
rect 2720 990 2840 1000
rect 3720 990 3840 1000
rect 4120 990 4160 1000
rect 5440 990 5520 1000
rect 5600 990 5640 1000
rect 6400 990 6440 1000
rect 6800 990 6840 1000
rect 7400 990 7440 1000
rect 7920 990 7960 1000
rect 8120 990 8360 1000
rect 8560 990 9000 1000
rect 9080 990 9120 1000
rect 9760 990 9800 1000
rect 800 980 840 990
rect 1480 980 1560 990
rect 2000 980 2040 990
rect 2280 980 2680 990
rect 2720 980 2840 990
rect 3720 980 3840 990
rect 4120 980 4160 990
rect 5440 980 5520 990
rect 5600 980 5640 990
rect 6400 980 6440 990
rect 6800 980 6840 990
rect 7400 980 7440 990
rect 7920 980 7960 990
rect 8120 980 8360 990
rect 8560 980 9000 990
rect 9080 980 9120 990
rect 9760 980 9800 990
rect 1360 970 1400 980
rect 1440 970 1520 980
rect 2000 970 2040 980
rect 2720 970 2840 980
rect 3760 970 3800 980
rect 5320 970 5960 980
rect 6400 970 6480 980
rect 7400 970 7440 980
rect 7920 970 7960 980
rect 8120 970 8160 980
rect 8200 970 8360 980
rect 8560 970 8960 980
rect 9080 970 9160 980
rect 1360 960 1400 970
rect 1440 960 1520 970
rect 2000 960 2040 970
rect 2720 960 2840 970
rect 3760 960 3800 970
rect 5320 960 5960 970
rect 6400 960 6480 970
rect 7400 960 7440 970
rect 7920 960 7960 970
rect 8120 960 8160 970
rect 8200 960 8360 970
rect 8560 960 8960 970
rect 9080 960 9160 970
rect 1360 950 1400 960
rect 1440 950 1520 960
rect 2000 950 2040 960
rect 2720 950 2840 960
rect 3760 950 3800 960
rect 5320 950 5960 960
rect 6400 950 6480 960
rect 7400 950 7440 960
rect 7920 950 7960 960
rect 8120 950 8160 960
rect 8200 950 8360 960
rect 8560 950 8960 960
rect 9080 950 9160 960
rect 1360 940 1400 950
rect 1440 940 1520 950
rect 2000 940 2040 950
rect 2720 940 2840 950
rect 3760 940 3800 950
rect 5320 940 5960 950
rect 6400 940 6480 950
rect 7400 940 7440 950
rect 7920 940 7960 950
rect 8120 940 8160 950
rect 8200 940 8360 950
rect 8560 940 8960 950
rect 9080 940 9160 950
rect 680 930 720 940
rect 760 930 800 940
rect 1320 930 1360 940
rect 1400 930 1480 940
rect 2000 930 2040 940
rect 2720 930 2760 940
rect 5320 930 5360 940
rect 5480 930 5520 940
rect 5560 930 6040 940
rect 6200 930 6280 940
rect 6400 930 6480 940
rect 7400 930 7440 940
rect 8120 930 8160 940
rect 8200 930 8400 940
rect 8600 930 8920 940
rect 9080 930 9160 940
rect 680 920 720 930
rect 760 920 800 930
rect 1320 920 1360 930
rect 1400 920 1480 930
rect 2000 920 2040 930
rect 2720 920 2760 930
rect 5320 920 5360 930
rect 5480 920 5520 930
rect 5560 920 6040 930
rect 6200 920 6280 930
rect 6400 920 6480 930
rect 7400 920 7440 930
rect 8120 920 8160 930
rect 8200 920 8400 930
rect 8600 920 8920 930
rect 9080 920 9160 930
rect 680 910 720 920
rect 760 910 800 920
rect 1320 910 1360 920
rect 1400 910 1480 920
rect 2000 910 2040 920
rect 2720 910 2760 920
rect 5320 910 5360 920
rect 5480 910 5520 920
rect 5560 910 6040 920
rect 6200 910 6280 920
rect 6400 910 6480 920
rect 7400 910 7440 920
rect 8120 910 8160 920
rect 8200 910 8400 920
rect 8600 910 8920 920
rect 9080 910 9160 920
rect 680 900 720 910
rect 760 900 800 910
rect 1320 900 1360 910
rect 1400 900 1480 910
rect 2000 900 2040 910
rect 2720 900 2760 910
rect 5320 900 5360 910
rect 5480 900 5520 910
rect 5560 900 6040 910
rect 6200 900 6280 910
rect 6400 900 6480 910
rect 7400 900 7440 910
rect 8120 900 8160 910
rect 8200 900 8400 910
rect 8600 900 8920 910
rect 9080 900 9160 910
rect 760 890 920 900
rect 1360 890 1440 900
rect 2000 890 2040 900
rect 2680 890 2720 900
rect 5320 890 5360 900
rect 5400 890 5680 900
rect 5800 890 6040 900
rect 6200 890 6280 900
rect 6400 890 6480 900
rect 7400 890 7440 900
rect 7960 890 8000 900
rect 8120 890 8160 900
rect 8200 890 8440 900
rect 8640 890 8880 900
rect 9080 890 9160 900
rect 9440 890 9480 900
rect 760 880 920 890
rect 1360 880 1440 890
rect 2000 880 2040 890
rect 2680 880 2720 890
rect 5320 880 5360 890
rect 5400 880 5680 890
rect 5800 880 6040 890
rect 6200 880 6280 890
rect 6400 880 6480 890
rect 7400 880 7440 890
rect 7960 880 8000 890
rect 8120 880 8160 890
rect 8200 880 8440 890
rect 8640 880 8880 890
rect 9080 880 9160 890
rect 9440 880 9480 890
rect 760 870 920 880
rect 1360 870 1440 880
rect 2000 870 2040 880
rect 2680 870 2720 880
rect 5320 870 5360 880
rect 5400 870 5680 880
rect 5800 870 6040 880
rect 6200 870 6280 880
rect 6400 870 6480 880
rect 7400 870 7440 880
rect 7960 870 8000 880
rect 8120 870 8160 880
rect 8200 870 8440 880
rect 8640 870 8880 880
rect 9080 870 9160 880
rect 9440 870 9480 880
rect 760 860 920 870
rect 1360 860 1440 870
rect 2000 860 2040 870
rect 2680 860 2720 870
rect 5320 860 5360 870
rect 5400 860 5680 870
rect 5800 860 6040 870
rect 6200 860 6280 870
rect 6400 860 6480 870
rect 7400 860 7440 870
rect 7960 860 8000 870
rect 8120 860 8160 870
rect 8200 860 8440 870
rect 8640 860 8880 870
rect 9080 860 9160 870
rect 9440 860 9480 870
rect 640 850 680 860
rect 760 850 920 860
rect 1320 850 1400 860
rect 2640 850 2680 860
rect 5360 850 5440 860
rect 5760 850 6040 860
rect 6200 850 6280 860
rect 6440 850 6480 860
rect 7360 850 7440 860
rect 7960 850 8000 860
rect 8120 850 8160 860
rect 8200 850 8480 860
rect 8640 850 8840 860
rect 9080 850 9160 860
rect 9400 850 9440 860
rect 640 840 680 850
rect 760 840 920 850
rect 1320 840 1400 850
rect 2640 840 2680 850
rect 5360 840 5440 850
rect 5760 840 6040 850
rect 6200 840 6280 850
rect 6440 840 6480 850
rect 7360 840 7440 850
rect 7960 840 8000 850
rect 8120 840 8160 850
rect 8200 840 8480 850
rect 8640 840 8840 850
rect 9080 840 9160 850
rect 9400 840 9440 850
rect 640 830 680 840
rect 760 830 920 840
rect 1320 830 1400 840
rect 2640 830 2680 840
rect 5360 830 5440 840
rect 5760 830 6040 840
rect 6200 830 6280 840
rect 6440 830 6480 840
rect 7360 830 7440 840
rect 7960 830 8000 840
rect 8120 830 8160 840
rect 8200 830 8480 840
rect 8640 830 8840 840
rect 9080 830 9160 840
rect 9400 830 9440 840
rect 640 820 680 830
rect 760 820 920 830
rect 1320 820 1400 830
rect 2640 820 2680 830
rect 5360 820 5440 830
rect 5760 820 6040 830
rect 6200 820 6280 830
rect 6440 820 6480 830
rect 7360 820 7440 830
rect 7960 820 8000 830
rect 8120 820 8160 830
rect 8200 820 8480 830
rect 8640 820 8840 830
rect 9080 820 9160 830
rect 9400 820 9440 830
rect 640 810 680 820
rect 760 810 840 820
rect 1160 810 1200 820
rect 1280 810 1360 820
rect 2560 810 2600 820
rect 3920 810 4000 820
rect 5480 810 5520 820
rect 5760 810 6040 820
rect 6160 810 6280 820
rect 6440 810 6520 820
rect 7360 810 7400 820
rect 7960 810 8000 820
rect 8120 810 8160 820
rect 8240 810 8840 820
rect 9160 810 9200 820
rect 9400 810 9440 820
rect 640 800 680 810
rect 760 800 840 810
rect 1160 800 1200 810
rect 1280 800 1360 810
rect 2560 800 2600 810
rect 3920 800 4000 810
rect 5480 800 5520 810
rect 5760 800 6040 810
rect 6160 800 6280 810
rect 6440 800 6520 810
rect 7360 800 7400 810
rect 7960 800 8000 810
rect 8120 800 8160 810
rect 8240 800 8840 810
rect 9160 800 9200 810
rect 9400 800 9440 810
rect 640 790 680 800
rect 760 790 840 800
rect 1160 790 1200 800
rect 1280 790 1360 800
rect 2560 790 2600 800
rect 3920 790 4000 800
rect 5480 790 5520 800
rect 5760 790 6040 800
rect 6160 790 6280 800
rect 6440 790 6520 800
rect 7360 790 7400 800
rect 7960 790 8000 800
rect 8120 790 8160 800
rect 8240 790 8840 800
rect 9160 790 9200 800
rect 9400 790 9440 800
rect 640 780 680 790
rect 760 780 840 790
rect 1160 780 1200 790
rect 1280 780 1360 790
rect 2560 780 2600 790
rect 3920 780 4000 790
rect 5480 780 5520 790
rect 5760 780 6040 790
rect 6160 780 6280 790
rect 6440 780 6520 790
rect 7360 780 7400 790
rect 7960 780 8000 790
rect 8120 780 8160 790
rect 8240 780 8840 790
rect 9160 780 9200 790
rect 9400 780 9440 790
rect 720 770 800 780
rect 1120 770 1160 780
rect 1240 770 1280 780
rect 2040 770 2080 780
rect 3520 770 3560 780
rect 3880 770 3920 780
rect 5760 770 6280 780
rect 6480 770 6520 780
rect 7360 770 7400 780
rect 7960 770 8000 780
rect 8120 770 8160 780
rect 8240 770 8800 780
rect 9160 770 9200 780
rect 9360 770 9400 780
rect 720 760 800 770
rect 1120 760 1160 770
rect 1240 760 1280 770
rect 2040 760 2080 770
rect 3520 760 3560 770
rect 3880 760 3920 770
rect 5760 760 6280 770
rect 6480 760 6520 770
rect 7360 760 7400 770
rect 7960 760 8000 770
rect 8120 760 8160 770
rect 8240 760 8800 770
rect 9160 760 9200 770
rect 9360 760 9400 770
rect 720 750 800 760
rect 1120 750 1160 760
rect 1240 750 1280 760
rect 2040 750 2080 760
rect 3520 750 3560 760
rect 3880 750 3920 760
rect 5760 750 6280 760
rect 6480 750 6520 760
rect 7360 750 7400 760
rect 7960 750 8000 760
rect 8120 750 8160 760
rect 8240 750 8800 760
rect 9160 750 9200 760
rect 9360 750 9400 760
rect 720 740 800 750
rect 1120 740 1160 750
rect 1240 740 1280 750
rect 2040 740 2080 750
rect 3520 740 3560 750
rect 3880 740 3920 750
rect 5760 740 6280 750
rect 6480 740 6520 750
rect 7360 740 7400 750
rect 7960 740 8000 750
rect 8120 740 8160 750
rect 8240 740 8800 750
rect 9160 740 9200 750
rect 9360 740 9400 750
rect 600 730 640 740
rect 720 730 760 740
rect 1200 730 1280 740
rect 3360 730 3400 740
rect 3920 730 3960 740
rect 4000 730 4040 740
rect 5760 730 6280 740
rect 6480 730 6560 740
rect 6840 730 6880 740
rect 7360 730 7400 740
rect 8120 730 8160 740
rect 8240 730 8760 740
rect 9160 730 9200 740
rect 600 720 640 730
rect 720 720 760 730
rect 1200 720 1280 730
rect 3360 720 3400 730
rect 3920 720 3960 730
rect 4000 720 4040 730
rect 5760 720 6280 730
rect 6480 720 6560 730
rect 6840 720 6880 730
rect 7360 720 7400 730
rect 8120 720 8160 730
rect 8240 720 8760 730
rect 9160 720 9200 730
rect 600 710 640 720
rect 720 710 760 720
rect 1200 710 1280 720
rect 3360 710 3400 720
rect 3920 710 3960 720
rect 4000 710 4040 720
rect 5760 710 6280 720
rect 6480 710 6560 720
rect 6840 710 6880 720
rect 7360 710 7400 720
rect 8120 710 8160 720
rect 8240 710 8760 720
rect 9160 710 9200 720
rect 600 700 640 710
rect 720 700 760 710
rect 1200 700 1280 710
rect 3360 700 3400 710
rect 3920 700 3960 710
rect 4000 700 4040 710
rect 5760 700 6280 710
rect 6480 700 6560 710
rect 6840 700 6880 710
rect 7360 700 7400 710
rect 8120 700 8160 710
rect 8240 700 8760 710
rect 9160 700 9200 710
rect 600 690 640 700
rect 680 690 760 700
rect 1000 690 1040 700
rect 1200 690 1320 700
rect 2080 690 2120 700
rect 2360 690 2400 700
rect 4120 690 4160 700
rect 4760 690 4800 700
rect 5520 690 5640 700
rect 5760 690 6280 700
rect 6520 690 6560 700
rect 7360 690 7400 700
rect 8000 690 8040 700
rect 8120 690 8160 700
rect 8280 690 8760 700
rect 9160 690 9200 700
rect 9320 690 9360 700
rect 600 680 640 690
rect 680 680 760 690
rect 1000 680 1040 690
rect 1200 680 1320 690
rect 2080 680 2120 690
rect 2360 680 2400 690
rect 4120 680 4160 690
rect 4760 680 4800 690
rect 5520 680 5640 690
rect 5760 680 6280 690
rect 6520 680 6560 690
rect 7360 680 7400 690
rect 8000 680 8040 690
rect 8120 680 8160 690
rect 8280 680 8760 690
rect 9160 680 9200 690
rect 9320 680 9360 690
rect 600 670 640 680
rect 680 670 760 680
rect 1000 670 1040 680
rect 1200 670 1320 680
rect 2080 670 2120 680
rect 2360 670 2400 680
rect 4120 670 4160 680
rect 4760 670 4800 680
rect 5520 670 5640 680
rect 5760 670 6280 680
rect 6520 670 6560 680
rect 7360 670 7400 680
rect 8000 670 8040 680
rect 8120 670 8160 680
rect 8280 670 8760 680
rect 9160 670 9200 680
rect 9320 670 9360 680
rect 600 660 640 670
rect 680 660 760 670
rect 1000 660 1040 670
rect 1200 660 1320 670
rect 2080 660 2120 670
rect 2360 660 2400 670
rect 4120 660 4160 670
rect 4760 660 4800 670
rect 5520 660 5640 670
rect 5760 660 6280 670
rect 6520 660 6560 670
rect 7360 660 7400 670
rect 8000 660 8040 670
rect 8120 660 8160 670
rect 8280 660 8760 670
rect 9160 660 9200 670
rect 9320 660 9360 670
rect 480 650 720 660
rect 760 650 1000 660
rect 1160 650 1280 660
rect 2280 650 2320 660
rect 3240 650 3280 660
rect 4920 650 4960 660
rect 5560 650 5680 660
rect 5760 650 6280 660
rect 6520 650 6600 660
rect 7320 650 7400 660
rect 8000 650 8040 660
rect 8120 650 8160 660
rect 8320 650 8720 660
rect 9120 650 9160 660
rect 480 640 720 650
rect 760 640 1000 650
rect 1160 640 1280 650
rect 2280 640 2320 650
rect 3240 640 3280 650
rect 4920 640 4960 650
rect 5560 640 5680 650
rect 5760 640 6280 650
rect 6520 640 6600 650
rect 7320 640 7400 650
rect 8000 640 8040 650
rect 8120 640 8160 650
rect 8320 640 8720 650
rect 9120 640 9160 650
rect 480 630 720 640
rect 760 630 1000 640
rect 1160 630 1280 640
rect 2280 630 2320 640
rect 3240 630 3280 640
rect 4920 630 4960 640
rect 5560 630 5680 640
rect 5760 630 6280 640
rect 6520 630 6600 640
rect 7320 630 7400 640
rect 8000 630 8040 640
rect 8120 630 8160 640
rect 8320 630 8720 640
rect 9120 630 9160 640
rect 480 620 720 630
rect 760 620 1000 630
rect 1160 620 1280 630
rect 2280 620 2320 630
rect 3240 620 3280 630
rect 4920 620 4960 630
rect 5560 620 5680 630
rect 5760 620 6280 630
rect 6520 620 6600 630
rect 7320 620 7400 630
rect 8000 620 8040 630
rect 8120 620 8160 630
rect 8320 620 8720 630
rect 9120 620 9160 630
rect 360 610 440 620
rect 640 610 720 620
rect 760 610 920 620
rect 1080 610 1240 620
rect 1320 610 1440 620
rect 2120 610 2160 620
rect 2200 610 2240 620
rect 5600 610 5680 620
rect 5840 610 6320 620
rect 6560 610 6600 620
rect 6880 610 6920 620
rect 7320 610 7400 620
rect 8040 610 8160 620
rect 8360 610 8680 620
rect 9080 610 9160 620
rect 9280 610 9320 620
rect 360 600 440 610
rect 640 600 720 610
rect 760 600 920 610
rect 1080 600 1240 610
rect 1320 600 1440 610
rect 2120 600 2160 610
rect 2200 600 2240 610
rect 5600 600 5680 610
rect 5840 600 6320 610
rect 6560 600 6600 610
rect 6880 600 6920 610
rect 7320 600 7400 610
rect 8040 600 8160 610
rect 8360 600 8680 610
rect 9080 600 9160 610
rect 9280 600 9320 610
rect 360 590 440 600
rect 640 590 720 600
rect 760 590 920 600
rect 1080 590 1240 600
rect 1320 590 1440 600
rect 2120 590 2160 600
rect 2200 590 2240 600
rect 5600 590 5680 600
rect 5840 590 6320 600
rect 6560 590 6600 600
rect 6880 590 6920 600
rect 7320 590 7400 600
rect 8040 590 8160 600
rect 8360 590 8680 600
rect 9080 590 9160 600
rect 9280 590 9320 600
rect 360 580 440 590
rect 640 580 720 590
rect 760 580 920 590
rect 1080 580 1240 590
rect 1320 580 1440 590
rect 2120 580 2160 590
rect 2200 580 2240 590
rect 5600 580 5680 590
rect 5840 580 6320 590
rect 6560 580 6600 590
rect 6880 580 6920 590
rect 7320 580 7400 590
rect 8040 580 8160 590
rect 8360 580 8680 590
rect 9080 580 9160 590
rect 9280 580 9320 590
rect 320 570 360 580
rect 640 570 920 580
rect 1040 570 1200 580
rect 1240 570 1280 580
rect 1440 570 1480 580
rect 4480 570 4560 580
rect 4680 570 4720 580
rect 5600 570 5680 580
rect 5880 570 6320 580
rect 6560 570 6640 580
rect 6880 570 6920 580
rect 7320 570 7360 580
rect 8080 570 8120 580
rect 8440 570 8560 580
rect 9040 570 9200 580
rect 9240 570 9280 580
rect 320 560 360 570
rect 640 560 920 570
rect 1040 560 1200 570
rect 1240 560 1280 570
rect 1440 560 1480 570
rect 4480 560 4560 570
rect 4680 560 4720 570
rect 5600 560 5680 570
rect 5880 560 6320 570
rect 6560 560 6640 570
rect 6880 560 6920 570
rect 7320 560 7360 570
rect 8080 560 8120 570
rect 8440 560 8560 570
rect 9040 560 9200 570
rect 9240 560 9280 570
rect 320 550 360 560
rect 640 550 920 560
rect 1040 550 1200 560
rect 1240 550 1280 560
rect 1440 550 1480 560
rect 4480 550 4560 560
rect 4680 550 4720 560
rect 5600 550 5680 560
rect 5880 550 6320 560
rect 6560 550 6640 560
rect 6880 550 6920 560
rect 7320 550 7360 560
rect 8080 550 8120 560
rect 8440 550 8560 560
rect 9040 550 9200 560
rect 9240 550 9280 560
rect 320 540 360 550
rect 640 540 920 550
rect 1040 540 1200 550
rect 1240 540 1280 550
rect 1440 540 1480 550
rect 4480 540 4560 550
rect 4680 540 4720 550
rect 5600 540 5680 550
rect 5880 540 6320 550
rect 6560 540 6640 550
rect 6880 540 6920 550
rect 7320 540 7360 550
rect 8080 540 8120 550
rect 8440 540 8560 550
rect 9040 540 9200 550
rect 9240 540 9280 550
rect 200 530 360 540
rect 640 530 680 540
rect 720 530 760 540
rect 800 530 840 540
rect 880 530 960 540
rect 1040 530 1080 540
rect 1200 530 1240 540
rect 1480 530 1520 540
rect 2920 530 2960 540
rect 4360 530 4480 540
rect 4520 530 4560 540
rect 4640 530 4680 540
rect 4720 530 4760 540
rect 5920 530 6320 540
rect 6600 530 6640 540
rect 7280 530 7360 540
rect 9160 530 9200 540
rect 9240 530 9280 540
rect 200 520 360 530
rect 640 520 680 530
rect 720 520 760 530
rect 800 520 840 530
rect 880 520 960 530
rect 1040 520 1080 530
rect 1200 520 1240 530
rect 1480 520 1520 530
rect 2920 520 2960 530
rect 4360 520 4480 530
rect 4520 520 4560 530
rect 4640 520 4680 530
rect 4720 520 4760 530
rect 5920 520 6320 530
rect 6600 520 6640 530
rect 7280 520 7360 530
rect 9160 520 9200 530
rect 9240 520 9280 530
rect 200 510 360 520
rect 640 510 680 520
rect 720 510 760 520
rect 800 510 840 520
rect 880 510 960 520
rect 1040 510 1080 520
rect 1200 510 1240 520
rect 1480 510 1520 520
rect 2920 510 2960 520
rect 4360 510 4480 520
rect 4520 510 4560 520
rect 4640 510 4680 520
rect 4720 510 4760 520
rect 5920 510 6320 520
rect 6600 510 6640 520
rect 7280 510 7360 520
rect 9160 510 9200 520
rect 9240 510 9280 520
rect 200 500 360 510
rect 640 500 680 510
rect 720 500 760 510
rect 800 500 840 510
rect 880 500 960 510
rect 1040 500 1080 510
rect 1200 500 1240 510
rect 1480 500 1520 510
rect 2920 500 2960 510
rect 4360 500 4480 510
rect 4520 500 4560 510
rect 4640 500 4680 510
rect 4720 500 4760 510
rect 5920 500 6320 510
rect 6600 500 6640 510
rect 7280 500 7360 510
rect 9160 500 9200 510
rect 9240 500 9280 510
rect 120 490 160 500
rect 320 490 360 500
rect 520 490 640 500
rect 920 490 1080 500
rect 1520 490 1560 500
rect 4240 490 4320 500
rect 4560 490 4680 500
rect 4720 490 4760 500
rect 5800 490 5840 500
rect 5920 490 6320 500
rect 6600 490 6680 500
rect 7280 490 7360 500
rect 9080 490 9160 500
rect 120 480 160 490
rect 320 480 360 490
rect 520 480 640 490
rect 920 480 1080 490
rect 1520 480 1560 490
rect 4240 480 4320 490
rect 4560 480 4680 490
rect 4720 480 4760 490
rect 5800 480 5840 490
rect 5920 480 6320 490
rect 6600 480 6680 490
rect 7280 480 7360 490
rect 9080 480 9160 490
rect 120 470 160 480
rect 320 470 360 480
rect 520 470 640 480
rect 920 470 1080 480
rect 1520 470 1560 480
rect 4240 470 4320 480
rect 4560 470 4680 480
rect 4720 470 4760 480
rect 5800 470 5840 480
rect 5920 470 6320 480
rect 6600 470 6680 480
rect 7280 470 7360 480
rect 9080 470 9160 480
rect 120 460 160 470
rect 320 460 360 470
rect 520 460 640 470
rect 920 460 1080 470
rect 1520 460 1560 470
rect 4240 460 4320 470
rect 4560 460 4680 470
rect 4720 460 4760 470
rect 5800 460 5840 470
rect 5920 460 6320 470
rect 6600 460 6680 470
rect 7280 460 7360 470
rect 9080 460 9160 470
rect 80 450 120 460
rect 360 450 440 460
rect 480 450 560 460
rect 600 450 680 460
rect 1560 450 1720 460
rect 1840 450 1960 460
rect 2280 450 2320 460
rect 2560 450 2640 460
rect 4200 450 4280 460
rect 4560 450 4680 460
rect 4720 450 4760 460
rect 4960 450 5000 460
rect 5800 450 5880 460
rect 5960 450 6280 460
rect 6640 450 6720 460
rect 7240 450 7360 460
rect 9000 450 9120 460
rect 9160 450 9200 460
rect 80 440 120 450
rect 360 440 440 450
rect 480 440 560 450
rect 600 440 680 450
rect 1560 440 1720 450
rect 1840 440 1960 450
rect 2280 440 2320 450
rect 2560 440 2640 450
rect 4200 440 4280 450
rect 4560 440 4680 450
rect 4720 440 4760 450
rect 4960 440 5000 450
rect 5800 440 5880 450
rect 5960 440 6280 450
rect 6640 440 6720 450
rect 7240 440 7360 450
rect 9000 440 9120 450
rect 9160 440 9200 450
rect 80 430 120 440
rect 360 430 440 440
rect 480 430 560 440
rect 600 430 680 440
rect 1560 430 1720 440
rect 1840 430 1960 440
rect 2280 430 2320 440
rect 2560 430 2640 440
rect 4200 430 4280 440
rect 4560 430 4680 440
rect 4720 430 4760 440
rect 4960 430 5000 440
rect 5800 430 5880 440
rect 5960 430 6280 440
rect 6640 430 6720 440
rect 7240 430 7360 440
rect 9000 430 9120 440
rect 9160 430 9200 440
rect 80 420 120 430
rect 360 420 440 430
rect 480 420 560 430
rect 600 420 680 430
rect 1560 420 1720 430
rect 1840 420 1960 430
rect 2280 420 2320 430
rect 2560 420 2640 430
rect 4200 420 4280 430
rect 4560 420 4680 430
rect 4720 420 4760 430
rect 4960 420 5000 430
rect 5800 420 5880 430
rect 5960 420 6280 430
rect 6640 420 6720 430
rect 7240 420 7360 430
rect 9000 420 9120 430
rect 9160 420 9200 430
rect 480 410 680 420
rect 4200 410 4280 420
rect 4320 410 4360 420
rect 4960 410 5000 420
rect 6000 410 6280 420
rect 6680 410 6720 420
rect 7240 410 7360 420
rect 9000 410 9120 420
rect 9320 410 9360 420
rect 480 400 680 410
rect 4200 400 4280 410
rect 4320 400 4360 410
rect 4960 400 5000 410
rect 6000 400 6280 410
rect 6680 400 6720 410
rect 7240 400 7360 410
rect 9000 400 9120 410
rect 9320 400 9360 410
rect 480 390 680 400
rect 4200 390 4280 400
rect 4320 390 4360 400
rect 4960 390 5000 400
rect 6000 390 6280 400
rect 6680 390 6720 400
rect 7240 390 7360 400
rect 9000 390 9120 400
rect 9320 390 9360 400
rect 480 380 680 390
rect 4200 380 4280 390
rect 4320 380 4360 390
rect 4960 380 5000 390
rect 6000 380 6280 390
rect 6680 380 6720 390
rect 7240 380 7360 390
rect 9000 380 9120 390
rect 9320 380 9360 390
rect 440 370 680 380
rect 1040 370 1080 380
rect 4200 370 4320 380
rect 4360 370 4400 380
rect 4560 370 4600 380
rect 4960 370 5000 380
rect 5800 370 5840 380
rect 6000 370 6280 380
rect 6720 370 6760 380
rect 7200 370 7320 380
rect 8800 370 8840 380
rect 8960 370 9040 380
rect 9080 370 9160 380
rect 9240 370 9320 380
rect 9360 370 9400 380
rect 440 360 680 370
rect 1040 360 1080 370
rect 4200 360 4320 370
rect 4360 360 4400 370
rect 4560 360 4600 370
rect 4960 360 5000 370
rect 5800 360 5840 370
rect 6000 360 6280 370
rect 6720 360 6760 370
rect 7200 360 7320 370
rect 8800 360 8840 370
rect 8960 360 9040 370
rect 9080 360 9160 370
rect 9240 360 9320 370
rect 9360 360 9400 370
rect 440 350 680 360
rect 1040 350 1080 360
rect 4200 350 4320 360
rect 4360 350 4400 360
rect 4560 350 4600 360
rect 4960 350 5000 360
rect 5800 350 5840 360
rect 6000 350 6280 360
rect 6720 350 6760 360
rect 7200 350 7320 360
rect 8800 350 8840 360
rect 8960 350 9040 360
rect 9080 350 9160 360
rect 9240 350 9320 360
rect 9360 350 9400 360
rect 440 340 680 350
rect 1040 340 1080 350
rect 4200 340 4320 350
rect 4360 340 4400 350
rect 4560 340 4600 350
rect 4960 340 5000 350
rect 5800 340 5840 350
rect 6000 340 6280 350
rect 6720 340 6760 350
rect 7200 340 7320 350
rect 8800 340 8840 350
rect 8960 340 9040 350
rect 9080 340 9160 350
rect 9240 340 9320 350
rect 9360 340 9400 350
rect 0 330 40 340
rect 400 330 480 340
rect 720 330 800 340
rect 4200 330 4240 340
rect 4400 330 4560 340
rect 4680 330 4760 340
rect 4960 330 5000 340
rect 6000 330 6280 340
rect 6760 330 6840 340
rect 7160 330 7320 340
rect 9040 330 9080 340
rect 9120 330 9160 340
rect 9360 330 9400 340
rect 0 320 40 330
rect 400 320 480 330
rect 720 320 800 330
rect 4200 320 4240 330
rect 4400 320 4560 330
rect 4680 320 4760 330
rect 4960 320 5000 330
rect 6000 320 6280 330
rect 6760 320 6840 330
rect 7160 320 7320 330
rect 9040 320 9080 330
rect 9120 320 9160 330
rect 9360 320 9400 330
rect 0 310 40 320
rect 400 310 480 320
rect 720 310 800 320
rect 4200 310 4240 320
rect 4400 310 4560 320
rect 4680 310 4760 320
rect 4960 310 5000 320
rect 6000 310 6280 320
rect 6760 310 6840 320
rect 7160 310 7320 320
rect 9040 310 9080 320
rect 9120 310 9160 320
rect 9360 310 9400 320
rect 0 300 40 310
rect 400 300 480 310
rect 720 300 800 310
rect 4200 300 4240 310
rect 4400 300 4560 310
rect 4680 300 4760 310
rect 4960 300 5000 310
rect 6000 300 6280 310
rect 6760 300 6840 310
rect 7160 300 7320 310
rect 9040 300 9080 310
rect 9120 300 9160 310
rect 9360 300 9400 310
rect 0 290 40 300
rect 400 290 440 300
rect 640 290 680 300
rect 840 290 1040 300
rect 4120 290 4200 300
rect 4520 290 4680 300
rect 6000 290 6040 300
rect 6120 290 6280 300
rect 6800 290 6920 300
rect 7040 290 7320 300
rect 8880 290 8920 300
rect 9080 290 9120 300
rect 9200 290 9240 300
rect 9280 290 9400 300
rect 0 280 40 290
rect 400 280 440 290
rect 640 280 680 290
rect 840 280 1040 290
rect 4120 280 4200 290
rect 4520 280 4680 290
rect 6000 280 6040 290
rect 6120 280 6280 290
rect 6800 280 6920 290
rect 7040 280 7320 290
rect 8880 280 8920 290
rect 9080 280 9120 290
rect 9200 280 9240 290
rect 9280 280 9400 290
rect 0 270 40 280
rect 400 270 440 280
rect 640 270 680 280
rect 840 270 1040 280
rect 4120 270 4200 280
rect 4520 270 4680 280
rect 6000 270 6040 280
rect 6120 270 6280 280
rect 6800 270 6920 280
rect 7040 270 7320 280
rect 8880 270 8920 280
rect 9080 270 9120 280
rect 9200 270 9240 280
rect 9280 270 9400 280
rect 0 260 40 270
rect 400 260 440 270
rect 640 260 680 270
rect 840 260 1040 270
rect 4120 260 4200 270
rect 4520 260 4680 270
rect 6000 260 6040 270
rect 6120 260 6280 270
rect 6800 260 6920 270
rect 7040 260 7320 270
rect 8880 260 8920 270
rect 9080 260 9120 270
rect 9200 260 9240 270
rect 9280 260 9400 270
rect 120 250 200 260
rect 400 250 440 260
rect 640 250 680 260
rect 880 250 1000 260
rect 4120 250 4160 260
rect 4560 250 4640 260
rect 6120 250 6280 260
rect 6840 250 7320 260
rect 9000 250 9040 260
rect 9080 250 9120 260
rect 9200 250 9320 260
rect 120 240 200 250
rect 400 240 440 250
rect 640 240 680 250
rect 880 240 1000 250
rect 4120 240 4160 250
rect 4560 240 4640 250
rect 6120 240 6280 250
rect 6840 240 7320 250
rect 9000 240 9040 250
rect 9080 240 9120 250
rect 9200 240 9320 250
rect 120 230 200 240
rect 400 230 440 240
rect 640 230 680 240
rect 880 230 1000 240
rect 4120 230 4160 240
rect 4560 230 4640 240
rect 6120 230 6280 240
rect 6840 230 7320 240
rect 9000 230 9040 240
rect 9080 230 9120 240
rect 9200 230 9320 240
rect 120 220 200 230
rect 400 220 440 230
rect 640 220 680 230
rect 880 220 1000 230
rect 4120 220 4160 230
rect 4560 220 4640 230
rect 6120 220 6280 230
rect 6840 220 7320 230
rect 9000 220 9040 230
rect 9080 220 9120 230
rect 9200 220 9320 230
rect 80 210 160 220
rect 200 210 240 220
rect 360 210 440 220
rect 600 210 680 220
rect 880 210 1000 220
rect 4160 210 4240 220
rect 4320 210 4400 220
rect 4560 210 4600 220
rect 6080 210 6320 220
rect 6880 210 7320 220
rect 8600 210 8640 220
rect 8680 210 8720 220
rect 8840 210 8880 220
rect 8920 210 8960 220
rect 9040 210 9080 220
rect 9160 210 9280 220
rect 9800 210 9840 220
rect 80 200 160 210
rect 200 200 240 210
rect 360 200 440 210
rect 600 200 680 210
rect 880 200 1000 210
rect 4160 200 4240 210
rect 4320 200 4400 210
rect 4560 200 4600 210
rect 6080 200 6320 210
rect 6880 200 7320 210
rect 8600 200 8640 210
rect 8680 200 8720 210
rect 8840 200 8880 210
rect 8920 200 8960 210
rect 9040 200 9080 210
rect 9160 200 9280 210
rect 9800 200 9840 210
rect 80 190 160 200
rect 200 190 240 200
rect 360 190 440 200
rect 600 190 680 200
rect 880 190 1000 200
rect 4160 190 4240 200
rect 4320 190 4400 200
rect 4560 190 4600 200
rect 6080 190 6320 200
rect 6880 190 7320 200
rect 8600 190 8640 200
rect 8680 190 8720 200
rect 8840 190 8880 200
rect 8920 190 8960 200
rect 9040 190 9080 200
rect 9160 190 9280 200
rect 9800 190 9840 200
rect 80 180 160 190
rect 200 180 240 190
rect 360 180 440 190
rect 600 180 680 190
rect 880 180 1000 190
rect 4160 180 4240 190
rect 4320 180 4400 190
rect 4560 180 4600 190
rect 6080 180 6320 190
rect 6880 180 7320 190
rect 8600 180 8640 190
rect 8680 180 8720 190
rect 8840 180 8880 190
rect 8920 180 8960 190
rect 9040 180 9080 190
rect 9160 180 9280 190
rect 9800 180 9840 190
rect 120 170 160 180
rect 280 170 360 180
rect 440 170 720 180
rect 800 170 1000 180
rect 4200 170 4560 180
rect 4840 170 4920 180
rect 5000 170 5040 180
rect 6080 170 6320 180
rect 6960 170 7320 180
rect 8560 170 8760 180
rect 8880 170 8920 180
rect 9160 170 9200 180
rect 9280 170 9320 180
rect 9760 170 9800 180
rect 9840 170 9990 180
rect 120 160 160 170
rect 280 160 360 170
rect 440 160 720 170
rect 800 160 1000 170
rect 4200 160 4560 170
rect 4840 160 4920 170
rect 5000 160 5040 170
rect 6080 160 6320 170
rect 6960 160 7320 170
rect 8560 160 8760 170
rect 8880 160 8920 170
rect 9160 160 9200 170
rect 9280 160 9320 170
rect 9760 160 9800 170
rect 9840 160 9990 170
rect 120 150 160 160
rect 280 150 360 160
rect 440 150 720 160
rect 800 150 1000 160
rect 4200 150 4560 160
rect 4840 150 4920 160
rect 5000 150 5040 160
rect 6080 150 6320 160
rect 6960 150 7320 160
rect 8560 150 8760 160
rect 8880 150 8920 160
rect 9160 150 9200 160
rect 9280 150 9320 160
rect 9760 150 9800 160
rect 9840 150 9990 160
rect 120 140 160 150
rect 280 140 360 150
rect 440 140 720 150
rect 800 140 1000 150
rect 4200 140 4560 150
rect 4840 140 4920 150
rect 5000 140 5040 150
rect 6080 140 6320 150
rect 6960 140 7320 150
rect 8560 140 8760 150
rect 8880 140 8920 150
rect 9160 140 9200 150
rect 9280 140 9320 150
rect 9760 140 9800 150
rect 9840 140 9990 150
rect 120 130 160 140
rect 240 130 320 140
rect 560 130 1000 140
rect 4240 130 4280 140
rect 4440 130 4560 140
rect 4600 130 4640 140
rect 4680 130 4720 140
rect 4800 130 4880 140
rect 4920 130 4960 140
rect 5960 130 6000 140
rect 6080 130 6320 140
rect 7000 130 7320 140
rect 8560 130 8720 140
rect 8800 130 8840 140
rect 8920 130 8960 140
rect 9160 130 9200 140
rect 9320 130 9360 140
rect 9720 130 9760 140
rect 9880 130 9990 140
rect 120 120 160 130
rect 240 120 320 130
rect 560 120 1000 130
rect 4240 120 4280 130
rect 4440 120 4560 130
rect 4600 120 4640 130
rect 4680 120 4720 130
rect 4800 120 4880 130
rect 4920 120 4960 130
rect 5960 120 6000 130
rect 6080 120 6320 130
rect 7000 120 7320 130
rect 8560 120 8720 130
rect 8800 120 8840 130
rect 8920 120 8960 130
rect 9160 120 9200 130
rect 9320 120 9360 130
rect 9720 120 9760 130
rect 9880 120 9990 130
rect 120 110 160 120
rect 240 110 320 120
rect 560 110 1000 120
rect 4240 110 4280 120
rect 4440 110 4560 120
rect 4600 110 4640 120
rect 4680 110 4720 120
rect 4800 110 4880 120
rect 4920 110 4960 120
rect 5960 110 6000 120
rect 6080 110 6320 120
rect 7000 110 7320 120
rect 8560 110 8720 120
rect 8800 110 8840 120
rect 8920 110 8960 120
rect 9160 110 9200 120
rect 9320 110 9360 120
rect 9720 110 9760 120
rect 9880 110 9990 120
rect 120 100 160 110
rect 240 100 320 110
rect 560 100 1000 110
rect 4240 100 4280 110
rect 4440 100 4560 110
rect 4600 100 4640 110
rect 4680 100 4720 110
rect 4800 100 4880 110
rect 4920 100 4960 110
rect 5960 100 6000 110
rect 6080 100 6320 110
rect 7000 100 7320 110
rect 8560 100 8720 110
rect 8800 100 8840 110
rect 8920 100 8960 110
rect 9160 100 9200 110
rect 9320 100 9360 110
rect 9720 100 9760 110
rect 9880 100 9990 110
rect 120 90 160 100
rect 280 90 320 100
rect 640 90 680 100
rect 840 90 1000 100
rect 4280 90 4320 100
rect 4520 90 4840 100
rect 4880 90 4920 100
rect 5880 90 6000 100
rect 6080 90 6400 100
rect 7040 90 7320 100
rect 8600 90 8720 100
rect 9000 90 9080 100
rect 9160 90 9200 100
rect 9360 90 9440 100
rect 9760 90 9800 100
rect 9880 90 9920 100
rect 9960 90 9990 100
rect 120 80 160 90
rect 280 80 320 90
rect 640 80 680 90
rect 840 80 1000 90
rect 4280 80 4320 90
rect 4520 80 4840 90
rect 4880 80 4920 90
rect 5880 80 6000 90
rect 6080 80 6400 90
rect 7040 80 7320 90
rect 8600 80 8720 90
rect 9000 80 9080 90
rect 9160 80 9200 90
rect 9360 80 9440 90
rect 9760 80 9800 90
rect 9880 80 9920 90
rect 9960 80 9990 90
rect 120 70 160 80
rect 280 70 320 80
rect 640 70 680 80
rect 840 70 1000 80
rect 4280 70 4320 80
rect 4520 70 4840 80
rect 4880 70 4920 80
rect 5880 70 6000 80
rect 6080 70 6400 80
rect 7040 70 7320 80
rect 8600 70 8720 80
rect 9000 70 9080 80
rect 9160 70 9200 80
rect 9360 70 9440 80
rect 9760 70 9800 80
rect 9880 70 9920 80
rect 9960 70 9990 80
rect 120 60 160 70
rect 280 60 320 70
rect 640 60 680 70
rect 840 60 1000 70
rect 4280 60 4320 70
rect 4520 60 4840 70
rect 4880 60 4920 70
rect 5880 60 6000 70
rect 6080 60 6400 70
rect 7040 60 7320 70
rect 8600 60 8720 70
rect 9000 60 9080 70
rect 9160 60 9200 70
rect 9360 60 9440 70
rect 9760 60 9800 70
rect 9880 60 9920 70
rect 9960 60 9990 70
rect 120 50 160 60
rect 280 50 320 60
rect 880 50 1000 60
rect 4520 50 4560 60
rect 4600 50 4800 60
rect 4840 50 4920 60
rect 5040 50 5080 60
rect 6080 50 6440 60
rect 7120 50 7320 60
rect 8720 50 8760 60
rect 8920 50 8960 60
rect 9160 50 9200 60
rect 9440 50 9480 60
rect 9760 50 9800 60
rect 9880 50 9920 60
rect 120 40 160 50
rect 280 40 320 50
rect 880 40 1000 50
rect 4520 40 4560 50
rect 4600 40 4800 50
rect 4840 40 4920 50
rect 5040 40 5080 50
rect 6080 40 6440 50
rect 7120 40 7320 50
rect 8720 40 8760 50
rect 8920 40 8960 50
rect 9160 40 9200 50
rect 9440 40 9480 50
rect 9760 40 9800 50
rect 9880 40 9920 50
rect 120 30 160 40
rect 280 30 320 40
rect 880 30 1000 40
rect 4520 30 4560 40
rect 4600 30 4800 40
rect 4840 30 4920 40
rect 5040 30 5080 40
rect 6080 30 6440 40
rect 7120 30 7320 40
rect 8720 30 8760 40
rect 8920 30 8960 40
rect 9160 30 9200 40
rect 9440 30 9480 40
rect 9760 30 9800 40
rect 9880 30 9920 40
rect 120 20 160 30
rect 280 20 320 30
rect 880 20 1000 30
rect 4520 20 4560 30
rect 4600 20 4800 30
rect 4840 20 4920 30
rect 5040 20 5080 30
rect 6080 20 6440 30
rect 7120 20 7320 30
rect 8720 20 8760 30
rect 8920 20 8960 30
rect 9160 20 9200 30
rect 9440 20 9480 30
rect 9760 20 9800 30
rect 9880 20 9920 30
rect 80 10 160 20
rect 280 10 320 20
rect 680 10 720 20
rect 920 10 1000 20
rect 4360 10 4400 20
rect 4600 10 4920 20
rect 6080 10 6440 20
rect 7160 10 7280 20
rect 8560 10 8600 20
rect 9000 10 9040 20
rect 9440 10 9480 20
rect 80 0 160 10
rect 280 0 320 10
rect 680 0 720 10
rect 920 0 1000 10
rect 4360 0 4400 10
rect 4600 0 4920 10
rect 6080 0 6440 10
rect 7160 0 7280 10
rect 8560 0 8600 10
rect 9000 0 9040 10
rect 9440 0 9480 10
<< metal3 >>
rect 2120 7490 2160 7500
rect 3320 7490 3360 7500
rect 3680 7490 3840 7500
rect 9520 7490 9760 7500
rect 2120 7480 2160 7490
rect 3320 7480 3360 7490
rect 3680 7480 3840 7490
rect 9520 7480 9760 7490
rect 2120 7470 2160 7480
rect 3320 7470 3360 7480
rect 3680 7470 3840 7480
rect 9520 7470 9760 7480
rect 2120 7460 2160 7470
rect 3320 7460 3360 7470
rect 3680 7460 3840 7470
rect 9520 7460 9760 7470
rect 2080 7450 2120 7460
rect 3640 7450 3680 7460
rect 3800 7450 3840 7460
rect 9560 7450 9640 7460
rect 2080 7440 2120 7450
rect 3640 7440 3680 7450
rect 3800 7440 3840 7450
rect 9560 7440 9640 7450
rect 2080 7430 2120 7440
rect 3640 7430 3680 7440
rect 3800 7430 3840 7440
rect 9560 7430 9640 7440
rect 2080 7420 2120 7430
rect 3640 7420 3680 7430
rect 3800 7420 3840 7430
rect 9560 7420 9640 7430
rect 3320 7410 3360 7420
rect 3800 7410 3880 7420
rect 9560 7410 9640 7420
rect 3320 7400 3360 7410
rect 3800 7400 3880 7410
rect 9560 7400 9640 7410
rect 3320 7390 3360 7400
rect 3800 7390 3880 7400
rect 9560 7390 9640 7400
rect 3320 7380 3360 7390
rect 3800 7380 3880 7390
rect 9560 7380 9640 7390
rect 3840 7370 3880 7380
rect 9560 7370 9640 7380
rect 3840 7360 3880 7370
rect 9560 7360 9640 7370
rect 3840 7350 3880 7360
rect 9560 7350 9640 7360
rect 3840 7340 3880 7350
rect 9560 7340 9640 7350
rect 2000 7330 2040 7340
rect 9560 7330 9640 7340
rect 9840 7330 9880 7340
rect 2000 7320 2040 7330
rect 9560 7320 9640 7330
rect 9840 7320 9880 7330
rect 2000 7310 2040 7320
rect 9560 7310 9640 7320
rect 9840 7310 9880 7320
rect 2000 7300 2040 7310
rect 9560 7300 9640 7310
rect 9840 7300 9880 7310
rect 3360 7290 3440 7300
rect 3840 7290 3920 7300
rect 9560 7290 9640 7300
rect 9840 7290 9880 7300
rect 3360 7280 3440 7290
rect 3840 7280 3920 7290
rect 9560 7280 9640 7290
rect 9840 7280 9880 7290
rect 3360 7270 3440 7280
rect 3840 7270 3920 7280
rect 9560 7270 9640 7280
rect 9840 7270 9880 7280
rect 3360 7260 3440 7270
rect 3840 7260 3920 7270
rect 9560 7260 9640 7270
rect 9840 7260 9880 7270
rect 1960 7250 2000 7260
rect 3800 7250 3840 7260
rect 3880 7250 3920 7260
rect 9560 7250 9640 7260
rect 1960 7240 2000 7250
rect 3800 7240 3840 7250
rect 3880 7240 3920 7250
rect 9560 7240 9640 7250
rect 1960 7230 2000 7240
rect 3800 7230 3840 7240
rect 3880 7230 3920 7240
rect 9560 7230 9640 7240
rect 1960 7220 2000 7230
rect 3800 7220 3840 7230
rect 3880 7220 3920 7230
rect 9560 7220 9640 7230
rect 1920 7210 1960 7220
rect 3400 7210 3440 7220
rect 3800 7210 3840 7220
rect 9560 7210 9600 7220
rect 1920 7200 1960 7210
rect 3400 7200 3440 7210
rect 3800 7200 3840 7210
rect 9560 7200 9600 7210
rect 1920 7190 1960 7200
rect 3400 7190 3440 7200
rect 3800 7190 3840 7200
rect 9560 7190 9600 7200
rect 1920 7180 1960 7190
rect 3400 7180 3440 7190
rect 3800 7180 3840 7190
rect 9560 7180 9600 7190
rect 3360 7170 3400 7180
rect 3720 7170 3760 7180
rect 3800 7170 3840 7180
rect 3920 7170 3960 7180
rect 9560 7170 9600 7180
rect 3360 7160 3400 7170
rect 3720 7160 3760 7170
rect 3800 7160 3840 7170
rect 3920 7160 3960 7170
rect 9560 7160 9600 7170
rect 3360 7150 3400 7160
rect 3720 7150 3760 7160
rect 3800 7150 3840 7160
rect 3920 7150 3960 7160
rect 9560 7150 9600 7160
rect 3360 7140 3400 7150
rect 3720 7140 3760 7150
rect 3800 7140 3840 7150
rect 3920 7140 3960 7150
rect 9560 7140 9600 7150
rect 3440 7130 3480 7140
rect 3720 7130 3840 7140
rect 3920 7130 3960 7140
rect 9560 7130 9600 7140
rect 3440 7120 3480 7130
rect 3720 7120 3840 7130
rect 3920 7120 3960 7130
rect 9560 7120 9600 7130
rect 3440 7110 3480 7120
rect 3720 7110 3840 7120
rect 3920 7110 3960 7120
rect 9560 7110 9600 7120
rect 3440 7100 3480 7110
rect 3720 7100 3840 7110
rect 3920 7100 3960 7110
rect 9560 7100 9600 7110
rect 1880 7090 1920 7100
rect 3520 7090 3640 7100
rect 3800 7090 3840 7100
rect 3920 7090 3960 7100
rect 1880 7080 1920 7090
rect 3520 7080 3640 7090
rect 3800 7080 3840 7090
rect 3920 7080 3960 7090
rect 1880 7070 1920 7080
rect 3520 7070 3640 7080
rect 3800 7070 3840 7080
rect 3920 7070 3960 7080
rect 1880 7060 1920 7070
rect 3520 7060 3640 7070
rect 3800 7060 3840 7070
rect 3920 7060 3960 7070
rect 1880 7050 1920 7060
rect 3520 7050 3560 7060
rect 3720 7050 3840 7060
rect 3920 7050 3960 7060
rect 9560 7050 9600 7060
rect 1880 7040 1920 7050
rect 3520 7040 3560 7050
rect 3720 7040 3840 7050
rect 3920 7040 3960 7050
rect 9560 7040 9600 7050
rect 1880 7030 1920 7040
rect 3520 7030 3560 7040
rect 3720 7030 3840 7040
rect 3920 7030 3960 7040
rect 9560 7030 9600 7040
rect 1880 7020 1920 7030
rect 3520 7020 3560 7030
rect 3720 7020 3840 7030
rect 3920 7020 3960 7030
rect 9560 7020 9600 7030
rect 1880 7010 1960 7020
rect 3600 7010 3680 7020
rect 3720 7010 3760 7020
rect 3800 7010 3840 7020
rect 3920 7010 4000 7020
rect 9560 7010 9600 7020
rect 1880 7000 1960 7010
rect 3600 7000 3680 7010
rect 3720 7000 3760 7010
rect 3800 7000 3840 7010
rect 3920 7000 4000 7010
rect 9560 7000 9600 7010
rect 1880 6990 1960 7000
rect 3600 6990 3680 7000
rect 3720 6990 3760 7000
rect 3800 6990 3840 7000
rect 3920 6990 4000 7000
rect 9560 6990 9600 7000
rect 1880 6980 1960 6990
rect 3600 6980 3680 6990
rect 3720 6980 3760 6990
rect 3800 6980 3840 6990
rect 3920 6980 4000 6990
rect 9560 6980 9600 6990
rect 1920 6970 1960 6980
rect 3160 6970 3280 6980
rect 3680 6970 3760 6980
rect 3800 6970 3840 6980
rect 3920 6970 4000 6980
rect 9600 6970 9640 6980
rect 1920 6960 1960 6970
rect 3160 6960 3280 6970
rect 3680 6960 3760 6970
rect 3800 6960 3840 6970
rect 3920 6960 4000 6970
rect 9600 6960 9640 6970
rect 1920 6950 1960 6960
rect 3160 6950 3280 6960
rect 3680 6950 3760 6960
rect 3800 6950 3840 6960
rect 3920 6950 4000 6960
rect 9600 6950 9640 6960
rect 1920 6940 1960 6950
rect 3160 6940 3280 6950
rect 3680 6940 3760 6950
rect 3800 6940 3840 6950
rect 3920 6940 4000 6950
rect 9600 6940 9640 6950
rect 1880 6930 1920 6940
rect 2480 6930 2560 6940
rect 3200 6930 3440 6940
rect 3800 6930 4000 6940
rect 1880 6920 1920 6930
rect 2480 6920 2560 6930
rect 3200 6920 3440 6930
rect 3800 6920 4000 6930
rect 1880 6910 1920 6920
rect 2480 6910 2560 6920
rect 3200 6910 3440 6920
rect 3800 6910 4000 6920
rect 1880 6900 1920 6910
rect 2480 6900 2560 6910
rect 3200 6900 3440 6910
rect 3800 6900 4000 6910
rect 2520 6890 2640 6900
rect 2920 6890 2960 6900
rect 3080 6890 3120 6900
rect 3160 6890 3400 6900
rect 3480 6890 3520 6900
rect 3880 6890 4000 6900
rect 2520 6880 2640 6890
rect 2920 6880 2960 6890
rect 3080 6880 3120 6890
rect 3160 6880 3400 6890
rect 3480 6880 3520 6890
rect 3880 6880 4000 6890
rect 2520 6870 2640 6880
rect 2920 6870 2960 6880
rect 3080 6870 3120 6880
rect 3160 6870 3400 6880
rect 3480 6870 3520 6880
rect 3880 6870 4000 6880
rect 2520 6860 2640 6870
rect 2920 6860 2960 6870
rect 3080 6860 3120 6870
rect 3160 6860 3400 6870
rect 3480 6860 3520 6870
rect 3880 6860 4000 6870
rect 2560 6850 2800 6860
rect 3040 6850 3440 6860
rect 3560 6850 3600 6860
rect 3880 6850 3960 6860
rect 2560 6840 2800 6850
rect 3040 6840 3440 6850
rect 3560 6840 3600 6850
rect 3880 6840 3960 6850
rect 2560 6830 2800 6840
rect 3040 6830 3440 6840
rect 3560 6830 3600 6840
rect 3880 6830 3960 6840
rect 2560 6820 2800 6830
rect 3040 6820 3440 6830
rect 3560 6820 3600 6830
rect 3880 6820 3960 6830
rect 1840 6810 1880 6820
rect 2760 6810 3280 6820
rect 3880 6810 3960 6820
rect 1840 6800 1880 6810
rect 2760 6800 3280 6810
rect 3880 6800 3960 6810
rect 1840 6790 1880 6800
rect 2760 6790 3280 6800
rect 3880 6790 3960 6800
rect 1840 6780 1880 6790
rect 2760 6780 3280 6790
rect 3880 6780 3960 6790
rect 1840 6770 1880 6780
rect 3040 6770 3400 6780
rect 3680 6770 3720 6780
rect 3920 6770 3960 6780
rect 9560 6770 9600 6780
rect 1840 6760 1880 6770
rect 3040 6760 3400 6770
rect 3680 6760 3720 6770
rect 3920 6760 3960 6770
rect 9560 6760 9600 6770
rect 1840 6750 1880 6760
rect 3040 6750 3400 6760
rect 3680 6750 3720 6760
rect 3920 6750 3960 6760
rect 9560 6750 9600 6760
rect 1840 6740 1880 6750
rect 3040 6740 3400 6750
rect 3680 6740 3720 6750
rect 3920 6740 3960 6750
rect 9560 6740 9600 6750
rect 1840 6730 1880 6740
rect 2280 6730 2480 6740
rect 3280 6730 3400 6740
rect 3920 6730 3960 6740
rect 9520 6730 9600 6740
rect 1840 6720 1880 6730
rect 2280 6720 2480 6730
rect 3280 6720 3400 6730
rect 3920 6720 3960 6730
rect 9520 6720 9600 6730
rect 1840 6710 1880 6720
rect 2280 6710 2480 6720
rect 3280 6710 3400 6720
rect 3920 6710 3960 6720
rect 9520 6710 9600 6720
rect 1840 6700 1880 6710
rect 2280 6700 2480 6710
rect 3280 6700 3400 6710
rect 3920 6700 3960 6710
rect 9520 6700 9600 6710
rect 1800 6690 1880 6700
rect 2240 6690 2280 6700
rect 2480 6690 2520 6700
rect 3440 6690 3520 6700
rect 9560 6690 9600 6700
rect 9960 6690 9990 6700
rect 1800 6680 1880 6690
rect 2240 6680 2280 6690
rect 2480 6680 2520 6690
rect 3440 6680 3520 6690
rect 9560 6680 9600 6690
rect 9960 6680 9990 6690
rect 1800 6670 1880 6680
rect 2240 6670 2280 6680
rect 2480 6670 2520 6680
rect 3440 6670 3520 6680
rect 9560 6670 9600 6680
rect 9960 6670 9990 6680
rect 1800 6660 1880 6670
rect 2240 6660 2280 6670
rect 2480 6660 2520 6670
rect 3440 6660 3520 6670
rect 9560 6660 9600 6670
rect 9960 6660 9990 6670
rect 1760 6650 1840 6660
rect 2520 6650 2560 6660
rect 3560 6650 3640 6660
rect 3840 6650 3880 6660
rect 3960 6650 4000 6660
rect 9480 6650 9560 6660
rect 9800 6650 9880 6660
rect 1760 6640 1840 6650
rect 2520 6640 2560 6650
rect 3560 6640 3640 6650
rect 3840 6640 3880 6650
rect 3960 6640 4000 6650
rect 9480 6640 9560 6650
rect 9800 6640 9880 6650
rect 1760 6630 1840 6640
rect 2520 6630 2560 6640
rect 3560 6630 3640 6640
rect 3840 6630 3880 6640
rect 3960 6630 4000 6640
rect 9480 6630 9560 6640
rect 9800 6630 9880 6640
rect 1760 6620 1840 6630
rect 2520 6620 2560 6630
rect 3560 6620 3640 6630
rect 3840 6620 3880 6630
rect 3960 6620 4000 6630
rect 9480 6620 9560 6630
rect 9800 6620 9880 6630
rect 1560 6610 1600 6620
rect 1640 6610 1680 6620
rect 2200 6610 2240 6620
rect 2560 6610 2600 6620
rect 3680 6610 3720 6620
rect 3880 6610 3920 6620
rect 3960 6610 4000 6620
rect 9520 6610 9640 6620
rect 9680 6610 9760 6620
rect 1560 6600 1600 6610
rect 1640 6600 1680 6610
rect 2200 6600 2240 6610
rect 2560 6600 2600 6610
rect 3680 6600 3720 6610
rect 3880 6600 3920 6610
rect 3960 6600 4000 6610
rect 9520 6600 9640 6610
rect 9680 6600 9760 6610
rect 1560 6590 1600 6600
rect 1640 6590 1680 6600
rect 2200 6590 2240 6600
rect 2560 6590 2600 6600
rect 3680 6590 3720 6600
rect 3880 6590 3920 6600
rect 3960 6590 4000 6600
rect 9520 6590 9640 6600
rect 9680 6590 9760 6600
rect 1560 6580 1600 6590
rect 1640 6580 1680 6590
rect 2200 6580 2240 6590
rect 2560 6580 2600 6590
rect 3680 6580 3720 6590
rect 3880 6580 3920 6590
rect 3960 6580 4000 6590
rect 9520 6580 9640 6590
rect 9680 6580 9760 6590
rect 1360 6570 1400 6580
rect 1480 6570 1520 6580
rect 1640 6570 1800 6580
rect 2560 6570 2600 6580
rect 3760 6570 3800 6580
rect 6000 6570 6480 6580
rect 6560 6570 6600 6580
rect 9480 6570 9520 6580
rect 1360 6560 1400 6570
rect 1480 6560 1520 6570
rect 1640 6560 1800 6570
rect 2560 6560 2600 6570
rect 3760 6560 3800 6570
rect 6000 6560 6480 6570
rect 6560 6560 6600 6570
rect 9480 6560 9520 6570
rect 1360 6550 1400 6560
rect 1480 6550 1520 6560
rect 1640 6550 1800 6560
rect 2560 6550 2600 6560
rect 3760 6550 3800 6560
rect 6000 6550 6480 6560
rect 6560 6550 6600 6560
rect 9480 6550 9520 6560
rect 1360 6540 1400 6550
rect 1480 6540 1520 6550
rect 1640 6540 1800 6550
rect 2560 6540 2600 6550
rect 3760 6540 3800 6550
rect 6000 6540 6480 6550
rect 6560 6540 6600 6550
rect 9480 6540 9520 6550
rect 1320 6530 1360 6540
rect 2240 6530 2280 6540
rect 2520 6530 2560 6540
rect 3840 6530 3880 6540
rect 4000 6530 4040 6540
rect 5840 6530 5880 6540
rect 5960 6530 6320 6540
rect 6560 6530 6680 6540
rect 9920 6530 9990 6540
rect 1320 6520 1360 6530
rect 2240 6520 2280 6530
rect 2520 6520 2560 6530
rect 3840 6520 3880 6530
rect 4000 6520 4040 6530
rect 5840 6520 5880 6530
rect 5960 6520 6320 6530
rect 6560 6520 6680 6530
rect 9920 6520 9990 6530
rect 1320 6510 1360 6520
rect 2240 6510 2280 6520
rect 2520 6510 2560 6520
rect 3840 6510 3880 6520
rect 4000 6510 4040 6520
rect 5840 6510 5880 6520
rect 5960 6510 6320 6520
rect 6560 6510 6680 6520
rect 9920 6510 9990 6520
rect 1320 6500 1360 6510
rect 2240 6500 2280 6510
rect 2520 6500 2560 6510
rect 3840 6500 3880 6510
rect 4000 6500 4040 6510
rect 5840 6500 5880 6510
rect 5960 6500 6320 6510
rect 6560 6500 6680 6510
rect 9920 6500 9990 6510
rect 1240 6490 1280 6500
rect 2120 6490 2160 6500
rect 2240 6490 2280 6500
rect 3960 6490 4040 6500
rect 5800 6490 5880 6500
rect 5960 6490 6080 6500
rect 6600 6490 6720 6500
rect 9800 6490 9880 6500
rect 1240 6480 1280 6490
rect 2120 6480 2160 6490
rect 2240 6480 2280 6490
rect 3960 6480 4040 6490
rect 5800 6480 5880 6490
rect 5960 6480 6080 6490
rect 6600 6480 6720 6490
rect 9800 6480 9880 6490
rect 1240 6470 1280 6480
rect 2120 6470 2160 6480
rect 2240 6470 2280 6480
rect 3960 6470 4040 6480
rect 5800 6470 5880 6480
rect 5960 6470 6080 6480
rect 6600 6470 6720 6480
rect 9800 6470 9880 6480
rect 1240 6460 1280 6470
rect 2120 6460 2160 6470
rect 2240 6460 2280 6470
rect 3960 6460 4040 6470
rect 5800 6460 5880 6470
rect 5960 6460 6080 6470
rect 6600 6460 6720 6470
rect 9800 6460 9880 6470
rect 1320 6450 1360 6460
rect 1680 6450 1760 6460
rect 2120 6450 2160 6460
rect 2280 6450 2320 6460
rect 2360 6450 2400 6460
rect 2520 6450 2560 6460
rect 3960 6450 4000 6460
rect 5720 6450 6080 6460
rect 6600 6450 6800 6460
rect 1320 6440 1360 6450
rect 1680 6440 1760 6450
rect 2120 6440 2160 6450
rect 2280 6440 2320 6450
rect 2360 6440 2400 6450
rect 2520 6440 2560 6450
rect 3960 6440 4000 6450
rect 5720 6440 6080 6450
rect 6600 6440 6800 6450
rect 1320 6430 1360 6440
rect 1680 6430 1760 6440
rect 2120 6430 2160 6440
rect 2280 6430 2320 6440
rect 2360 6430 2400 6440
rect 2520 6430 2560 6440
rect 3960 6430 4000 6440
rect 5720 6430 6080 6440
rect 6600 6430 6800 6440
rect 1320 6420 1360 6430
rect 1680 6420 1760 6430
rect 2120 6420 2160 6430
rect 2280 6420 2320 6430
rect 2360 6420 2400 6430
rect 2520 6420 2560 6430
rect 3960 6420 4000 6430
rect 5720 6420 6080 6430
rect 6600 6420 6800 6430
rect 1200 6410 1360 6420
rect 1720 6410 1960 6420
rect 2040 6410 2120 6420
rect 2360 6410 2400 6420
rect 5680 6410 6120 6420
rect 6720 6410 6840 6420
rect 1200 6400 1360 6410
rect 1720 6400 1960 6410
rect 2040 6400 2120 6410
rect 2360 6400 2400 6410
rect 5680 6400 6120 6410
rect 6720 6400 6840 6410
rect 1200 6390 1360 6400
rect 1720 6390 1960 6400
rect 2040 6390 2120 6400
rect 2360 6390 2400 6400
rect 5680 6390 6120 6400
rect 6720 6390 6840 6400
rect 1200 6380 1360 6390
rect 1720 6380 1960 6390
rect 2040 6380 2120 6390
rect 2360 6380 2400 6390
rect 5680 6380 6120 6390
rect 6720 6380 6840 6390
rect 1240 6370 1280 6380
rect 1600 6370 1720 6380
rect 1840 6370 1880 6380
rect 1960 6370 2040 6380
rect 4080 6370 4120 6380
rect 5640 6370 5800 6380
rect 5840 6370 6280 6380
rect 6320 6370 6360 6380
rect 6800 6370 6840 6380
rect 9600 6370 9640 6380
rect 1240 6360 1280 6370
rect 1600 6360 1720 6370
rect 1840 6360 1880 6370
rect 1960 6360 2040 6370
rect 4080 6360 4120 6370
rect 5640 6360 5800 6370
rect 5840 6360 6280 6370
rect 6320 6360 6360 6370
rect 6800 6360 6840 6370
rect 9600 6360 9640 6370
rect 1240 6350 1280 6360
rect 1600 6350 1720 6360
rect 1840 6350 1880 6360
rect 1960 6350 2040 6360
rect 4080 6350 4120 6360
rect 5640 6350 5800 6360
rect 5840 6350 6280 6360
rect 6320 6350 6360 6360
rect 6800 6350 6840 6360
rect 9600 6350 9640 6360
rect 1240 6340 1280 6350
rect 1600 6340 1720 6350
rect 1840 6340 1880 6350
rect 1960 6340 2040 6350
rect 4080 6340 4120 6350
rect 5640 6340 5800 6350
rect 5840 6340 6280 6350
rect 6320 6340 6360 6350
rect 6800 6340 6840 6350
rect 9600 6340 9640 6350
rect 1200 6330 1320 6340
rect 1600 6330 1640 6340
rect 1840 6330 1880 6340
rect 4120 6330 4160 6340
rect 5400 6330 5480 6340
rect 5640 6330 5680 6340
rect 5800 6330 5840 6340
rect 6400 6330 6440 6340
rect 6800 6330 6840 6340
rect 9320 6330 9520 6340
rect 1200 6320 1320 6330
rect 1600 6320 1640 6330
rect 1840 6320 1880 6330
rect 4120 6320 4160 6330
rect 5400 6320 5480 6330
rect 5640 6320 5680 6330
rect 5800 6320 5840 6330
rect 6400 6320 6440 6330
rect 6800 6320 6840 6330
rect 9320 6320 9520 6330
rect 1200 6310 1320 6320
rect 1600 6310 1640 6320
rect 1840 6310 1880 6320
rect 4120 6310 4160 6320
rect 5400 6310 5480 6320
rect 5640 6310 5680 6320
rect 5800 6310 5840 6320
rect 6400 6310 6440 6320
rect 6800 6310 6840 6320
rect 9320 6310 9520 6320
rect 1200 6300 1320 6310
rect 1600 6300 1640 6310
rect 1840 6300 1880 6310
rect 4120 6300 4160 6310
rect 5400 6300 5480 6310
rect 5640 6300 5680 6310
rect 5800 6300 5840 6310
rect 6400 6300 6440 6310
rect 6800 6300 6840 6310
rect 9320 6300 9520 6310
rect 1200 6290 1240 6300
rect 1280 6290 1320 6300
rect 4160 6290 4200 6300
rect 5640 6290 5720 6300
rect 6440 6290 6520 6300
rect 6800 6290 6840 6300
rect 9280 6290 9320 6300
rect 9400 6290 9440 6300
rect 9480 6290 9520 6300
rect 9960 6290 9990 6300
rect 1200 6280 1240 6290
rect 1280 6280 1320 6290
rect 4160 6280 4200 6290
rect 5640 6280 5720 6290
rect 6440 6280 6520 6290
rect 6800 6280 6840 6290
rect 9280 6280 9320 6290
rect 9400 6280 9440 6290
rect 9480 6280 9520 6290
rect 9960 6280 9990 6290
rect 1200 6270 1240 6280
rect 1280 6270 1320 6280
rect 4160 6270 4200 6280
rect 5640 6270 5720 6280
rect 6440 6270 6520 6280
rect 6800 6270 6840 6280
rect 9280 6270 9320 6280
rect 9400 6270 9440 6280
rect 9480 6270 9520 6280
rect 9960 6270 9990 6280
rect 1200 6260 1240 6270
rect 1280 6260 1320 6270
rect 4160 6260 4200 6270
rect 5640 6260 5720 6270
rect 6440 6260 6520 6270
rect 6800 6260 6840 6270
rect 9280 6260 9320 6270
rect 9400 6260 9440 6270
rect 9480 6260 9520 6270
rect 9960 6260 9990 6270
rect 1200 6250 1400 6260
rect 4200 6250 4240 6260
rect 5560 6250 5640 6260
rect 6520 6250 6560 6260
rect 6840 6250 6880 6260
rect 9240 6250 9320 6260
rect 9440 6250 9480 6260
rect 9600 6250 9640 6260
rect 9800 6250 9840 6260
rect 9920 6250 9960 6260
rect 1200 6240 1400 6250
rect 4200 6240 4240 6250
rect 5560 6240 5640 6250
rect 6520 6240 6560 6250
rect 6840 6240 6880 6250
rect 9240 6240 9320 6250
rect 9440 6240 9480 6250
rect 9600 6240 9640 6250
rect 9800 6240 9840 6250
rect 9920 6240 9960 6250
rect 1200 6230 1400 6240
rect 4200 6230 4240 6240
rect 5560 6230 5640 6240
rect 6520 6230 6560 6240
rect 6840 6230 6880 6240
rect 9240 6230 9320 6240
rect 9440 6230 9480 6240
rect 9600 6230 9640 6240
rect 9800 6230 9840 6240
rect 9920 6230 9960 6240
rect 1200 6220 1400 6230
rect 4200 6220 4240 6230
rect 5560 6220 5640 6230
rect 6520 6220 6560 6230
rect 6840 6220 6880 6230
rect 9240 6220 9320 6230
rect 9440 6220 9480 6230
rect 9600 6220 9640 6230
rect 9800 6220 9840 6230
rect 9920 6220 9960 6230
rect 1160 6210 1320 6220
rect 1760 6210 1800 6220
rect 5280 6210 5320 6220
rect 5520 6210 5560 6220
rect 6560 6210 6640 6220
rect 6800 6210 6840 6220
rect 6880 6210 6920 6220
rect 9240 6210 9320 6220
rect 9600 6210 9640 6220
rect 9800 6210 9840 6220
rect 1160 6200 1320 6210
rect 1760 6200 1800 6210
rect 5280 6200 5320 6210
rect 5520 6200 5560 6210
rect 6560 6200 6640 6210
rect 6800 6200 6840 6210
rect 6880 6200 6920 6210
rect 9240 6200 9320 6210
rect 9600 6200 9640 6210
rect 9800 6200 9840 6210
rect 1160 6190 1320 6200
rect 1760 6190 1800 6200
rect 5280 6190 5320 6200
rect 5520 6190 5560 6200
rect 6560 6190 6640 6200
rect 6800 6190 6840 6200
rect 6880 6190 6920 6200
rect 9240 6190 9320 6200
rect 9600 6190 9640 6200
rect 9800 6190 9840 6200
rect 1160 6180 1320 6190
rect 1760 6180 1800 6190
rect 5280 6180 5320 6190
rect 5520 6180 5560 6190
rect 6560 6180 6640 6190
rect 6800 6180 6840 6190
rect 6880 6180 6920 6190
rect 9240 6180 9320 6190
rect 9600 6180 9640 6190
rect 9800 6180 9840 6190
rect 1200 6170 1280 6180
rect 1760 6170 1800 6180
rect 5240 6170 5280 6180
rect 5440 6170 5480 6180
rect 6640 6170 6680 6180
rect 6880 6170 6960 6180
rect 9200 6170 9240 6180
rect 1200 6160 1280 6170
rect 1760 6160 1800 6170
rect 5240 6160 5280 6170
rect 5440 6160 5480 6170
rect 6640 6160 6680 6170
rect 6880 6160 6960 6170
rect 9200 6160 9240 6170
rect 1200 6150 1280 6160
rect 1760 6150 1800 6160
rect 5240 6150 5280 6160
rect 5440 6150 5480 6160
rect 6640 6150 6680 6160
rect 6880 6150 6960 6160
rect 9200 6150 9240 6160
rect 1200 6140 1280 6150
rect 1760 6140 1800 6150
rect 5240 6140 5280 6150
rect 5440 6140 5480 6150
rect 6640 6140 6680 6150
rect 6880 6140 6960 6150
rect 9200 6140 9240 6150
rect 1120 6130 1160 6140
rect 1200 6130 1280 6140
rect 1640 6130 1680 6140
rect 1720 6130 1800 6140
rect 4280 6130 4320 6140
rect 5240 6130 5280 6140
rect 5400 6130 5440 6140
rect 6640 6130 6680 6140
rect 6920 6130 7000 6140
rect 9120 6130 9160 6140
rect 9840 6130 9960 6140
rect 1120 6120 1160 6130
rect 1200 6120 1280 6130
rect 1640 6120 1680 6130
rect 1720 6120 1800 6130
rect 4280 6120 4320 6130
rect 5240 6120 5280 6130
rect 5400 6120 5440 6130
rect 6640 6120 6680 6130
rect 6920 6120 7000 6130
rect 9120 6120 9160 6130
rect 9840 6120 9960 6130
rect 1120 6110 1160 6120
rect 1200 6110 1280 6120
rect 1640 6110 1680 6120
rect 1720 6110 1800 6120
rect 4280 6110 4320 6120
rect 5240 6110 5280 6120
rect 5400 6110 5440 6120
rect 6640 6110 6680 6120
rect 6920 6110 7000 6120
rect 9120 6110 9160 6120
rect 9840 6110 9960 6120
rect 1120 6100 1160 6110
rect 1200 6100 1280 6110
rect 1640 6100 1680 6110
rect 1720 6100 1800 6110
rect 4280 6100 4320 6110
rect 5240 6100 5280 6110
rect 5400 6100 5440 6110
rect 6640 6100 6680 6110
rect 6920 6100 7000 6110
rect 9120 6100 9160 6110
rect 9840 6100 9960 6110
rect 1120 6090 1280 6100
rect 1680 6090 1760 6100
rect 5200 6090 5240 6100
rect 6680 6090 6720 6100
rect 6960 6090 7000 6100
rect 9000 6090 9080 6100
rect 9840 6090 9960 6100
rect 1120 6080 1280 6090
rect 1680 6080 1760 6090
rect 5200 6080 5240 6090
rect 6680 6080 6720 6090
rect 6960 6080 7000 6090
rect 9000 6080 9080 6090
rect 9840 6080 9960 6090
rect 1120 6070 1280 6080
rect 1680 6070 1760 6080
rect 5200 6070 5240 6080
rect 6680 6070 6720 6080
rect 6960 6070 7000 6080
rect 9000 6070 9080 6080
rect 9840 6070 9960 6080
rect 1120 6060 1280 6070
rect 1680 6060 1760 6070
rect 5200 6060 5240 6070
rect 6680 6060 6720 6070
rect 6960 6060 7000 6070
rect 9000 6060 9080 6070
rect 9840 6060 9960 6070
rect 800 6050 960 6060
rect 1040 6050 1200 6060
rect 1240 6050 1280 6060
rect 1720 6050 1760 6060
rect 2440 6050 2480 6060
rect 4320 6050 4360 6060
rect 5200 6050 5240 6060
rect 5360 6050 5400 6060
rect 6960 6050 7000 6060
rect 8840 6050 8920 6060
rect 9200 6050 9240 6060
rect 9280 6050 9320 6060
rect 800 6040 960 6050
rect 1040 6040 1200 6050
rect 1240 6040 1280 6050
rect 1720 6040 1760 6050
rect 2440 6040 2480 6050
rect 4320 6040 4360 6050
rect 5200 6040 5240 6050
rect 5360 6040 5400 6050
rect 6960 6040 7000 6050
rect 8840 6040 8920 6050
rect 9200 6040 9240 6050
rect 9280 6040 9320 6050
rect 800 6030 960 6040
rect 1040 6030 1200 6040
rect 1240 6030 1280 6040
rect 1720 6030 1760 6040
rect 2440 6030 2480 6040
rect 4320 6030 4360 6040
rect 5200 6030 5240 6040
rect 5360 6030 5400 6040
rect 6960 6030 7000 6040
rect 8840 6030 8920 6040
rect 9200 6030 9240 6040
rect 9280 6030 9320 6040
rect 800 6020 960 6030
rect 1040 6020 1200 6030
rect 1240 6020 1280 6030
rect 1720 6020 1760 6030
rect 2440 6020 2480 6030
rect 4320 6020 4360 6030
rect 5200 6020 5240 6030
rect 5360 6020 5400 6030
rect 6960 6020 7000 6030
rect 8840 6020 8920 6030
rect 9200 6020 9240 6030
rect 9280 6020 9320 6030
rect 760 6010 840 6020
rect 960 6010 1040 6020
rect 1080 6010 1120 6020
rect 1720 6010 1800 6020
rect 2480 6010 2520 6020
rect 5160 6010 5200 6020
rect 5360 6010 5400 6020
rect 6720 6010 6760 6020
rect 6960 6010 7000 6020
rect 8720 6010 8760 6020
rect 9080 6010 9200 6020
rect 9440 6010 9480 6020
rect 9880 6010 9960 6020
rect 760 6000 840 6010
rect 960 6000 1040 6010
rect 1080 6000 1120 6010
rect 1720 6000 1800 6010
rect 2480 6000 2520 6010
rect 5160 6000 5200 6010
rect 5360 6000 5400 6010
rect 6720 6000 6760 6010
rect 6960 6000 7000 6010
rect 8720 6000 8760 6010
rect 9080 6000 9200 6010
rect 9440 6000 9480 6010
rect 9880 6000 9960 6010
rect 760 5990 840 6000
rect 960 5990 1040 6000
rect 1080 5990 1120 6000
rect 1720 5990 1800 6000
rect 2480 5990 2520 6000
rect 5160 5990 5200 6000
rect 5360 5990 5400 6000
rect 6720 5990 6760 6000
rect 6960 5990 7000 6000
rect 8720 5990 8760 6000
rect 9080 5990 9200 6000
rect 9440 5990 9480 6000
rect 9880 5990 9960 6000
rect 760 5980 840 5990
rect 960 5980 1040 5990
rect 1080 5980 1120 5990
rect 1720 5980 1800 5990
rect 2480 5980 2520 5990
rect 5160 5980 5200 5990
rect 5360 5980 5400 5990
rect 6720 5980 6760 5990
rect 6960 5980 7000 5990
rect 8720 5980 8760 5990
rect 9080 5980 9200 5990
rect 9440 5980 9480 5990
rect 9880 5980 9960 5990
rect 720 5970 920 5980
rect 1720 5970 1800 5980
rect 2480 5970 2520 5980
rect 3760 5970 3800 5980
rect 4080 5970 4120 5980
rect 6720 5970 6760 5980
rect 8600 5970 8640 5980
rect 8960 5970 9040 5980
rect 9120 5970 9160 5980
rect 9280 5970 9320 5980
rect 9400 5970 9440 5980
rect 9480 5970 9520 5980
rect 9920 5970 9960 5980
rect 720 5960 920 5970
rect 1720 5960 1800 5970
rect 2480 5960 2520 5970
rect 3760 5960 3800 5970
rect 4080 5960 4120 5970
rect 6720 5960 6760 5970
rect 8600 5960 8640 5970
rect 8960 5960 9040 5970
rect 9120 5960 9160 5970
rect 9280 5960 9320 5970
rect 9400 5960 9440 5970
rect 9480 5960 9520 5970
rect 9920 5960 9960 5970
rect 720 5950 920 5960
rect 1720 5950 1800 5960
rect 2480 5950 2520 5960
rect 3760 5950 3800 5960
rect 4080 5950 4120 5960
rect 6720 5950 6760 5960
rect 8600 5950 8640 5960
rect 8960 5950 9040 5960
rect 9120 5950 9160 5960
rect 9280 5950 9320 5960
rect 9400 5950 9440 5960
rect 9480 5950 9520 5960
rect 9920 5950 9960 5960
rect 720 5940 920 5950
rect 1720 5940 1800 5950
rect 2480 5940 2520 5950
rect 3760 5940 3800 5950
rect 4080 5940 4120 5950
rect 6720 5940 6760 5950
rect 8600 5940 8640 5950
rect 8960 5940 9040 5950
rect 9120 5940 9160 5950
rect 9280 5940 9320 5950
rect 9400 5940 9440 5950
rect 9480 5940 9520 5950
rect 9920 5940 9960 5950
rect 680 5930 720 5940
rect 760 5930 840 5940
rect 920 5930 960 5940
rect 1720 5930 1760 5940
rect 2440 5930 2560 5940
rect 3160 5930 3200 5940
rect 3880 5930 3920 5940
rect 4160 5930 4200 5940
rect 4320 5930 4360 5940
rect 5120 5930 5160 5940
rect 6760 5930 6800 5940
rect 8480 5930 8520 5940
rect 8800 5930 8840 5940
rect 8920 5930 9000 5940
rect 9240 5930 9280 5940
rect 9360 5930 9440 5940
rect 9880 5930 9920 5940
rect 680 5920 720 5930
rect 760 5920 840 5930
rect 920 5920 960 5930
rect 1720 5920 1760 5930
rect 2440 5920 2560 5930
rect 3160 5920 3200 5930
rect 3880 5920 3920 5930
rect 4160 5920 4200 5930
rect 4320 5920 4360 5930
rect 5120 5920 5160 5930
rect 6760 5920 6800 5930
rect 8480 5920 8520 5930
rect 8800 5920 8840 5930
rect 8920 5920 9000 5930
rect 9240 5920 9280 5930
rect 9360 5920 9440 5930
rect 9880 5920 9920 5930
rect 680 5910 720 5920
rect 760 5910 840 5920
rect 920 5910 960 5920
rect 1720 5910 1760 5920
rect 2440 5910 2560 5920
rect 3160 5910 3200 5920
rect 3880 5910 3920 5920
rect 4160 5910 4200 5920
rect 4320 5910 4360 5920
rect 5120 5910 5160 5920
rect 6760 5910 6800 5920
rect 8480 5910 8520 5920
rect 8800 5910 8840 5920
rect 8920 5910 9000 5920
rect 9240 5910 9280 5920
rect 9360 5910 9440 5920
rect 9880 5910 9920 5920
rect 680 5900 720 5910
rect 760 5900 840 5910
rect 920 5900 960 5910
rect 1720 5900 1760 5910
rect 2440 5900 2560 5910
rect 3160 5900 3200 5910
rect 3880 5900 3920 5910
rect 4160 5900 4200 5910
rect 4320 5900 4360 5910
rect 5120 5900 5160 5910
rect 6760 5900 6800 5910
rect 8480 5900 8520 5910
rect 8800 5900 8840 5910
rect 8920 5900 9000 5910
rect 9240 5900 9280 5910
rect 9360 5900 9440 5910
rect 9880 5900 9920 5910
rect 640 5890 680 5900
rect 800 5890 840 5900
rect 920 5890 960 5900
rect 1840 5890 1880 5900
rect 2320 5890 2600 5900
rect 3120 5890 3240 5900
rect 5320 5890 5360 5900
rect 6760 5890 6800 5900
rect 8320 5890 8400 5900
rect 8640 5890 8760 5900
rect 8880 5890 8920 5900
rect 8960 5890 9000 5900
rect 9200 5890 9240 5900
rect 9320 5890 9360 5900
rect 640 5880 680 5890
rect 800 5880 840 5890
rect 920 5880 960 5890
rect 1840 5880 1880 5890
rect 2320 5880 2600 5890
rect 3120 5880 3240 5890
rect 5320 5880 5360 5890
rect 6760 5880 6800 5890
rect 8320 5880 8400 5890
rect 8640 5880 8760 5890
rect 8880 5880 8920 5890
rect 8960 5880 9000 5890
rect 9200 5880 9240 5890
rect 9320 5880 9360 5890
rect 640 5870 680 5880
rect 800 5870 840 5880
rect 920 5870 960 5880
rect 1840 5870 1880 5880
rect 2320 5870 2600 5880
rect 3120 5870 3240 5880
rect 5320 5870 5360 5880
rect 6760 5870 6800 5880
rect 8320 5870 8400 5880
rect 8640 5870 8760 5880
rect 8880 5870 8920 5880
rect 8960 5870 9000 5880
rect 9200 5870 9240 5880
rect 9320 5870 9360 5880
rect 640 5860 680 5870
rect 800 5860 840 5870
rect 920 5860 960 5870
rect 1840 5860 1880 5870
rect 2320 5860 2600 5870
rect 3120 5860 3240 5870
rect 5320 5860 5360 5870
rect 6760 5860 6800 5870
rect 8320 5860 8400 5870
rect 8640 5860 8760 5870
rect 8880 5860 8920 5870
rect 8960 5860 9000 5870
rect 9200 5860 9240 5870
rect 9320 5860 9360 5870
rect 560 5850 640 5860
rect 920 5850 960 5860
rect 1840 5850 1880 5860
rect 2280 5850 2320 5860
rect 2360 5850 2600 5860
rect 3040 5850 3240 5860
rect 3760 5850 3880 5860
rect 3920 5850 3960 5860
rect 5080 5850 5120 5860
rect 5320 5850 5360 5860
rect 6760 5850 6800 5860
rect 8200 5850 8240 5860
rect 8640 5850 8680 5860
rect 560 5840 640 5850
rect 920 5840 960 5850
rect 1840 5840 1880 5850
rect 2280 5840 2320 5850
rect 2360 5840 2600 5850
rect 3040 5840 3240 5850
rect 3760 5840 3880 5850
rect 3920 5840 3960 5850
rect 5080 5840 5120 5850
rect 5320 5840 5360 5850
rect 6760 5840 6800 5850
rect 8200 5840 8240 5850
rect 8640 5840 8680 5850
rect 560 5830 640 5840
rect 920 5830 960 5840
rect 1840 5830 1880 5840
rect 2280 5830 2320 5840
rect 2360 5830 2600 5840
rect 3040 5830 3240 5840
rect 3760 5830 3880 5840
rect 3920 5830 3960 5840
rect 5080 5830 5120 5840
rect 5320 5830 5360 5840
rect 6760 5830 6800 5840
rect 8200 5830 8240 5840
rect 8640 5830 8680 5840
rect 560 5820 640 5830
rect 920 5820 960 5830
rect 1840 5820 1880 5830
rect 2280 5820 2320 5830
rect 2360 5820 2600 5830
rect 3040 5820 3240 5830
rect 3760 5820 3880 5830
rect 3920 5820 3960 5830
rect 5080 5820 5120 5830
rect 5320 5820 5360 5830
rect 6760 5820 6800 5830
rect 8200 5820 8240 5830
rect 8640 5820 8680 5830
rect 600 5810 640 5820
rect 720 5810 760 5820
rect 840 5810 880 5820
rect 1880 5810 1920 5820
rect 2240 5810 2280 5820
rect 2360 5810 2400 5820
rect 2480 5810 2600 5820
rect 2960 5810 3120 5820
rect 3160 5810 3240 5820
rect 3840 5810 3920 5820
rect 5080 5810 5120 5820
rect 5320 5810 5360 5820
rect 8080 5810 8160 5820
rect 8800 5810 8880 5820
rect 9000 5810 9080 5820
rect 9920 5810 9960 5820
rect 600 5800 640 5810
rect 720 5800 760 5810
rect 840 5800 880 5810
rect 1880 5800 1920 5810
rect 2240 5800 2280 5810
rect 2360 5800 2400 5810
rect 2480 5800 2600 5810
rect 2960 5800 3120 5810
rect 3160 5800 3240 5810
rect 3840 5800 3920 5810
rect 5080 5800 5120 5810
rect 5320 5800 5360 5810
rect 8080 5800 8160 5810
rect 8800 5800 8880 5810
rect 9000 5800 9080 5810
rect 9920 5800 9960 5810
rect 600 5790 640 5800
rect 720 5790 760 5800
rect 840 5790 880 5800
rect 1880 5790 1920 5800
rect 2240 5790 2280 5800
rect 2360 5790 2400 5800
rect 2480 5790 2600 5800
rect 2960 5790 3120 5800
rect 3160 5790 3240 5800
rect 3840 5790 3920 5800
rect 5080 5790 5120 5800
rect 5320 5790 5360 5800
rect 8080 5790 8160 5800
rect 8800 5790 8880 5800
rect 9000 5790 9080 5800
rect 9920 5790 9960 5800
rect 600 5780 640 5790
rect 720 5780 760 5790
rect 840 5780 880 5790
rect 1880 5780 1920 5790
rect 2240 5780 2280 5790
rect 2360 5780 2400 5790
rect 2480 5780 2600 5790
rect 2960 5780 3120 5790
rect 3160 5780 3240 5790
rect 3840 5780 3920 5790
rect 5080 5780 5120 5790
rect 5320 5780 5360 5790
rect 8080 5780 8160 5790
rect 8800 5780 8880 5790
rect 9000 5780 9080 5790
rect 9920 5780 9960 5790
rect 560 5770 720 5780
rect 760 5770 880 5780
rect 1880 5770 1960 5780
rect 2200 5770 2240 5780
rect 2320 5770 2600 5780
rect 2960 5770 3040 5780
rect 3200 5770 3240 5780
rect 3960 5770 4000 5780
rect 6800 5770 6840 5780
rect 7920 5770 8000 5780
rect 8400 5770 8440 5780
rect 8680 5770 8760 5780
rect 8920 5770 8960 5780
rect 560 5760 720 5770
rect 760 5760 880 5770
rect 1880 5760 1960 5770
rect 2200 5760 2240 5770
rect 2320 5760 2600 5770
rect 2960 5760 3040 5770
rect 3200 5760 3240 5770
rect 3960 5760 4000 5770
rect 6800 5760 6840 5770
rect 7920 5760 8000 5770
rect 8400 5760 8440 5770
rect 8680 5760 8760 5770
rect 8920 5760 8960 5770
rect 560 5750 720 5760
rect 760 5750 880 5760
rect 1880 5750 1960 5760
rect 2200 5750 2240 5760
rect 2320 5750 2600 5760
rect 2960 5750 3040 5760
rect 3200 5750 3240 5760
rect 3960 5750 4000 5760
rect 6800 5750 6840 5760
rect 7920 5750 8000 5760
rect 8400 5750 8440 5760
rect 8680 5750 8760 5760
rect 8920 5750 8960 5760
rect 560 5740 720 5750
rect 760 5740 880 5750
rect 1880 5740 1960 5750
rect 2200 5740 2240 5750
rect 2320 5740 2600 5750
rect 2960 5740 3040 5750
rect 3200 5740 3240 5750
rect 3960 5740 4000 5750
rect 6800 5740 6840 5750
rect 7920 5740 8000 5750
rect 8400 5740 8440 5750
rect 8680 5740 8760 5750
rect 8920 5740 8960 5750
rect 600 5730 680 5740
rect 720 5730 800 5740
rect 1920 5730 1960 5740
rect 2280 5730 2520 5740
rect 2840 5730 3040 5740
rect 3200 5730 3240 5740
rect 5280 5730 5320 5740
rect 6800 5730 6840 5740
rect 6960 5730 7000 5740
rect 7760 5730 7880 5740
rect 8200 5730 8240 5740
rect 8680 5730 8760 5740
rect 600 5720 680 5730
rect 720 5720 800 5730
rect 1920 5720 1960 5730
rect 2280 5720 2520 5730
rect 2840 5720 3040 5730
rect 3200 5720 3240 5730
rect 5280 5720 5320 5730
rect 6800 5720 6840 5730
rect 6960 5720 7000 5730
rect 7760 5720 7880 5730
rect 8200 5720 8240 5730
rect 8680 5720 8760 5730
rect 600 5710 680 5720
rect 720 5710 800 5720
rect 1920 5710 1960 5720
rect 2280 5710 2520 5720
rect 2840 5710 3040 5720
rect 3200 5710 3240 5720
rect 5280 5710 5320 5720
rect 6800 5710 6840 5720
rect 6960 5710 7000 5720
rect 7760 5710 7880 5720
rect 8200 5710 8240 5720
rect 8680 5710 8760 5720
rect 600 5700 680 5710
rect 720 5700 800 5710
rect 1920 5700 1960 5710
rect 2280 5700 2520 5710
rect 2840 5700 3040 5710
rect 3200 5700 3240 5710
rect 5280 5700 5320 5710
rect 6800 5700 6840 5710
rect 6960 5700 7000 5710
rect 7760 5700 7880 5710
rect 8200 5700 8240 5710
rect 8680 5700 8760 5710
rect 1920 5690 1960 5700
rect 2160 5690 2200 5700
rect 2280 5690 2480 5700
rect 2800 5690 2840 5700
rect 2920 5690 3000 5700
rect 3160 5690 3240 5700
rect 5280 5690 5320 5700
rect 6960 5690 7000 5700
rect 7680 5690 7720 5700
rect 8120 5690 8280 5700
rect 1920 5680 1960 5690
rect 2160 5680 2200 5690
rect 2280 5680 2480 5690
rect 2800 5680 2840 5690
rect 2920 5680 3000 5690
rect 3160 5680 3240 5690
rect 5280 5680 5320 5690
rect 6960 5680 7000 5690
rect 7680 5680 7720 5690
rect 8120 5680 8280 5690
rect 1920 5670 1960 5680
rect 2160 5670 2200 5680
rect 2280 5670 2480 5680
rect 2800 5670 2840 5680
rect 2920 5670 3000 5680
rect 3160 5670 3240 5680
rect 5280 5670 5320 5680
rect 6960 5670 7000 5680
rect 7680 5670 7720 5680
rect 8120 5670 8280 5680
rect 1920 5660 1960 5670
rect 2160 5660 2200 5670
rect 2280 5660 2480 5670
rect 2800 5660 2840 5670
rect 2920 5660 3000 5670
rect 3160 5660 3240 5670
rect 5280 5660 5320 5670
rect 6960 5660 7000 5670
rect 7680 5660 7720 5670
rect 8120 5660 8280 5670
rect 520 5650 640 5660
rect 1960 5650 2000 5660
rect 2160 5650 2200 5660
rect 2240 5650 2360 5660
rect 2400 5650 2480 5660
rect 2720 5650 2840 5660
rect 3160 5650 3240 5660
rect 3800 5650 3840 5660
rect 3920 5650 3960 5660
rect 5080 5650 5120 5660
rect 5600 5650 5800 5660
rect 6960 5650 7000 5660
rect 7520 5650 7640 5660
rect 8080 5650 8120 5660
rect 8160 5650 8320 5660
rect 8400 5650 8440 5660
rect 520 5640 640 5650
rect 1960 5640 2000 5650
rect 2160 5640 2200 5650
rect 2240 5640 2360 5650
rect 2400 5640 2480 5650
rect 2720 5640 2840 5650
rect 3160 5640 3240 5650
rect 3800 5640 3840 5650
rect 3920 5640 3960 5650
rect 5080 5640 5120 5650
rect 5600 5640 5800 5650
rect 6960 5640 7000 5650
rect 7520 5640 7640 5650
rect 8080 5640 8120 5650
rect 8160 5640 8320 5650
rect 8400 5640 8440 5650
rect 520 5630 640 5640
rect 1960 5630 2000 5640
rect 2160 5630 2200 5640
rect 2240 5630 2360 5640
rect 2400 5630 2480 5640
rect 2720 5630 2840 5640
rect 3160 5630 3240 5640
rect 3800 5630 3840 5640
rect 3920 5630 3960 5640
rect 5080 5630 5120 5640
rect 5600 5630 5800 5640
rect 6960 5630 7000 5640
rect 7520 5630 7640 5640
rect 8080 5630 8120 5640
rect 8160 5630 8320 5640
rect 8400 5630 8440 5640
rect 520 5620 640 5630
rect 1960 5620 2000 5630
rect 2160 5620 2200 5630
rect 2240 5620 2360 5630
rect 2400 5620 2480 5630
rect 2720 5620 2840 5630
rect 3160 5620 3240 5630
rect 3800 5620 3840 5630
rect 3920 5620 3960 5630
rect 5080 5620 5120 5630
rect 5600 5620 5800 5630
rect 6960 5620 7000 5630
rect 7520 5620 7640 5630
rect 8080 5620 8120 5630
rect 8160 5620 8320 5630
rect 8400 5620 8440 5630
rect 520 5610 720 5620
rect 1960 5610 2040 5620
rect 2080 5610 2160 5620
rect 2240 5610 2360 5620
rect 2400 5610 2440 5620
rect 2720 5610 2920 5620
rect 3160 5610 3240 5620
rect 5080 5610 5120 5620
rect 5480 5610 5560 5620
rect 5840 5610 6080 5620
rect 6160 5610 6560 5620
rect 6840 5610 6880 5620
rect 6960 5610 7000 5620
rect 7400 5610 7440 5620
rect 8160 5610 8280 5620
rect 8360 5610 8400 5620
rect 9000 5610 9080 5620
rect 520 5600 720 5610
rect 1960 5600 2040 5610
rect 2080 5600 2160 5610
rect 2240 5600 2360 5610
rect 2400 5600 2440 5610
rect 2720 5600 2920 5610
rect 3160 5600 3240 5610
rect 5080 5600 5120 5610
rect 5480 5600 5560 5610
rect 5840 5600 6080 5610
rect 6160 5600 6560 5610
rect 6840 5600 6880 5610
rect 6960 5600 7000 5610
rect 7400 5600 7440 5610
rect 8160 5600 8280 5610
rect 8360 5600 8400 5610
rect 9000 5600 9080 5610
rect 520 5590 720 5600
rect 1960 5590 2040 5600
rect 2080 5590 2160 5600
rect 2240 5590 2360 5600
rect 2400 5590 2440 5600
rect 2720 5590 2920 5600
rect 3160 5590 3240 5600
rect 5080 5590 5120 5600
rect 5480 5590 5560 5600
rect 5840 5590 6080 5600
rect 6160 5590 6560 5600
rect 6840 5590 6880 5600
rect 6960 5590 7000 5600
rect 7400 5590 7440 5600
rect 8160 5590 8280 5600
rect 8360 5590 8400 5600
rect 9000 5590 9080 5600
rect 520 5580 720 5590
rect 1960 5580 2040 5590
rect 2080 5580 2160 5590
rect 2240 5580 2360 5590
rect 2400 5580 2440 5590
rect 2720 5580 2920 5590
rect 3160 5580 3240 5590
rect 5080 5580 5120 5590
rect 5480 5580 5560 5590
rect 5840 5580 6080 5590
rect 6160 5580 6560 5590
rect 6840 5580 6880 5590
rect 6960 5580 7000 5590
rect 7400 5580 7440 5590
rect 8160 5580 8280 5590
rect 8360 5580 8400 5590
rect 9000 5580 9080 5590
rect 520 5570 640 5580
rect 1960 5570 2160 5580
rect 2240 5570 2400 5580
rect 2680 5570 2880 5580
rect 2920 5570 3000 5580
rect 3160 5570 3240 5580
rect 3760 5570 3800 5580
rect 5080 5570 5120 5580
rect 5440 5570 5520 5580
rect 5920 5570 6200 5580
rect 6560 5570 6640 5580
rect 7280 5570 7320 5580
rect 7640 5570 7680 5580
rect 7720 5570 7760 5580
rect 7840 5570 7880 5580
rect 8080 5570 8240 5580
rect 8880 5570 8920 5580
rect 9000 5570 9080 5580
rect 520 5560 640 5570
rect 1960 5560 2160 5570
rect 2240 5560 2400 5570
rect 2680 5560 2880 5570
rect 2920 5560 3000 5570
rect 3160 5560 3240 5570
rect 3760 5560 3800 5570
rect 5080 5560 5120 5570
rect 5440 5560 5520 5570
rect 5920 5560 6200 5570
rect 6560 5560 6640 5570
rect 7280 5560 7320 5570
rect 7640 5560 7680 5570
rect 7720 5560 7760 5570
rect 7840 5560 7880 5570
rect 8080 5560 8240 5570
rect 8880 5560 8920 5570
rect 9000 5560 9080 5570
rect 520 5550 640 5560
rect 1960 5550 2160 5560
rect 2240 5550 2400 5560
rect 2680 5550 2880 5560
rect 2920 5550 3000 5560
rect 3160 5550 3240 5560
rect 3760 5550 3800 5560
rect 5080 5550 5120 5560
rect 5440 5550 5520 5560
rect 5920 5550 6200 5560
rect 6560 5550 6640 5560
rect 7280 5550 7320 5560
rect 7640 5550 7680 5560
rect 7720 5550 7760 5560
rect 7840 5550 7880 5560
rect 8080 5550 8240 5560
rect 8880 5550 8920 5560
rect 9000 5550 9080 5560
rect 520 5540 640 5550
rect 1960 5540 2160 5550
rect 2240 5540 2400 5550
rect 2680 5540 2880 5550
rect 2920 5540 3000 5550
rect 3160 5540 3240 5550
rect 3760 5540 3800 5550
rect 5080 5540 5120 5550
rect 5440 5540 5520 5550
rect 5920 5540 6200 5550
rect 6560 5540 6640 5550
rect 7280 5540 7320 5550
rect 7640 5540 7680 5550
rect 7720 5540 7760 5550
rect 7840 5540 7880 5550
rect 8080 5540 8240 5550
rect 8880 5540 8920 5550
rect 9000 5540 9080 5550
rect 440 5530 520 5540
rect 1960 5530 2160 5540
rect 2240 5530 2400 5540
rect 2680 5530 2840 5540
rect 3000 5530 3040 5540
rect 3160 5530 3200 5540
rect 3640 5530 3760 5540
rect 5080 5530 5120 5540
rect 5240 5530 5280 5540
rect 5400 5530 5640 5540
rect 5960 5530 6040 5540
rect 6120 5530 6160 5540
rect 6600 5530 6720 5540
rect 7280 5530 7400 5540
rect 7600 5530 7720 5540
rect 7920 5530 7960 5540
rect 8040 5530 8120 5540
rect 8800 5530 8840 5540
rect 9080 5530 9120 5540
rect 440 5520 520 5530
rect 1960 5520 2160 5530
rect 2240 5520 2400 5530
rect 2680 5520 2840 5530
rect 3000 5520 3040 5530
rect 3160 5520 3200 5530
rect 3640 5520 3760 5530
rect 5080 5520 5120 5530
rect 5240 5520 5280 5530
rect 5400 5520 5640 5530
rect 5960 5520 6040 5530
rect 6120 5520 6160 5530
rect 6600 5520 6720 5530
rect 7280 5520 7400 5530
rect 7600 5520 7720 5530
rect 7920 5520 7960 5530
rect 8040 5520 8120 5530
rect 8800 5520 8840 5530
rect 9080 5520 9120 5530
rect 440 5510 520 5520
rect 1960 5510 2160 5520
rect 2240 5510 2400 5520
rect 2680 5510 2840 5520
rect 3000 5510 3040 5520
rect 3160 5510 3200 5520
rect 3640 5510 3760 5520
rect 5080 5510 5120 5520
rect 5240 5510 5280 5520
rect 5400 5510 5640 5520
rect 5960 5510 6040 5520
rect 6120 5510 6160 5520
rect 6600 5510 6720 5520
rect 7280 5510 7400 5520
rect 7600 5510 7720 5520
rect 7920 5510 7960 5520
rect 8040 5510 8120 5520
rect 8800 5510 8840 5520
rect 9080 5510 9120 5520
rect 440 5500 520 5510
rect 1960 5500 2160 5510
rect 2240 5500 2400 5510
rect 2680 5500 2840 5510
rect 3000 5500 3040 5510
rect 3160 5500 3200 5510
rect 3640 5500 3760 5510
rect 5080 5500 5120 5510
rect 5240 5500 5280 5510
rect 5400 5500 5640 5510
rect 5960 5500 6040 5510
rect 6120 5500 6160 5510
rect 6600 5500 6720 5510
rect 7280 5500 7400 5510
rect 7600 5500 7720 5510
rect 7920 5500 7960 5510
rect 8040 5500 8120 5510
rect 8800 5500 8840 5510
rect 9080 5500 9120 5510
rect 400 5490 440 5500
rect 2000 5490 2160 5500
rect 2240 5490 2360 5500
rect 2600 5490 2760 5500
rect 3000 5490 3080 5500
rect 3120 5490 3200 5500
rect 3600 5490 3680 5500
rect 5080 5490 5120 5500
rect 5240 5490 5280 5500
rect 5400 5490 5520 5500
rect 5960 5490 6000 5500
rect 6120 5490 6160 5500
rect 6520 5490 6720 5500
rect 6880 5490 6920 5500
rect 7240 5490 7400 5500
rect 7560 5490 7680 5500
rect 7720 5490 7760 5500
rect 7840 5490 7880 5500
rect 7920 5490 7960 5500
rect 8600 5490 8640 5500
rect 8680 5490 8760 5500
rect 8840 5490 8880 5500
rect 9040 5490 9080 5500
rect 400 5480 440 5490
rect 2000 5480 2160 5490
rect 2240 5480 2360 5490
rect 2600 5480 2760 5490
rect 3000 5480 3080 5490
rect 3120 5480 3200 5490
rect 3600 5480 3680 5490
rect 5080 5480 5120 5490
rect 5240 5480 5280 5490
rect 5400 5480 5520 5490
rect 5960 5480 6000 5490
rect 6120 5480 6160 5490
rect 6520 5480 6720 5490
rect 6880 5480 6920 5490
rect 7240 5480 7400 5490
rect 7560 5480 7680 5490
rect 7720 5480 7760 5490
rect 7840 5480 7880 5490
rect 7920 5480 7960 5490
rect 8600 5480 8640 5490
rect 8680 5480 8760 5490
rect 8840 5480 8880 5490
rect 9040 5480 9080 5490
rect 400 5470 440 5480
rect 2000 5470 2160 5480
rect 2240 5470 2360 5480
rect 2600 5470 2760 5480
rect 3000 5470 3080 5480
rect 3120 5470 3200 5480
rect 3600 5470 3680 5480
rect 5080 5470 5120 5480
rect 5240 5470 5280 5480
rect 5400 5470 5520 5480
rect 5960 5470 6000 5480
rect 6120 5470 6160 5480
rect 6520 5470 6720 5480
rect 6880 5470 6920 5480
rect 7240 5470 7400 5480
rect 7560 5470 7680 5480
rect 7720 5470 7760 5480
rect 7840 5470 7880 5480
rect 7920 5470 7960 5480
rect 8600 5470 8640 5480
rect 8680 5470 8760 5480
rect 8840 5470 8880 5480
rect 9040 5470 9080 5480
rect 400 5460 440 5470
rect 2000 5460 2160 5470
rect 2240 5460 2360 5470
rect 2600 5460 2760 5470
rect 3000 5460 3080 5470
rect 3120 5460 3200 5470
rect 3600 5460 3680 5470
rect 5080 5460 5120 5470
rect 5240 5460 5280 5470
rect 5400 5460 5520 5470
rect 5960 5460 6000 5470
rect 6120 5460 6160 5470
rect 6520 5460 6720 5470
rect 6880 5460 6920 5470
rect 7240 5460 7400 5470
rect 7560 5460 7680 5470
rect 7720 5460 7760 5470
rect 7840 5460 7880 5470
rect 7920 5460 7960 5470
rect 8600 5460 8640 5470
rect 8680 5460 8760 5470
rect 8840 5460 8880 5470
rect 9040 5460 9080 5470
rect 560 5450 600 5460
rect 2000 5450 2160 5460
rect 2240 5450 2360 5460
rect 2680 5450 2760 5460
rect 3040 5450 3160 5460
rect 5080 5450 5120 5460
rect 5400 5450 5440 5460
rect 5960 5450 6000 5460
rect 6120 5450 6160 5460
rect 6560 5450 6720 5460
rect 6880 5450 6920 5460
rect 7200 5450 7240 5460
rect 7600 5450 7640 5460
rect 7720 5450 7840 5460
rect 7880 5450 7920 5460
rect 8560 5450 8800 5460
rect 8920 5450 9080 5460
rect 560 5440 600 5450
rect 2000 5440 2160 5450
rect 2240 5440 2360 5450
rect 2680 5440 2760 5450
rect 3040 5440 3160 5450
rect 5080 5440 5120 5450
rect 5400 5440 5440 5450
rect 5960 5440 6000 5450
rect 6120 5440 6160 5450
rect 6560 5440 6720 5450
rect 6880 5440 6920 5450
rect 7200 5440 7240 5450
rect 7600 5440 7640 5450
rect 7720 5440 7840 5450
rect 7880 5440 7920 5450
rect 8560 5440 8800 5450
rect 8920 5440 9080 5450
rect 560 5430 600 5440
rect 2000 5430 2160 5440
rect 2240 5430 2360 5440
rect 2680 5430 2760 5440
rect 3040 5430 3160 5440
rect 5080 5430 5120 5440
rect 5400 5430 5440 5440
rect 5960 5430 6000 5440
rect 6120 5430 6160 5440
rect 6560 5430 6720 5440
rect 6880 5430 6920 5440
rect 7200 5430 7240 5440
rect 7600 5430 7640 5440
rect 7720 5430 7840 5440
rect 7880 5430 7920 5440
rect 8560 5430 8800 5440
rect 8920 5430 9080 5440
rect 560 5420 600 5430
rect 2000 5420 2160 5430
rect 2240 5420 2360 5430
rect 2680 5420 2760 5430
rect 3040 5420 3160 5430
rect 5080 5420 5120 5430
rect 5400 5420 5440 5430
rect 5960 5420 6000 5430
rect 6120 5420 6160 5430
rect 6560 5420 6720 5430
rect 6880 5420 6920 5430
rect 7200 5420 7240 5430
rect 7600 5420 7640 5430
rect 7720 5420 7840 5430
rect 7880 5420 7920 5430
rect 8560 5420 8800 5430
rect 8920 5420 9080 5430
rect 400 5410 440 5420
rect 480 5410 520 5420
rect 2040 5410 2160 5420
rect 2240 5410 2360 5420
rect 3560 5410 3600 5420
rect 5920 5410 5960 5420
rect 6120 5410 6160 5420
rect 6680 5410 6720 5420
rect 6880 5410 6960 5420
rect 7240 5410 7320 5420
rect 7560 5410 7600 5420
rect 7680 5410 7760 5420
rect 8400 5410 8440 5420
rect 8600 5410 8640 5420
rect 8680 5410 8720 5420
rect 8760 5410 8800 5420
rect 8920 5410 8960 5420
rect 9000 5410 9080 5420
rect 9480 5410 9600 5420
rect 400 5400 440 5410
rect 480 5400 520 5410
rect 2040 5400 2160 5410
rect 2240 5400 2360 5410
rect 3560 5400 3600 5410
rect 5920 5400 5960 5410
rect 6120 5400 6160 5410
rect 6680 5400 6720 5410
rect 6880 5400 6960 5410
rect 7240 5400 7320 5410
rect 7560 5400 7600 5410
rect 7680 5400 7760 5410
rect 8400 5400 8440 5410
rect 8600 5400 8640 5410
rect 8680 5400 8720 5410
rect 8760 5400 8800 5410
rect 8920 5400 8960 5410
rect 9000 5400 9080 5410
rect 9480 5400 9600 5410
rect 400 5390 440 5400
rect 480 5390 520 5400
rect 2040 5390 2160 5400
rect 2240 5390 2360 5400
rect 3560 5390 3600 5400
rect 5920 5390 5960 5400
rect 6120 5390 6160 5400
rect 6680 5390 6720 5400
rect 6880 5390 6960 5400
rect 7240 5390 7320 5400
rect 7560 5390 7600 5400
rect 7680 5390 7760 5400
rect 8400 5390 8440 5400
rect 8600 5390 8640 5400
rect 8680 5390 8720 5400
rect 8760 5390 8800 5400
rect 8920 5390 8960 5400
rect 9000 5390 9080 5400
rect 9480 5390 9600 5400
rect 400 5380 440 5390
rect 480 5380 520 5390
rect 2040 5380 2160 5390
rect 2240 5380 2360 5390
rect 3560 5380 3600 5390
rect 5920 5380 5960 5390
rect 6120 5380 6160 5390
rect 6680 5380 6720 5390
rect 6880 5380 6960 5390
rect 7240 5380 7320 5390
rect 7560 5380 7600 5390
rect 7680 5380 7760 5390
rect 8400 5380 8440 5390
rect 8600 5380 8640 5390
rect 8680 5380 8720 5390
rect 8760 5380 8800 5390
rect 8920 5380 8960 5390
rect 9000 5380 9080 5390
rect 9480 5380 9600 5390
rect 280 5370 360 5380
rect 440 5370 560 5380
rect 2040 5370 2160 5380
rect 2240 5370 2360 5380
rect 5360 5370 5400 5380
rect 5920 5370 5960 5380
rect 6720 5370 6760 5380
rect 6920 5370 6960 5380
rect 7240 5370 7320 5380
rect 7520 5370 7560 5380
rect 8520 5370 8600 5380
rect 8680 5370 8720 5380
rect 9280 5370 9360 5380
rect 9400 5370 9440 5380
rect 280 5360 360 5370
rect 440 5360 560 5370
rect 2040 5360 2160 5370
rect 2240 5360 2360 5370
rect 5360 5360 5400 5370
rect 5920 5360 5960 5370
rect 6720 5360 6760 5370
rect 6920 5360 6960 5370
rect 7240 5360 7320 5370
rect 7520 5360 7560 5370
rect 8520 5360 8600 5370
rect 8680 5360 8720 5370
rect 9280 5360 9360 5370
rect 9400 5360 9440 5370
rect 280 5350 360 5360
rect 440 5350 560 5360
rect 2040 5350 2160 5360
rect 2240 5350 2360 5360
rect 5360 5350 5400 5360
rect 5920 5350 5960 5360
rect 6720 5350 6760 5360
rect 6920 5350 6960 5360
rect 7240 5350 7320 5360
rect 7520 5350 7560 5360
rect 8520 5350 8600 5360
rect 8680 5350 8720 5360
rect 9280 5350 9360 5360
rect 9400 5350 9440 5360
rect 280 5340 360 5350
rect 440 5340 560 5350
rect 2040 5340 2160 5350
rect 2240 5340 2360 5350
rect 5360 5340 5400 5350
rect 5920 5340 5960 5350
rect 6720 5340 6760 5350
rect 6920 5340 6960 5350
rect 7240 5340 7320 5350
rect 7520 5340 7560 5350
rect 8520 5340 8600 5350
rect 8680 5340 8720 5350
rect 9280 5340 9360 5350
rect 9400 5340 9440 5350
rect 320 5330 560 5340
rect 2120 5330 2160 5340
rect 2240 5330 2360 5340
rect 5080 5330 5120 5340
rect 5200 5330 5240 5340
rect 5640 5330 5680 5340
rect 5880 5330 5920 5340
rect 6760 5330 6800 5340
rect 7240 5330 7280 5340
rect 8040 5330 8120 5340
rect 8280 5330 8320 5340
rect 8520 5330 8600 5340
rect 8680 5330 8760 5340
rect 9240 5330 9320 5340
rect 9400 5330 9480 5340
rect 320 5320 560 5330
rect 2120 5320 2160 5330
rect 2240 5320 2360 5330
rect 5080 5320 5120 5330
rect 5200 5320 5240 5330
rect 5640 5320 5680 5330
rect 5880 5320 5920 5330
rect 6760 5320 6800 5330
rect 7240 5320 7280 5330
rect 8040 5320 8120 5330
rect 8280 5320 8320 5330
rect 8520 5320 8600 5330
rect 8680 5320 8760 5330
rect 9240 5320 9320 5330
rect 9400 5320 9480 5330
rect 320 5310 560 5320
rect 2120 5310 2160 5320
rect 2240 5310 2360 5320
rect 5080 5310 5120 5320
rect 5200 5310 5240 5320
rect 5640 5310 5680 5320
rect 5880 5310 5920 5320
rect 6760 5310 6800 5320
rect 7240 5310 7280 5320
rect 8040 5310 8120 5320
rect 8280 5310 8320 5320
rect 8520 5310 8600 5320
rect 8680 5310 8760 5320
rect 9240 5310 9320 5320
rect 9400 5310 9480 5320
rect 320 5300 560 5310
rect 2120 5300 2160 5310
rect 2240 5300 2360 5310
rect 5080 5300 5120 5310
rect 5200 5300 5240 5310
rect 5640 5300 5680 5310
rect 5880 5300 5920 5310
rect 6760 5300 6800 5310
rect 7240 5300 7280 5310
rect 8040 5300 8120 5310
rect 8280 5300 8320 5310
rect 8520 5300 8600 5310
rect 8680 5300 8760 5310
rect 9240 5300 9320 5310
rect 9400 5300 9480 5310
rect 200 5290 600 5300
rect 2160 5290 2200 5300
rect 2240 5290 2360 5300
rect 2480 5290 2560 5300
rect 3520 5290 3560 5300
rect 5200 5290 5240 5300
rect 5560 5290 5680 5300
rect 5840 5290 5920 5300
rect 6160 5290 6200 5300
rect 6440 5290 6800 5300
rect 7240 5290 7280 5300
rect 8160 5290 8240 5300
rect 8360 5290 8520 5300
rect 8560 5290 8600 5300
rect 9040 5290 9080 5300
rect 9280 5290 9400 5300
rect 9440 5290 9480 5300
rect 9520 5290 9560 5300
rect 9960 5290 9990 5300
rect 200 5280 600 5290
rect 2160 5280 2200 5290
rect 2240 5280 2360 5290
rect 2480 5280 2560 5290
rect 3520 5280 3560 5290
rect 5200 5280 5240 5290
rect 5560 5280 5680 5290
rect 5840 5280 5920 5290
rect 6160 5280 6200 5290
rect 6440 5280 6800 5290
rect 7240 5280 7280 5290
rect 8160 5280 8240 5290
rect 8360 5280 8520 5290
rect 8560 5280 8600 5290
rect 9040 5280 9080 5290
rect 9280 5280 9400 5290
rect 9440 5280 9480 5290
rect 9520 5280 9560 5290
rect 9960 5280 9990 5290
rect 200 5270 600 5280
rect 2160 5270 2200 5280
rect 2240 5270 2360 5280
rect 2480 5270 2560 5280
rect 3520 5270 3560 5280
rect 5200 5270 5240 5280
rect 5560 5270 5680 5280
rect 5840 5270 5920 5280
rect 6160 5270 6200 5280
rect 6440 5270 6800 5280
rect 7240 5270 7280 5280
rect 8160 5270 8240 5280
rect 8360 5270 8520 5280
rect 8560 5270 8600 5280
rect 9040 5270 9080 5280
rect 9280 5270 9400 5280
rect 9440 5270 9480 5280
rect 9520 5270 9560 5280
rect 9960 5270 9990 5280
rect 200 5260 600 5270
rect 2160 5260 2200 5270
rect 2240 5260 2360 5270
rect 2480 5260 2560 5270
rect 3520 5260 3560 5270
rect 5200 5260 5240 5270
rect 5560 5260 5680 5270
rect 5840 5260 5920 5270
rect 6160 5260 6200 5270
rect 6440 5260 6800 5270
rect 7240 5260 7280 5270
rect 8160 5260 8240 5270
rect 8360 5260 8520 5270
rect 8560 5260 8600 5270
rect 9040 5260 9080 5270
rect 9280 5260 9400 5270
rect 9440 5260 9480 5270
rect 9520 5260 9560 5270
rect 9960 5260 9990 5270
rect 160 5250 600 5260
rect 2160 5250 2200 5260
rect 2240 5250 2400 5260
rect 2480 5250 2600 5260
rect 2640 5250 2680 5260
rect 2720 5250 2800 5260
rect 5040 5250 5080 5260
rect 5200 5250 5240 5260
rect 5560 5250 5680 5260
rect 5720 5250 5800 5260
rect 6200 5250 6320 5260
rect 6560 5250 6600 5260
rect 7240 5250 7280 5260
rect 8000 5250 8040 5260
rect 8160 5250 8240 5260
rect 8320 5250 8360 5260
rect 8400 5250 8440 5260
rect 8920 5250 9000 5260
rect 9120 5250 9200 5260
rect 9280 5250 9400 5260
rect 9720 5250 9760 5260
rect 9840 5250 9880 5260
rect 9960 5250 9990 5260
rect 160 5240 600 5250
rect 2160 5240 2200 5250
rect 2240 5240 2400 5250
rect 2480 5240 2600 5250
rect 2640 5240 2680 5250
rect 2720 5240 2800 5250
rect 5040 5240 5080 5250
rect 5200 5240 5240 5250
rect 5560 5240 5680 5250
rect 5720 5240 5800 5250
rect 6200 5240 6320 5250
rect 6560 5240 6600 5250
rect 7240 5240 7280 5250
rect 8000 5240 8040 5250
rect 8160 5240 8240 5250
rect 8320 5240 8360 5250
rect 8400 5240 8440 5250
rect 8920 5240 9000 5250
rect 9120 5240 9200 5250
rect 9280 5240 9400 5250
rect 9720 5240 9760 5250
rect 9840 5240 9880 5250
rect 9960 5240 9990 5250
rect 160 5230 600 5240
rect 2160 5230 2200 5240
rect 2240 5230 2400 5240
rect 2480 5230 2600 5240
rect 2640 5230 2680 5240
rect 2720 5230 2800 5240
rect 5040 5230 5080 5240
rect 5200 5230 5240 5240
rect 5560 5230 5680 5240
rect 5720 5230 5800 5240
rect 6200 5230 6320 5240
rect 6560 5230 6600 5240
rect 7240 5230 7280 5240
rect 8000 5230 8040 5240
rect 8160 5230 8240 5240
rect 8320 5230 8360 5240
rect 8400 5230 8440 5240
rect 8920 5230 9000 5240
rect 9120 5230 9200 5240
rect 9280 5230 9400 5240
rect 9720 5230 9760 5240
rect 9840 5230 9880 5240
rect 9960 5230 9990 5240
rect 160 5220 600 5230
rect 2160 5220 2200 5230
rect 2240 5220 2400 5230
rect 2480 5220 2600 5230
rect 2640 5220 2680 5230
rect 2720 5220 2800 5230
rect 5040 5220 5080 5230
rect 5200 5220 5240 5230
rect 5560 5220 5680 5230
rect 5720 5220 5800 5230
rect 6200 5220 6320 5230
rect 6560 5220 6600 5230
rect 7240 5220 7280 5230
rect 8000 5220 8040 5230
rect 8160 5220 8240 5230
rect 8320 5220 8360 5230
rect 8400 5220 8440 5230
rect 8920 5220 9000 5230
rect 9120 5220 9200 5230
rect 9280 5220 9400 5230
rect 9720 5220 9760 5230
rect 9840 5220 9880 5230
rect 9960 5220 9990 5230
rect 80 5210 600 5220
rect 2240 5210 2400 5220
rect 2440 5210 2560 5220
rect 2640 5210 2680 5220
rect 2760 5210 2880 5220
rect 3480 5210 3520 5220
rect 5040 5210 5080 5220
rect 5200 5210 5240 5220
rect 6200 5210 6280 5220
rect 6360 5210 6560 5220
rect 7200 5210 7280 5220
rect 8000 5210 8040 5220
rect 8080 5210 8120 5220
rect 8160 5210 8280 5220
rect 8320 5210 8360 5220
rect 8760 5210 8800 5220
rect 8920 5210 8960 5220
rect 9040 5210 9120 5220
rect 9160 5210 9200 5220
rect 9880 5210 9990 5220
rect 80 5200 600 5210
rect 2240 5200 2400 5210
rect 2440 5200 2560 5210
rect 2640 5200 2680 5210
rect 2760 5200 2880 5210
rect 3480 5200 3520 5210
rect 5040 5200 5080 5210
rect 5200 5200 5240 5210
rect 6200 5200 6280 5210
rect 6360 5200 6560 5210
rect 7200 5200 7280 5210
rect 8000 5200 8040 5210
rect 8080 5200 8120 5210
rect 8160 5200 8280 5210
rect 8320 5200 8360 5210
rect 8760 5200 8800 5210
rect 8920 5200 8960 5210
rect 9040 5200 9120 5210
rect 9160 5200 9200 5210
rect 9880 5200 9990 5210
rect 80 5190 600 5200
rect 2240 5190 2400 5200
rect 2440 5190 2560 5200
rect 2640 5190 2680 5200
rect 2760 5190 2880 5200
rect 3480 5190 3520 5200
rect 5040 5190 5080 5200
rect 5200 5190 5240 5200
rect 6200 5190 6280 5200
rect 6360 5190 6560 5200
rect 7200 5190 7280 5200
rect 8000 5190 8040 5200
rect 8080 5190 8120 5200
rect 8160 5190 8280 5200
rect 8320 5190 8360 5200
rect 8760 5190 8800 5200
rect 8920 5190 8960 5200
rect 9040 5190 9120 5200
rect 9160 5190 9200 5200
rect 9880 5190 9990 5200
rect 80 5180 600 5190
rect 2240 5180 2400 5190
rect 2440 5180 2560 5190
rect 2640 5180 2680 5190
rect 2760 5180 2880 5190
rect 3480 5180 3520 5190
rect 5040 5180 5080 5190
rect 5200 5180 5240 5190
rect 6200 5180 6280 5190
rect 6360 5180 6560 5190
rect 7200 5180 7280 5190
rect 8000 5180 8040 5190
rect 8080 5180 8120 5190
rect 8160 5180 8280 5190
rect 8320 5180 8360 5190
rect 8760 5180 8800 5190
rect 8920 5180 8960 5190
rect 9040 5180 9120 5190
rect 9160 5180 9200 5190
rect 9880 5180 9990 5190
rect 40 5170 600 5180
rect 2200 5170 2400 5180
rect 2440 5170 2560 5180
rect 2680 5170 2720 5180
rect 2800 5170 2840 5180
rect 5200 5170 5240 5180
rect 7280 5170 7320 5180
rect 8080 5170 8120 5180
rect 8160 5170 8200 5180
rect 8600 5170 8640 5180
rect 8680 5170 8720 5180
rect 8800 5170 8840 5180
rect 8920 5170 8960 5180
rect 9080 5170 9120 5180
rect 9400 5170 9480 5180
rect 9560 5170 9640 5180
rect 9800 5170 9840 5180
rect 9880 5170 9920 5180
rect 9960 5170 9990 5180
rect 40 5160 600 5170
rect 2200 5160 2400 5170
rect 2440 5160 2560 5170
rect 2680 5160 2720 5170
rect 2800 5160 2840 5170
rect 5200 5160 5240 5170
rect 7280 5160 7320 5170
rect 8080 5160 8120 5170
rect 8160 5160 8200 5170
rect 8600 5160 8640 5170
rect 8680 5160 8720 5170
rect 8800 5160 8840 5170
rect 8920 5160 8960 5170
rect 9080 5160 9120 5170
rect 9400 5160 9480 5170
rect 9560 5160 9640 5170
rect 9800 5160 9840 5170
rect 9880 5160 9920 5170
rect 9960 5160 9990 5170
rect 40 5150 600 5160
rect 2200 5150 2400 5160
rect 2440 5150 2560 5160
rect 2680 5150 2720 5160
rect 2800 5150 2840 5160
rect 5200 5150 5240 5160
rect 7280 5150 7320 5160
rect 8080 5150 8120 5160
rect 8160 5150 8200 5160
rect 8600 5150 8640 5160
rect 8680 5150 8720 5160
rect 8800 5150 8840 5160
rect 8920 5150 8960 5160
rect 9080 5150 9120 5160
rect 9400 5150 9480 5160
rect 9560 5150 9640 5160
rect 9800 5150 9840 5160
rect 9880 5150 9920 5160
rect 9960 5150 9990 5160
rect 40 5140 600 5150
rect 2200 5140 2400 5150
rect 2440 5140 2560 5150
rect 2680 5140 2720 5150
rect 2800 5140 2840 5150
rect 5200 5140 5240 5150
rect 7280 5140 7320 5150
rect 8080 5140 8120 5150
rect 8160 5140 8200 5150
rect 8600 5140 8640 5150
rect 8680 5140 8720 5150
rect 8800 5140 8840 5150
rect 8920 5140 8960 5150
rect 9080 5140 9120 5150
rect 9400 5140 9480 5150
rect 9560 5140 9640 5150
rect 9800 5140 9840 5150
rect 9880 5140 9920 5150
rect 9960 5140 9990 5150
rect 0 5130 520 5140
rect 2200 5130 2560 5140
rect 2640 5130 2760 5140
rect 5200 5130 5240 5140
rect 7280 5130 7320 5140
rect 8440 5130 8520 5140
rect 8680 5130 8720 5140
rect 8760 5130 8800 5140
rect 8840 5130 8880 5140
rect 8920 5130 8960 5140
rect 9280 5130 9320 5140
rect 9360 5130 9440 5140
rect 9720 5130 9800 5140
rect 0 5120 520 5130
rect 2200 5120 2560 5130
rect 2640 5120 2760 5130
rect 5200 5120 5240 5130
rect 7280 5120 7320 5130
rect 8440 5120 8520 5130
rect 8680 5120 8720 5130
rect 8760 5120 8800 5130
rect 8840 5120 8880 5130
rect 8920 5120 8960 5130
rect 9280 5120 9320 5130
rect 9360 5120 9440 5130
rect 9720 5120 9800 5130
rect 0 5110 520 5120
rect 2200 5110 2560 5120
rect 2640 5110 2760 5120
rect 5200 5110 5240 5120
rect 7280 5110 7320 5120
rect 8440 5110 8520 5120
rect 8680 5110 8720 5120
rect 8760 5110 8800 5120
rect 8840 5110 8880 5120
rect 8920 5110 8960 5120
rect 9280 5110 9320 5120
rect 9360 5110 9440 5120
rect 9720 5110 9800 5120
rect 0 5100 520 5110
rect 2200 5100 2560 5110
rect 2640 5100 2760 5110
rect 5200 5100 5240 5110
rect 7280 5100 7320 5110
rect 8440 5100 8520 5110
rect 8680 5100 8720 5110
rect 8760 5100 8800 5110
rect 8840 5100 8880 5110
rect 8920 5100 8960 5110
rect 9280 5100 9320 5110
rect 9360 5100 9440 5110
rect 9720 5100 9800 5110
rect 0 5090 440 5100
rect 2280 5090 2440 5100
rect 2480 5090 2800 5100
rect 3400 5090 3440 5100
rect 5120 5090 5160 5100
rect 5200 5090 5240 5100
rect 7280 5090 7320 5100
rect 8280 5090 8320 5100
rect 8360 5090 8400 5100
rect 8440 5090 8520 5100
rect 8680 5090 8720 5100
rect 8760 5090 8800 5100
rect 9120 5090 9200 5100
rect 9240 5090 9280 5100
rect 9360 5090 9400 5100
rect 9440 5090 9480 5100
rect 9520 5090 9560 5100
rect 0 5080 440 5090
rect 2280 5080 2440 5090
rect 2480 5080 2800 5090
rect 3400 5080 3440 5090
rect 5120 5080 5160 5090
rect 5200 5080 5240 5090
rect 7280 5080 7320 5090
rect 8280 5080 8320 5090
rect 8360 5080 8400 5090
rect 8440 5080 8520 5090
rect 8680 5080 8720 5090
rect 8760 5080 8800 5090
rect 9120 5080 9200 5090
rect 9240 5080 9280 5090
rect 9360 5080 9400 5090
rect 9440 5080 9480 5090
rect 9520 5080 9560 5090
rect 0 5070 440 5080
rect 2280 5070 2440 5080
rect 2480 5070 2800 5080
rect 3400 5070 3440 5080
rect 5120 5070 5160 5080
rect 5200 5070 5240 5080
rect 7280 5070 7320 5080
rect 8280 5070 8320 5080
rect 8360 5070 8400 5080
rect 8440 5070 8520 5080
rect 8680 5070 8720 5080
rect 8760 5070 8800 5080
rect 9120 5070 9200 5080
rect 9240 5070 9280 5080
rect 9360 5070 9400 5080
rect 9440 5070 9480 5080
rect 9520 5070 9560 5080
rect 0 5060 440 5070
rect 2280 5060 2440 5070
rect 2480 5060 2800 5070
rect 3400 5060 3440 5070
rect 5120 5060 5160 5070
rect 5200 5060 5240 5070
rect 7280 5060 7320 5070
rect 8280 5060 8320 5070
rect 8360 5060 8400 5070
rect 8440 5060 8520 5070
rect 8680 5060 8720 5070
rect 8760 5060 8800 5070
rect 9120 5060 9200 5070
rect 9240 5060 9280 5070
rect 9360 5060 9400 5070
rect 9440 5060 9480 5070
rect 9520 5060 9560 5070
rect 0 5050 360 5060
rect 2280 5050 2440 5060
rect 2520 5050 2640 5060
rect 5200 5050 5240 5060
rect 5680 5050 5800 5060
rect 7280 5050 7320 5060
rect 8240 5050 8280 5060
rect 8680 5050 8720 5060
rect 9040 5050 9080 5060
rect 9120 5050 9200 5060
rect 9400 5050 9440 5060
rect 9520 5050 9600 5060
rect 0 5040 360 5050
rect 2280 5040 2440 5050
rect 2520 5040 2640 5050
rect 5200 5040 5240 5050
rect 5680 5040 5800 5050
rect 7280 5040 7320 5050
rect 8240 5040 8280 5050
rect 8680 5040 8720 5050
rect 9040 5040 9080 5050
rect 9120 5040 9200 5050
rect 9400 5040 9440 5050
rect 9520 5040 9600 5050
rect 0 5030 360 5040
rect 2280 5030 2440 5040
rect 2520 5030 2640 5040
rect 5200 5030 5240 5040
rect 5680 5030 5800 5040
rect 7280 5030 7320 5040
rect 8240 5030 8280 5040
rect 8680 5030 8720 5040
rect 9040 5030 9080 5040
rect 9120 5030 9200 5040
rect 9400 5030 9440 5040
rect 9520 5030 9600 5040
rect 0 5020 360 5030
rect 2280 5020 2440 5030
rect 2520 5020 2640 5030
rect 5200 5020 5240 5030
rect 5680 5020 5800 5030
rect 7280 5020 7320 5030
rect 8240 5020 8280 5030
rect 8680 5020 8720 5030
rect 9040 5020 9080 5030
rect 9120 5020 9200 5030
rect 9400 5020 9440 5030
rect 9520 5020 9600 5030
rect 0 5010 360 5020
rect 2320 5010 2440 5020
rect 5160 5010 5240 5020
rect 5600 5010 5720 5020
rect 5760 5010 5800 5020
rect 6320 5010 6440 5020
rect 7280 5010 7320 5020
rect 8000 5010 8040 5020
rect 8120 5010 8200 5020
rect 8280 5010 8320 5020
rect 8360 5010 8400 5020
rect 8520 5010 8560 5020
rect 9160 5010 9200 5020
rect 9280 5010 9320 5020
rect 9400 5010 9480 5020
rect 0 5000 360 5010
rect 2320 5000 2440 5010
rect 5160 5000 5240 5010
rect 5600 5000 5720 5010
rect 5760 5000 5800 5010
rect 6320 5000 6440 5010
rect 7280 5000 7320 5010
rect 8000 5000 8040 5010
rect 8120 5000 8200 5010
rect 8280 5000 8320 5010
rect 8360 5000 8400 5010
rect 8520 5000 8560 5010
rect 9160 5000 9200 5010
rect 9280 5000 9320 5010
rect 9400 5000 9480 5010
rect 0 4990 360 5000
rect 2320 4990 2440 5000
rect 5160 4990 5240 5000
rect 5600 4990 5720 5000
rect 5760 4990 5800 5000
rect 6320 4990 6440 5000
rect 7280 4990 7320 5000
rect 8000 4990 8040 5000
rect 8120 4990 8200 5000
rect 8280 4990 8320 5000
rect 8360 4990 8400 5000
rect 8520 4990 8560 5000
rect 9160 4990 9200 5000
rect 9280 4990 9320 5000
rect 9400 4990 9480 5000
rect 0 4980 360 4990
rect 2320 4980 2440 4990
rect 5160 4980 5240 4990
rect 5600 4980 5720 4990
rect 5760 4980 5800 4990
rect 6320 4980 6440 4990
rect 7280 4980 7320 4990
rect 8000 4980 8040 4990
rect 8120 4980 8200 4990
rect 8280 4980 8320 4990
rect 8360 4980 8400 4990
rect 8520 4980 8560 4990
rect 9160 4980 9200 4990
rect 9280 4980 9320 4990
rect 9400 4980 9480 4990
rect 0 4970 240 4980
rect 280 4970 360 4980
rect 2320 4970 2480 4980
rect 3360 4970 3400 4980
rect 4360 4970 4440 4980
rect 4640 4970 4720 4980
rect 5200 4970 5240 4980
rect 5520 4970 5640 4980
rect 5760 4970 5880 4980
rect 5920 4970 5960 4980
rect 6040 4970 6200 4980
rect 6280 4970 6320 4980
rect 6400 4970 6560 4980
rect 7840 4970 7920 4980
rect 8120 4970 8160 4980
rect 8320 4970 8400 4980
rect 8640 4970 8840 4980
rect 8880 4970 8920 4980
rect 9000 4970 9080 4980
rect 9640 4970 9720 4980
rect 0 4960 240 4970
rect 280 4960 360 4970
rect 2320 4960 2480 4970
rect 3360 4960 3400 4970
rect 4360 4960 4440 4970
rect 4640 4960 4720 4970
rect 5200 4960 5240 4970
rect 5520 4960 5640 4970
rect 5760 4960 5880 4970
rect 5920 4960 5960 4970
rect 6040 4960 6200 4970
rect 6280 4960 6320 4970
rect 6400 4960 6560 4970
rect 7840 4960 7920 4970
rect 8120 4960 8160 4970
rect 8320 4960 8400 4970
rect 8640 4960 8840 4970
rect 8880 4960 8920 4970
rect 9000 4960 9080 4970
rect 9640 4960 9720 4970
rect 0 4950 240 4960
rect 280 4950 360 4960
rect 2320 4950 2480 4960
rect 3360 4950 3400 4960
rect 4360 4950 4440 4960
rect 4640 4950 4720 4960
rect 5200 4950 5240 4960
rect 5520 4950 5640 4960
rect 5760 4950 5880 4960
rect 5920 4950 5960 4960
rect 6040 4950 6200 4960
rect 6280 4950 6320 4960
rect 6400 4950 6560 4960
rect 7840 4950 7920 4960
rect 8120 4950 8160 4960
rect 8320 4950 8400 4960
rect 8640 4950 8840 4960
rect 8880 4950 8920 4960
rect 9000 4950 9080 4960
rect 9640 4950 9720 4960
rect 0 4940 240 4950
rect 280 4940 360 4950
rect 2320 4940 2480 4950
rect 3360 4940 3400 4950
rect 4360 4940 4440 4950
rect 4640 4940 4720 4950
rect 5200 4940 5240 4950
rect 5520 4940 5640 4950
rect 5760 4940 5880 4950
rect 5920 4940 5960 4950
rect 6040 4940 6200 4950
rect 6280 4940 6320 4950
rect 6400 4940 6560 4950
rect 7840 4940 7920 4950
rect 8120 4940 8160 4950
rect 8320 4940 8400 4950
rect 8640 4940 8840 4950
rect 8880 4940 8920 4950
rect 9000 4940 9080 4950
rect 9640 4940 9720 4950
rect 0 4930 80 4940
rect 2360 4930 2480 4940
rect 3360 4930 3400 4940
rect 3960 4930 4000 4940
rect 4040 4930 4200 4940
rect 4480 4930 4680 4940
rect 4800 4930 4840 4940
rect 5200 4930 5240 4940
rect 5440 4930 5560 4940
rect 5720 4930 5800 4940
rect 5960 4930 6120 4940
rect 6440 4930 6680 4940
rect 7840 4930 7960 4940
rect 8000 4930 8040 4940
rect 8120 4930 8200 4940
rect 8240 4930 8280 4940
rect 8520 4930 8560 4940
rect 8640 4930 8680 4940
rect 8760 4930 8800 4940
rect 8880 4930 9040 4940
rect 9120 4930 9160 4940
rect 9520 4930 9680 4940
rect 0 4920 80 4930
rect 2360 4920 2480 4930
rect 3360 4920 3400 4930
rect 3960 4920 4000 4930
rect 4040 4920 4200 4930
rect 4480 4920 4680 4930
rect 4800 4920 4840 4930
rect 5200 4920 5240 4930
rect 5440 4920 5560 4930
rect 5720 4920 5800 4930
rect 5960 4920 6120 4930
rect 6440 4920 6680 4930
rect 7840 4920 7960 4930
rect 8000 4920 8040 4930
rect 8120 4920 8200 4930
rect 8240 4920 8280 4930
rect 8520 4920 8560 4930
rect 8640 4920 8680 4930
rect 8760 4920 8800 4930
rect 8880 4920 9040 4930
rect 9120 4920 9160 4930
rect 9520 4920 9680 4930
rect 0 4910 80 4920
rect 2360 4910 2480 4920
rect 3360 4910 3400 4920
rect 3960 4910 4000 4920
rect 4040 4910 4200 4920
rect 4480 4910 4680 4920
rect 4800 4910 4840 4920
rect 5200 4910 5240 4920
rect 5440 4910 5560 4920
rect 5720 4910 5800 4920
rect 5960 4910 6120 4920
rect 6440 4910 6680 4920
rect 7840 4910 7960 4920
rect 8000 4910 8040 4920
rect 8120 4910 8200 4920
rect 8240 4910 8280 4920
rect 8520 4910 8560 4920
rect 8640 4910 8680 4920
rect 8760 4910 8800 4920
rect 8880 4910 9040 4920
rect 9120 4910 9160 4920
rect 9520 4910 9680 4920
rect 0 4900 80 4910
rect 2360 4900 2480 4910
rect 3360 4900 3400 4910
rect 3960 4900 4000 4910
rect 4040 4900 4200 4910
rect 4480 4900 4680 4910
rect 4800 4900 4840 4910
rect 5200 4900 5240 4910
rect 5440 4900 5560 4910
rect 5720 4900 5800 4910
rect 5960 4900 6120 4910
rect 6440 4900 6680 4910
rect 7840 4900 7960 4910
rect 8000 4900 8040 4910
rect 8120 4900 8200 4910
rect 8240 4900 8280 4910
rect 8520 4900 8560 4910
rect 8640 4900 8680 4910
rect 8760 4900 8800 4910
rect 8880 4900 9040 4910
rect 9120 4900 9160 4910
rect 9520 4900 9680 4910
rect 2360 4890 2560 4900
rect 3320 4890 3400 4900
rect 3680 4890 3760 4900
rect 3840 4890 3880 4900
rect 4840 4890 4920 4900
rect 5200 4890 5240 4900
rect 5360 4890 5520 4900
rect 5720 4890 5800 4900
rect 6480 4890 6720 4900
rect 7680 4890 7720 4900
rect 7800 4890 7840 4900
rect 8000 4890 8080 4900
rect 8520 4890 8640 4900
rect 8680 4890 8720 4900
rect 8800 4890 8840 4900
rect 8920 4890 8960 4900
rect 9080 4890 9120 4900
rect 9320 4890 9360 4900
rect 9400 4890 9480 4900
rect 9520 4890 9560 4900
rect 2360 4880 2560 4890
rect 3320 4880 3400 4890
rect 3680 4880 3760 4890
rect 3840 4880 3880 4890
rect 4840 4880 4920 4890
rect 5200 4880 5240 4890
rect 5360 4880 5520 4890
rect 5720 4880 5800 4890
rect 6480 4880 6720 4890
rect 7680 4880 7720 4890
rect 7800 4880 7840 4890
rect 8000 4880 8080 4890
rect 8520 4880 8640 4890
rect 8680 4880 8720 4890
rect 8800 4880 8840 4890
rect 8920 4880 8960 4890
rect 9080 4880 9120 4890
rect 9320 4880 9360 4890
rect 9400 4880 9480 4890
rect 9520 4880 9560 4890
rect 2360 4870 2560 4880
rect 3320 4870 3400 4880
rect 3680 4870 3760 4880
rect 3840 4870 3880 4880
rect 4840 4870 4920 4880
rect 5200 4870 5240 4880
rect 5360 4870 5520 4880
rect 5720 4870 5800 4880
rect 6480 4870 6720 4880
rect 7680 4870 7720 4880
rect 7800 4870 7840 4880
rect 8000 4870 8080 4880
rect 8520 4870 8640 4880
rect 8680 4870 8720 4880
rect 8800 4870 8840 4880
rect 8920 4870 8960 4880
rect 9080 4870 9120 4880
rect 9320 4870 9360 4880
rect 9400 4870 9480 4880
rect 9520 4870 9560 4880
rect 2360 4860 2560 4870
rect 3320 4860 3400 4870
rect 3680 4860 3760 4870
rect 3840 4860 3880 4870
rect 4840 4860 4920 4870
rect 5200 4860 5240 4870
rect 5360 4860 5520 4870
rect 5720 4860 5800 4870
rect 6480 4860 6720 4870
rect 7680 4860 7720 4870
rect 7800 4860 7840 4870
rect 8000 4860 8080 4870
rect 8520 4860 8640 4870
rect 8680 4860 8720 4870
rect 8800 4860 8840 4870
rect 8920 4860 8960 4870
rect 9080 4860 9120 4870
rect 9320 4860 9360 4870
rect 9400 4860 9480 4870
rect 9520 4860 9560 4870
rect 2400 4850 2640 4860
rect 3360 4850 3400 4860
rect 3640 4850 3680 4860
rect 4960 4850 5000 4860
rect 5160 4850 5240 4860
rect 5360 4850 5480 4860
rect 5720 4850 5840 4860
rect 6520 4850 6720 4860
rect 7320 4850 7360 4860
rect 7680 4850 7720 4860
rect 7800 4850 7840 4860
rect 7920 4850 7960 4860
rect 8640 4850 8720 4860
rect 8760 4850 8800 4860
rect 9400 4850 9440 4860
rect 9680 4850 9760 4860
rect 2400 4840 2640 4850
rect 3360 4840 3400 4850
rect 3640 4840 3680 4850
rect 4960 4840 5000 4850
rect 5160 4840 5240 4850
rect 5360 4840 5480 4850
rect 5720 4840 5840 4850
rect 6520 4840 6720 4850
rect 7320 4840 7360 4850
rect 7680 4840 7720 4850
rect 7800 4840 7840 4850
rect 7920 4840 7960 4850
rect 8640 4840 8720 4850
rect 8760 4840 8800 4850
rect 9400 4840 9440 4850
rect 9680 4840 9760 4850
rect 2400 4830 2640 4840
rect 3360 4830 3400 4840
rect 3640 4830 3680 4840
rect 4960 4830 5000 4840
rect 5160 4830 5240 4840
rect 5360 4830 5480 4840
rect 5720 4830 5840 4840
rect 6520 4830 6720 4840
rect 7320 4830 7360 4840
rect 7680 4830 7720 4840
rect 7800 4830 7840 4840
rect 7920 4830 7960 4840
rect 8640 4830 8720 4840
rect 8760 4830 8800 4840
rect 9400 4830 9440 4840
rect 9680 4830 9760 4840
rect 2400 4820 2640 4830
rect 3360 4820 3400 4830
rect 3640 4820 3680 4830
rect 4960 4820 5000 4830
rect 5160 4820 5240 4830
rect 5360 4820 5480 4830
rect 5720 4820 5840 4830
rect 6520 4820 6720 4830
rect 7320 4820 7360 4830
rect 7680 4820 7720 4830
rect 7800 4820 7840 4830
rect 7920 4820 7960 4830
rect 8640 4820 8720 4830
rect 8760 4820 8800 4830
rect 9400 4820 9440 4830
rect 9680 4820 9760 4830
rect 2400 4810 2680 4820
rect 3360 4810 3400 4820
rect 3600 4810 3640 4820
rect 5160 4810 5200 4820
rect 5360 4810 5440 4820
rect 5680 4810 5960 4820
rect 6560 4810 6720 4820
rect 7320 4810 7360 4820
rect 7720 4810 7760 4820
rect 8320 4810 8360 4820
rect 8480 4810 8520 4820
rect 8640 4810 8720 4820
rect 9000 4810 9040 4820
rect 9320 4810 9360 4820
rect 9400 4810 9440 4820
rect 9560 4810 9600 4820
rect 2400 4800 2680 4810
rect 3360 4800 3400 4810
rect 3600 4800 3640 4810
rect 5160 4800 5200 4810
rect 5360 4800 5440 4810
rect 5680 4800 5960 4810
rect 6560 4800 6720 4810
rect 7320 4800 7360 4810
rect 7720 4800 7760 4810
rect 8320 4800 8360 4810
rect 8480 4800 8520 4810
rect 8640 4800 8720 4810
rect 9000 4800 9040 4810
rect 9320 4800 9360 4810
rect 9400 4800 9440 4810
rect 9560 4800 9600 4810
rect 2400 4790 2680 4800
rect 3360 4790 3400 4800
rect 3600 4790 3640 4800
rect 5160 4790 5200 4800
rect 5360 4790 5440 4800
rect 5680 4790 5960 4800
rect 6560 4790 6720 4800
rect 7320 4790 7360 4800
rect 7720 4790 7760 4800
rect 8320 4790 8360 4800
rect 8480 4790 8520 4800
rect 8640 4790 8720 4800
rect 9000 4790 9040 4800
rect 9320 4790 9360 4800
rect 9400 4790 9440 4800
rect 9560 4790 9600 4800
rect 2400 4780 2680 4790
rect 3360 4780 3400 4790
rect 3600 4780 3640 4790
rect 5160 4780 5200 4790
rect 5360 4780 5440 4790
rect 5680 4780 5960 4790
rect 6560 4780 6720 4790
rect 7320 4780 7360 4790
rect 7720 4780 7760 4790
rect 8320 4780 8360 4790
rect 8480 4780 8520 4790
rect 8640 4780 8720 4790
rect 9000 4780 9040 4790
rect 9320 4780 9360 4790
rect 9400 4780 9440 4790
rect 9560 4780 9600 4790
rect 2480 4770 2720 4780
rect 3240 4770 3280 4780
rect 3520 4770 3600 4780
rect 5360 4770 5400 4780
rect 5640 4770 5760 4780
rect 5920 4770 6000 4780
rect 6640 4770 6720 4780
rect 8080 4770 8120 4780
rect 8800 4770 8880 4780
rect 9280 4770 9360 4780
rect 2480 4760 2720 4770
rect 3240 4760 3280 4770
rect 3520 4760 3600 4770
rect 5360 4760 5400 4770
rect 5640 4760 5760 4770
rect 5920 4760 6000 4770
rect 6640 4760 6720 4770
rect 8080 4760 8120 4770
rect 8800 4760 8880 4770
rect 9280 4760 9360 4770
rect 2480 4750 2720 4760
rect 3240 4750 3280 4760
rect 3520 4750 3600 4760
rect 5360 4750 5400 4760
rect 5640 4750 5760 4760
rect 5920 4750 6000 4760
rect 6640 4750 6720 4760
rect 8080 4750 8120 4760
rect 8800 4750 8880 4760
rect 9280 4750 9360 4760
rect 2480 4740 2720 4750
rect 3240 4740 3280 4750
rect 3520 4740 3600 4750
rect 5360 4740 5400 4750
rect 5640 4740 5760 4750
rect 5920 4740 6000 4750
rect 6640 4740 6720 4750
rect 8080 4740 8120 4750
rect 8800 4740 8880 4750
rect 9280 4740 9360 4750
rect 2560 4730 2720 4740
rect 3480 4730 3520 4740
rect 5120 4730 5160 4740
rect 5320 4730 5400 4740
rect 5640 4730 5760 4740
rect 5920 4730 6040 4740
rect 6240 4730 6320 4740
rect 6640 4730 6760 4740
rect 7760 4730 7800 4740
rect 7840 4730 7960 4740
rect 8040 4730 8080 4740
rect 8120 4730 8200 4740
rect 8240 4730 8320 4740
rect 8800 4730 8880 4740
rect 2560 4720 2720 4730
rect 3480 4720 3520 4730
rect 5120 4720 5160 4730
rect 5320 4720 5400 4730
rect 5640 4720 5760 4730
rect 5920 4720 6040 4730
rect 6240 4720 6320 4730
rect 6640 4720 6760 4730
rect 7760 4720 7800 4730
rect 7840 4720 7960 4730
rect 8040 4720 8080 4730
rect 8120 4720 8200 4730
rect 8240 4720 8320 4730
rect 8800 4720 8880 4730
rect 2560 4710 2720 4720
rect 3480 4710 3520 4720
rect 5120 4710 5160 4720
rect 5320 4710 5400 4720
rect 5640 4710 5760 4720
rect 5920 4710 6040 4720
rect 6240 4710 6320 4720
rect 6640 4710 6760 4720
rect 7760 4710 7800 4720
rect 7840 4710 7960 4720
rect 8040 4710 8080 4720
rect 8120 4710 8200 4720
rect 8240 4710 8320 4720
rect 8800 4710 8880 4720
rect 2560 4700 2720 4710
rect 3480 4700 3520 4710
rect 5120 4700 5160 4710
rect 5320 4700 5400 4710
rect 5640 4700 5760 4710
rect 5920 4700 6040 4710
rect 6240 4700 6320 4710
rect 6640 4700 6760 4710
rect 7760 4700 7800 4710
rect 7840 4700 7960 4710
rect 8040 4700 8080 4710
rect 8120 4700 8200 4710
rect 8240 4700 8320 4710
rect 8800 4700 8880 4710
rect 3360 4690 3400 4700
rect 5160 4690 5200 4700
rect 5320 4690 5400 4700
rect 5760 4690 6320 4700
rect 6640 4690 6760 4700
rect 7360 4690 7400 4700
rect 7600 4690 7680 4700
rect 7760 4690 7800 4700
rect 7840 4690 7880 4700
rect 8040 4690 8080 4700
rect 8160 4690 8200 4700
rect 8560 4690 8600 4700
rect 8800 4690 8840 4700
rect 8880 4690 9000 4700
rect 9800 4690 9840 4700
rect 3360 4680 3400 4690
rect 5160 4680 5200 4690
rect 5320 4680 5400 4690
rect 5760 4680 6320 4690
rect 6640 4680 6760 4690
rect 7360 4680 7400 4690
rect 7600 4680 7680 4690
rect 7760 4680 7800 4690
rect 7840 4680 7880 4690
rect 8040 4680 8080 4690
rect 8160 4680 8200 4690
rect 8560 4680 8600 4690
rect 8800 4680 8840 4690
rect 8880 4680 9000 4690
rect 9800 4680 9840 4690
rect 3360 4670 3400 4680
rect 5160 4670 5200 4680
rect 5320 4670 5400 4680
rect 5760 4670 6320 4680
rect 6640 4670 6760 4680
rect 7360 4670 7400 4680
rect 7600 4670 7680 4680
rect 7760 4670 7800 4680
rect 7840 4670 7880 4680
rect 8040 4670 8080 4680
rect 8160 4670 8200 4680
rect 8560 4670 8600 4680
rect 8800 4670 8840 4680
rect 8880 4670 9000 4680
rect 9800 4670 9840 4680
rect 3360 4660 3400 4670
rect 5160 4660 5200 4670
rect 5320 4660 5400 4670
rect 5760 4660 6320 4670
rect 6640 4660 6760 4670
rect 7360 4660 7400 4670
rect 7600 4660 7680 4670
rect 7760 4660 7800 4670
rect 7840 4660 7880 4670
rect 8040 4660 8080 4670
rect 8160 4660 8200 4670
rect 8560 4660 8600 4670
rect 8800 4660 8840 4670
rect 8880 4660 9000 4670
rect 9800 4660 9840 4670
rect 3320 4650 3400 4660
rect 3440 4650 3480 4660
rect 5280 4650 5400 4660
rect 6640 4650 6760 4660
rect 7360 4650 7400 4660
rect 7480 4650 7520 4660
rect 7560 4650 7600 4660
rect 7640 4650 7680 4660
rect 7720 4650 7760 4660
rect 7800 4650 7840 4660
rect 7920 4650 8080 4660
rect 8320 4650 8360 4660
rect 8480 4650 8520 4660
rect 8600 4650 8640 4660
rect 8840 4650 8920 4660
rect 8960 4650 9000 4660
rect 9240 4650 9280 4660
rect 9760 4650 9800 4660
rect 3320 4640 3400 4650
rect 3440 4640 3480 4650
rect 5280 4640 5400 4650
rect 6640 4640 6760 4650
rect 7360 4640 7400 4650
rect 7480 4640 7520 4650
rect 7560 4640 7600 4650
rect 7640 4640 7680 4650
rect 7720 4640 7760 4650
rect 7800 4640 7840 4650
rect 7920 4640 8080 4650
rect 8320 4640 8360 4650
rect 8480 4640 8520 4650
rect 8600 4640 8640 4650
rect 8840 4640 8920 4650
rect 8960 4640 9000 4650
rect 9240 4640 9280 4650
rect 9760 4640 9800 4650
rect 3320 4630 3400 4640
rect 3440 4630 3480 4640
rect 5280 4630 5400 4640
rect 6640 4630 6760 4640
rect 7360 4630 7400 4640
rect 7480 4630 7520 4640
rect 7560 4630 7600 4640
rect 7640 4630 7680 4640
rect 7720 4630 7760 4640
rect 7800 4630 7840 4640
rect 7920 4630 8080 4640
rect 8320 4630 8360 4640
rect 8480 4630 8520 4640
rect 8600 4630 8640 4640
rect 8840 4630 8920 4640
rect 8960 4630 9000 4640
rect 9240 4630 9280 4640
rect 9760 4630 9800 4640
rect 3320 4620 3400 4630
rect 3440 4620 3480 4630
rect 5280 4620 5400 4630
rect 6640 4620 6760 4630
rect 7360 4620 7400 4630
rect 7480 4620 7520 4630
rect 7560 4620 7600 4630
rect 7640 4620 7680 4630
rect 7720 4620 7760 4630
rect 7800 4620 7840 4630
rect 7920 4620 8080 4630
rect 8320 4620 8360 4630
rect 8480 4620 8520 4630
rect 8600 4620 8640 4630
rect 8840 4620 8920 4630
rect 8960 4620 9000 4630
rect 9240 4620 9280 4630
rect 9760 4620 9800 4630
rect 3280 4610 3400 4620
rect 5280 4610 5400 4620
rect 5920 4610 6000 4620
rect 6600 4610 6720 4620
rect 7360 4610 7400 4620
rect 7520 4610 7680 4620
rect 7720 4610 7760 4620
rect 7880 4610 7960 4620
rect 8160 4610 8240 4620
rect 8320 4610 8400 4620
rect 8480 4610 8520 4620
rect 8560 4610 8680 4620
rect 8960 4610 9000 4620
rect 9720 4610 9760 4620
rect 3280 4600 3400 4610
rect 5280 4600 5400 4610
rect 5920 4600 6000 4610
rect 6600 4600 6720 4610
rect 7360 4600 7400 4610
rect 7520 4600 7680 4610
rect 7720 4600 7760 4610
rect 7880 4600 7960 4610
rect 8160 4600 8240 4610
rect 8320 4600 8400 4610
rect 8480 4600 8520 4610
rect 8560 4600 8680 4610
rect 8960 4600 9000 4610
rect 9720 4600 9760 4610
rect 3280 4590 3400 4600
rect 5280 4590 5400 4600
rect 5920 4590 6000 4600
rect 6600 4590 6720 4600
rect 7360 4590 7400 4600
rect 7520 4590 7680 4600
rect 7720 4590 7760 4600
rect 7880 4590 7960 4600
rect 8160 4590 8240 4600
rect 8320 4590 8400 4600
rect 8480 4590 8520 4600
rect 8560 4590 8680 4600
rect 8960 4590 9000 4600
rect 9720 4590 9760 4600
rect 3280 4580 3400 4590
rect 5280 4580 5400 4590
rect 5920 4580 6000 4590
rect 6600 4580 6720 4590
rect 7360 4580 7400 4590
rect 7520 4580 7680 4590
rect 7720 4580 7760 4590
rect 7880 4580 7960 4590
rect 8160 4580 8240 4590
rect 8320 4580 8400 4590
rect 8480 4580 8520 4590
rect 8560 4580 8680 4590
rect 8960 4580 9000 4590
rect 9720 4580 9760 4590
rect 3240 4570 3280 4580
rect 3320 4570 3360 4580
rect 5280 4570 5440 4580
rect 5600 4570 5640 4580
rect 5800 4570 5880 4580
rect 6000 4570 6160 4580
rect 6560 4570 6720 4580
rect 7320 4570 7360 4580
rect 7480 4570 7560 4580
rect 7600 4570 7640 4580
rect 7680 4570 7720 4580
rect 8080 4570 8120 4580
rect 8360 4570 8400 4580
rect 8480 4570 8520 4580
rect 9680 4570 9720 4580
rect 9960 4570 9990 4580
rect 3240 4560 3280 4570
rect 3320 4560 3360 4570
rect 5280 4560 5440 4570
rect 5600 4560 5640 4570
rect 5800 4560 5880 4570
rect 6000 4560 6160 4570
rect 6560 4560 6720 4570
rect 7320 4560 7360 4570
rect 7480 4560 7560 4570
rect 7600 4560 7640 4570
rect 7680 4560 7720 4570
rect 8080 4560 8120 4570
rect 8360 4560 8400 4570
rect 8480 4560 8520 4570
rect 9680 4560 9720 4570
rect 9960 4560 9990 4570
rect 3240 4550 3280 4560
rect 3320 4550 3360 4560
rect 5280 4550 5440 4560
rect 5600 4550 5640 4560
rect 5800 4550 5880 4560
rect 6000 4550 6160 4560
rect 6560 4550 6720 4560
rect 7320 4550 7360 4560
rect 7480 4550 7560 4560
rect 7600 4550 7640 4560
rect 7680 4550 7720 4560
rect 8080 4550 8120 4560
rect 8360 4550 8400 4560
rect 8480 4550 8520 4560
rect 9680 4550 9720 4560
rect 9960 4550 9990 4560
rect 3240 4540 3280 4550
rect 3320 4540 3360 4550
rect 5280 4540 5440 4550
rect 5600 4540 5640 4550
rect 5800 4540 5880 4550
rect 6000 4540 6160 4550
rect 6560 4540 6720 4550
rect 7320 4540 7360 4550
rect 7480 4540 7560 4550
rect 7600 4540 7640 4550
rect 7680 4540 7720 4550
rect 8080 4540 8120 4550
rect 8360 4540 8400 4550
rect 8480 4540 8520 4550
rect 9680 4540 9720 4550
rect 9960 4540 9990 4550
rect 3240 4530 3280 4540
rect 3400 4530 3440 4540
rect 5280 4530 5480 4540
rect 5600 4530 5680 4540
rect 5840 4530 5880 4540
rect 6160 4530 6240 4540
rect 6520 4530 6720 4540
rect 7320 4530 7400 4540
rect 7480 4530 7560 4540
rect 7880 4530 7920 4540
rect 7960 4530 8040 4540
rect 8120 4530 8160 4540
rect 8200 4530 8240 4540
rect 8280 4530 8320 4540
rect 8480 4530 8520 4540
rect 8920 4530 8960 4540
rect 9200 4530 9240 4540
rect 9640 4530 9680 4540
rect 3240 4520 3280 4530
rect 3400 4520 3440 4530
rect 5280 4520 5480 4530
rect 5600 4520 5680 4530
rect 5840 4520 5880 4530
rect 6160 4520 6240 4530
rect 6520 4520 6720 4530
rect 7320 4520 7400 4530
rect 7480 4520 7560 4530
rect 7880 4520 7920 4530
rect 7960 4520 8040 4530
rect 8120 4520 8160 4530
rect 8200 4520 8240 4530
rect 8280 4520 8320 4530
rect 8480 4520 8520 4530
rect 8920 4520 8960 4530
rect 9200 4520 9240 4530
rect 9640 4520 9680 4530
rect 3240 4510 3280 4520
rect 3400 4510 3440 4520
rect 5280 4510 5480 4520
rect 5600 4510 5680 4520
rect 5840 4510 5880 4520
rect 6160 4510 6240 4520
rect 6520 4510 6720 4520
rect 7320 4510 7400 4520
rect 7480 4510 7560 4520
rect 7880 4510 7920 4520
rect 7960 4510 8040 4520
rect 8120 4510 8160 4520
rect 8200 4510 8240 4520
rect 8280 4510 8320 4520
rect 8480 4510 8520 4520
rect 8920 4510 8960 4520
rect 9200 4510 9240 4520
rect 9640 4510 9680 4520
rect 3240 4500 3280 4510
rect 3400 4500 3440 4510
rect 5280 4500 5480 4510
rect 5600 4500 5680 4510
rect 5840 4500 5880 4510
rect 6160 4500 6240 4510
rect 6520 4500 6720 4510
rect 7320 4500 7400 4510
rect 7480 4500 7560 4510
rect 7880 4500 7920 4510
rect 7960 4500 8040 4510
rect 8120 4500 8160 4510
rect 8200 4500 8240 4510
rect 8280 4500 8320 4510
rect 8480 4500 8520 4510
rect 8920 4500 8960 4510
rect 9200 4500 9240 4510
rect 9640 4500 9680 4510
rect 3000 4490 3040 4500
rect 5280 4490 5320 4500
rect 5360 4490 5480 4500
rect 5600 4490 5720 4500
rect 5800 4490 5920 4500
rect 6160 4490 6200 4500
rect 6520 4490 6720 4500
rect 7320 4490 7360 4500
rect 7400 4490 7440 4500
rect 8120 4490 8280 4500
rect 9200 4490 9240 4500
rect 9600 4490 9640 4500
rect 3000 4480 3040 4490
rect 5280 4480 5320 4490
rect 5360 4480 5480 4490
rect 5600 4480 5720 4490
rect 5800 4480 5920 4490
rect 6160 4480 6200 4490
rect 6520 4480 6720 4490
rect 7320 4480 7360 4490
rect 7400 4480 7440 4490
rect 8120 4480 8280 4490
rect 9200 4480 9240 4490
rect 9600 4480 9640 4490
rect 3000 4470 3040 4480
rect 5280 4470 5320 4480
rect 5360 4470 5480 4480
rect 5600 4470 5720 4480
rect 5800 4470 5920 4480
rect 6160 4470 6200 4480
rect 6520 4470 6720 4480
rect 7320 4470 7360 4480
rect 7400 4470 7440 4480
rect 8120 4470 8280 4480
rect 9200 4470 9240 4480
rect 9600 4470 9640 4480
rect 3000 4460 3040 4470
rect 5280 4460 5320 4470
rect 5360 4460 5480 4470
rect 5600 4460 5720 4470
rect 5800 4460 5920 4470
rect 6160 4460 6200 4470
rect 6520 4460 6720 4470
rect 7320 4460 7360 4470
rect 7400 4460 7440 4470
rect 8120 4460 8280 4470
rect 9200 4460 9240 4470
rect 9600 4460 9640 4470
rect 3000 4450 3040 4460
rect 3280 4450 3320 4460
rect 3360 4450 3400 4460
rect 5320 4450 5520 4460
rect 5600 4450 5760 4460
rect 5800 4450 6120 4460
rect 6520 4450 6680 4460
rect 7880 4450 7920 4460
rect 8080 4450 8160 4460
rect 8200 4450 8240 4460
rect 8880 4450 8920 4460
rect 9560 4450 9600 4460
rect 9840 4450 9880 4460
rect 3000 4440 3040 4450
rect 3280 4440 3320 4450
rect 3360 4440 3400 4450
rect 5320 4440 5520 4450
rect 5600 4440 5760 4450
rect 5800 4440 6120 4450
rect 6520 4440 6680 4450
rect 7880 4440 7920 4450
rect 8080 4440 8160 4450
rect 8200 4440 8240 4450
rect 8880 4440 8920 4450
rect 9560 4440 9600 4450
rect 9840 4440 9880 4450
rect 3000 4430 3040 4440
rect 3280 4430 3320 4440
rect 3360 4430 3400 4440
rect 5320 4430 5520 4440
rect 5600 4430 5760 4440
rect 5800 4430 6120 4440
rect 6520 4430 6680 4440
rect 7880 4430 7920 4440
rect 8080 4430 8160 4440
rect 8200 4430 8240 4440
rect 8880 4430 8920 4440
rect 9560 4430 9600 4440
rect 9840 4430 9880 4440
rect 3000 4420 3040 4430
rect 3280 4420 3320 4430
rect 3360 4420 3400 4430
rect 5320 4420 5520 4430
rect 5600 4420 5760 4430
rect 5800 4420 6120 4430
rect 6520 4420 6680 4430
rect 7880 4420 7920 4430
rect 8080 4420 8160 4430
rect 8200 4420 8240 4430
rect 8880 4420 8920 4430
rect 9560 4420 9600 4430
rect 9840 4420 9880 4430
rect 2960 4410 3000 4420
rect 3240 4410 3280 4420
rect 5320 4410 5400 4420
rect 5440 4410 5520 4420
rect 5560 4410 6000 4420
rect 6520 4410 6680 4420
rect 7320 4410 7360 4420
rect 7400 4410 7440 4420
rect 7800 4410 7840 4420
rect 8840 4410 8880 4420
rect 9520 4410 9560 4420
rect 2960 4400 3000 4410
rect 3240 4400 3280 4410
rect 5320 4400 5400 4410
rect 5440 4400 5520 4410
rect 5560 4400 6000 4410
rect 6520 4400 6680 4410
rect 7320 4400 7360 4410
rect 7400 4400 7440 4410
rect 7800 4400 7840 4410
rect 8840 4400 8880 4410
rect 9520 4400 9560 4410
rect 2960 4390 3000 4400
rect 3240 4390 3280 4400
rect 5320 4390 5400 4400
rect 5440 4390 5520 4400
rect 5560 4390 6000 4400
rect 6520 4390 6680 4400
rect 7320 4390 7360 4400
rect 7400 4390 7440 4400
rect 7800 4390 7840 4400
rect 8840 4390 8880 4400
rect 9520 4390 9560 4400
rect 2960 4380 3000 4390
rect 3240 4380 3280 4390
rect 5320 4380 5400 4390
rect 5440 4380 5520 4390
rect 5560 4380 6000 4390
rect 6520 4380 6680 4390
rect 7320 4380 7360 4390
rect 7400 4380 7440 4390
rect 7800 4380 7840 4390
rect 8840 4380 8880 4390
rect 9520 4380 9560 4390
rect 2960 4370 3000 4380
rect 3320 4370 3360 4380
rect 4600 4370 4760 4380
rect 5320 4370 5400 4380
rect 5480 4370 5800 4380
rect 5920 4370 5960 4380
rect 6480 4370 6680 4380
rect 7320 4370 7400 4380
rect 8680 4370 8720 4380
rect 8840 4370 8880 4380
rect 9160 4370 9200 4380
rect 9480 4370 9520 4380
rect 2960 4360 3000 4370
rect 3320 4360 3360 4370
rect 4600 4360 4760 4370
rect 5320 4360 5400 4370
rect 5480 4360 5800 4370
rect 5920 4360 5960 4370
rect 6480 4360 6680 4370
rect 7320 4360 7400 4370
rect 8680 4360 8720 4370
rect 8840 4360 8880 4370
rect 9160 4360 9200 4370
rect 9480 4360 9520 4370
rect 2960 4350 3000 4360
rect 3320 4350 3360 4360
rect 4600 4350 4760 4360
rect 5320 4350 5400 4360
rect 5480 4350 5800 4360
rect 5920 4350 5960 4360
rect 6480 4350 6680 4360
rect 7320 4350 7400 4360
rect 8680 4350 8720 4360
rect 8840 4350 8880 4360
rect 9160 4350 9200 4360
rect 9480 4350 9520 4360
rect 2960 4340 3000 4350
rect 3320 4340 3360 4350
rect 4600 4340 4760 4350
rect 5320 4340 5400 4350
rect 5480 4340 5800 4350
rect 5920 4340 5960 4350
rect 6480 4340 6680 4350
rect 7320 4340 7400 4350
rect 8680 4340 8720 4350
rect 8840 4340 8880 4350
rect 9160 4340 9200 4350
rect 9480 4340 9520 4350
rect 2920 4330 3000 4340
rect 4600 4330 4680 4340
rect 4760 4330 4880 4340
rect 5400 4330 5440 4340
rect 5480 4330 6120 4340
rect 6480 4330 6680 4340
rect 7280 4330 7360 4340
rect 8440 4330 8520 4340
rect 8680 4330 8760 4340
rect 9160 4330 9200 4340
rect 9440 4330 9480 4340
rect 9840 4330 9990 4340
rect 2920 4320 3000 4330
rect 4600 4320 4680 4330
rect 4760 4320 4880 4330
rect 5400 4320 5440 4330
rect 5480 4320 6120 4330
rect 6480 4320 6680 4330
rect 7280 4320 7360 4330
rect 8440 4320 8520 4330
rect 8680 4320 8760 4330
rect 9160 4320 9200 4330
rect 9440 4320 9480 4330
rect 9840 4320 9990 4330
rect 2920 4310 3000 4320
rect 4600 4310 4680 4320
rect 4760 4310 4880 4320
rect 5400 4310 5440 4320
rect 5480 4310 6120 4320
rect 6480 4310 6680 4320
rect 7280 4310 7360 4320
rect 8440 4310 8520 4320
rect 8680 4310 8760 4320
rect 9160 4310 9200 4320
rect 9440 4310 9480 4320
rect 9840 4310 9990 4320
rect 2920 4300 3000 4310
rect 4600 4300 4680 4310
rect 4760 4300 4880 4310
rect 5400 4300 5440 4310
rect 5480 4300 6120 4310
rect 6480 4300 6680 4310
rect 7280 4300 7360 4310
rect 8440 4300 8520 4310
rect 8680 4300 8760 4310
rect 9160 4300 9200 4310
rect 9440 4300 9480 4310
rect 9840 4300 9990 4310
rect 3200 4290 3240 4300
rect 4560 4290 4640 4300
rect 4840 4290 4920 4300
rect 5520 4290 5960 4300
rect 6440 4290 6640 4300
rect 7120 4290 7200 4300
rect 8840 4290 8880 4300
rect 9160 4290 9200 4300
rect 9400 4290 9440 4300
rect 9800 4290 9960 4300
rect 3200 4280 3240 4290
rect 4560 4280 4640 4290
rect 4840 4280 4920 4290
rect 5520 4280 5960 4290
rect 6440 4280 6640 4290
rect 7120 4280 7200 4290
rect 8840 4280 8880 4290
rect 9160 4280 9200 4290
rect 9400 4280 9440 4290
rect 9800 4280 9960 4290
rect 3200 4270 3240 4280
rect 4560 4270 4640 4280
rect 4840 4270 4920 4280
rect 5520 4270 5960 4280
rect 6440 4270 6640 4280
rect 7120 4270 7200 4280
rect 8840 4270 8880 4280
rect 9160 4270 9200 4280
rect 9400 4270 9440 4280
rect 9800 4270 9960 4280
rect 3200 4260 3240 4270
rect 4560 4260 4640 4270
rect 4840 4260 4920 4270
rect 5520 4260 5960 4270
rect 6440 4260 6640 4270
rect 7120 4260 7200 4270
rect 8840 4260 8880 4270
rect 9160 4260 9200 4270
rect 9400 4260 9440 4270
rect 9800 4260 9960 4270
rect 4160 4250 4320 4260
rect 4520 4250 4600 4260
rect 4840 4250 4920 4260
rect 5360 4250 5400 4260
rect 5520 4250 5640 4260
rect 5720 4250 6000 4260
rect 6280 4250 6320 4260
rect 6360 4250 6520 4260
rect 6560 4250 6680 4260
rect 7080 4250 7120 4260
rect 9160 4250 9200 4260
rect 9840 4250 9990 4260
rect 4160 4240 4320 4250
rect 4520 4240 4600 4250
rect 4840 4240 4920 4250
rect 5360 4240 5400 4250
rect 5520 4240 5640 4250
rect 5720 4240 6000 4250
rect 6280 4240 6320 4250
rect 6360 4240 6520 4250
rect 6560 4240 6680 4250
rect 7080 4240 7120 4250
rect 9160 4240 9200 4250
rect 9840 4240 9990 4250
rect 4160 4230 4320 4240
rect 4520 4230 4600 4240
rect 4840 4230 4920 4240
rect 5360 4230 5400 4240
rect 5520 4230 5640 4240
rect 5720 4230 6000 4240
rect 6280 4230 6320 4240
rect 6360 4230 6520 4240
rect 6560 4230 6680 4240
rect 7080 4230 7120 4240
rect 9160 4230 9200 4240
rect 9840 4230 9990 4240
rect 4160 4220 4320 4230
rect 4520 4220 4600 4230
rect 4840 4220 4920 4230
rect 5360 4220 5400 4230
rect 5520 4220 5640 4230
rect 5720 4220 6000 4230
rect 6280 4220 6320 4230
rect 6360 4220 6520 4230
rect 6560 4220 6680 4230
rect 7080 4220 7120 4230
rect 9160 4220 9200 4230
rect 9840 4220 9990 4230
rect 4160 4210 4240 4220
rect 4320 4210 4360 4220
rect 4480 4210 4960 4220
rect 5560 4210 5640 4220
rect 5920 4210 6480 4220
rect 6560 4210 6680 4220
rect 7280 4210 7360 4220
rect 7440 4210 7480 4220
rect 9160 4210 9280 4220
rect 9680 4210 9760 4220
rect 9840 4210 9920 4220
rect 9960 4210 9990 4220
rect 4160 4200 4240 4210
rect 4320 4200 4360 4210
rect 4480 4200 4960 4210
rect 5560 4200 5640 4210
rect 5920 4200 6480 4210
rect 6560 4200 6680 4210
rect 7280 4200 7360 4210
rect 7440 4200 7480 4210
rect 9160 4200 9280 4210
rect 9680 4200 9760 4210
rect 9840 4200 9920 4210
rect 9960 4200 9990 4210
rect 4160 4190 4240 4200
rect 4320 4190 4360 4200
rect 4480 4190 4960 4200
rect 5560 4190 5640 4200
rect 5920 4190 6480 4200
rect 6560 4190 6680 4200
rect 7280 4190 7360 4200
rect 7440 4190 7480 4200
rect 9160 4190 9280 4200
rect 9680 4190 9760 4200
rect 9840 4190 9920 4200
rect 9960 4190 9990 4200
rect 4160 4180 4240 4190
rect 4320 4180 4360 4190
rect 4480 4180 4960 4190
rect 5560 4180 5640 4190
rect 5920 4180 6480 4190
rect 6560 4180 6680 4190
rect 7280 4180 7360 4190
rect 7440 4180 7480 4190
rect 9160 4180 9280 4190
rect 9680 4180 9760 4190
rect 9840 4180 9920 4190
rect 9960 4180 9990 4190
rect 4120 4170 4200 4180
rect 4360 4170 4640 4180
rect 4720 4170 5000 4180
rect 5600 4170 5680 4180
rect 5920 4170 6440 4180
rect 6520 4170 6680 4180
rect 7440 4170 7480 4180
rect 8800 4170 8840 4180
rect 9640 4170 9680 4180
rect 9800 4170 9840 4180
rect 9880 4170 9920 4180
rect 9960 4170 9990 4180
rect 4120 4160 4200 4170
rect 4360 4160 4640 4170
rect 4720 4160 5000 4170
rect 5600 4160 5680 4170
rect 5920 4160 6440 4170
rect 6520 4160 6680 4170
rect 7440 4160 7480 4170
rect 8800 4160 8840 4170
rect 9640 4160 9680 4170
rect 9800 4160 9840 4170
rect 9880 4160 9920 4170
rect 9960 4160 9990 4170
rect 4120 4150 4200 4160
rect 4360 4150 4640 4160
rect 4720 4150 5000 4160
rect 5600 4150 5680 4160
rect 5920 4150 6440 4160
rect 6520 4150 6680 4160
rect 7440 4150 7480 4160
rect 8800 4150 8840 4160
rect 9640 4150 9680 4160
rect 9800 4150 9840 4160
rect 9880 4150 9920 4160
rect 9960 4150 9990 4160
rect 4120 4140 4200 4150
rect 4360 4140 4640 4150
rect 4720 4140 5000 4150
rect 5600 4140 5680 4150
rect 5920 4140 6440 4150
rect 6520 4140 6680 4150
rect 7440 4140 7480 4150
rect 8800 4140 8840 4150
rect 9640 4140 9680 4150
rect 9800 4140 9840 4150
rect 9880 4140 9920 4150
rect 9960 4140 9990 4150
rect 3240 4130 3280 4140
rect 4080 4130 4160 4140
rect 4400 4130 4560 4140
rect 5440 4130 5520 4140
rect 5640 4130 5720 4140
rect 5960 4130 6400 4140
rect 6480 4130 6680 4140
rect 9800 4130 9880 4140
rect 3240 4120 3280 4130
rect 4080 4120 4160 4130
rect 4400 4120 4560 4130
rect 5440 4120 5520 4130
rect 5640 4120 5720 4130
rect 5960 4120 6400 4130
rect 6480 4120 6680 4130
rect 9800 4120 9880 4130
rect 3240 4110 3280 4120
rect 4080 4110 4160 4120
rect 4400 4110 4560 4120
rect 5440 4110 5520 4120
rect 5640 4110 5720 4120
rect 5960 4110 6400 4120
rect 6480 4110 6680 4120
rect 9800 4110 9880 4120
rect 3240 4100 3280 4110
rect 4080 4100 4160 4110
rect 4400 4100 4560 4110
rect 5440 4100 5520 4110
rect 5640 4100 5720 4110
rect 5960 4100 6400 4110
rect 6480 4100 6680 4110
rect 9800 4100 9880 4110
rect 3160 4090 3280 4100
rect 4080 4090 4120 4100
rect 4440 4090 4560 4100
rect 4840 4090 4920 4100
rect 5040 4090 5080 4100
rect 5480 4090 5520 4100
rect 5680 4090 5840 4100
rect 5960 4090 6360 4100
rect 6440 4090 6640 4100
rect 7200 4090 7240 4100
rect 9600 4090 9760 4100
rect 9880 4090 9920 4100
rect 3160 4080 3280 4090
rect 4080 4080 4120 4090
rect 4440 4080 4560 4090
rect 4840 4080 4920 4090
rect 5040 4080 5080 4090
rect 5480 4080 5520 4090
rect 5680 4080 5840 4090
rect 5960 4080 6360 4090
rect 6440 4080 6640 4090
rect 7200 4080 7240 4090
rect 9600 4080 9760 4090
rect 9880 4080 9920 4090
rect 3160 4070 3280 4080
rect 4080 4070 4120 4080
rect 4440 4070 4560 4080
rect 4840 4070 4920 4080
rect 5040 4070 5080 4080
rect 5480 4070 5520 4080
rect 5680 4070 5840 4080
rect 5960 4070 6360 4080
rect 6440 4070 6640 4080
rect 7200 4070 7240 4080
rect 9600 4070 9760 4080
rect 9880 4070 9920 4080
rect 3160 4060 3280 4070
rect 4080 4060 4120 4070
rect 4440 4060 4560 4070
rect 4840 4060 4920 4070
rect 5040 4060 5080 4070
rect 5480 4060 5520 4070
rect 5680 4060 5840 4070
rect 5960 4060 6360 4070
rect 6440 4060 6640 4070
rect 7200 4060 7240 4070
rect 9600 4060 9760 4070
rect 9880 4060 9920 4070
rect 3080 4050 3280 4060
rect 4040 4050 4080 4060
rect 4160 4050 4280 4060
rect 4480 4050 4560 4060
rect 4760 4050 4800 4060
rect 4840 4050 4920 4060
rect 5040 4050 5080 4060
rect 5400 4050 5440 4060
rect 5480 4050 5520 4060
rect 5760 4050 6280 4060
rect 6400 4050 6640 4060
rect 8760 4050 8800 4060
rect 3080 4040 3280 4050
rect 4040 4040 4080 4050
rect 4160 4040 4280 4050
rect 4480 4040 4560 4050
rect 4760 4040 4800 4050
rect 4840 4040 4920 4050
rect 5040 4040 5080 4050
rect 5400 4040 5440 4050
rect 5480 4040 5520 4050
rect 5760 4040 6280 4050
rect 6400 4040 6640 4050
rect 8760 4040 8800 4050
rect 3080 4030 3280 4040
rect 4040 4030 4080 4040
rect 4160 4030 4280 4040
rect 4480 4030 4560 4040
rect 4760 4030 4800 4040
rect 4840 4030 4920 4040
rect 5040 4030 5080 4040
rect 5400 4030 5440 4040
rect 5480 4030 5520 4040
rect 5760 4030 6280 4040
rect 6400 4030 6640 4040
rect 8760 4030 8800 4040
rect 3080 4020 3280 4030
rect 4040 4020 4080 4030
rect 4160 4020 4280 4030
rect 4480 4020 4560 4030
rect 4760 4020 4800 4030
rect 4840 4020 4920 4030
rect 5040 4020 5080 4030
rect 5400 4020 5440 4030
rect 5480 4020 5520 4030
rect 5760 4020 6280 4030
rect 6400 4020 6640 4030
rect 8760 4020 8800 4030
rect 3120 4010 3280 4020
rect 4040 4010 4080 4020
rect 4160 4010 4320 4020
rect 4520 4010 4560 4020
rect 4720 4010 4880 4020
rect 5040 4010 5120 4020
rect 5400 4010 5440 4020
rect 6000 4010 6200 4020
rect 6400 4010 6600 4020
rect 7120 4010 7160 4020
rect 8360 4010 8400 4020
rect 8440 4010 8480 4020
rect 8560 4010 8640 4020
rect 3120 4000 3280 4010
rect 4040 4000 4080 4010
rect 4160 4000 4320 4010
rect 4520 4000 4560 4010
rect 4720 4000 4880 4010
rect 5040 4000 5120 4010
rect 5400 4000 5440 4010
rect 6000 4000 6200 4010
rect 6400 4000 6600 4010
rect 7120 4000 7160 4010
rect 8360 4000 8400 4010
rect 8440 4000 8480 4010
rect 8560 4000 8640 4010
rect 3120 3990 3280 4000
rect 4040 3990 4080 4000
rect 4160 3990 4320 4000
rect 4520 3990 4560 4000
rect 4720 3990 4880 4000
rect 5040 3990 5120 4000
rect 5400 3990 5440 4000
rect 6000 3990 6200 4000
rect 6400 3990 6600 4000
rect 7120 3990 7160 4000
rect 8360 3990 8400 4000
rect 8440 3990 8480 4000
rect 8560 3990 8640 4000
rect 3120 3980 3280 3990
rect 4040 3980 4080 3990
rect 4160 3980 4320 3990
rect 4520 3980 4560 3990
rect 4720 3980 4880 3990
rect 5040 3980 5120 3990
rect 5400 3980 5440 3990
rect 6000 3980 6200 3990
rect 6400 3980 6600 3990
rect 7120 3980 7160 3990
rect 8360 3980 8400 3990
rect 8440 3980 8480 3990
rect 8560 3980 8640 3990
rect 3200 3970 3240 3980
rect 4000 3970 4040 3980
rect 4120 3970 4160 3980
rect 4280 3970 4360 3980
rect 4520 3970 4720 3980
rect 4800 3970 4840 3980
rect 5440 3970 5480 3980
rect 6400 3970 6600 3980
rect 7120 3970 7160 3980
rect 8240 3970 8280 3980
rect 8320 3970 8360 3980
rect 8440 3970 8520 3980
rect 8560 3970 8600 3980
rect 8640 3970 8760 3980
rect 9680 3970 9720 3980
rect 3200 3960 3240 3970
rect 4000 3960 4040 3970
rect 4120 3960 4160 3970
rect 4280 3960 4360 3970
rect 4520 3960 4720 3970
rect 4800 3960 4840 3970
rect 5440 3960 5480 3970
rect 6400 3960 6600 3970
rect 7120 3960 7160 3970
rect 8240 3960 8280 3970
rect 8320 3960 8360 3970
rect 8440 3960 8520 3970
rect 8560 3960 8600 3970
rect 8640 3960 8760 3970
rect 9680 3960 9720 3970
rect 3200 3950 3240 3960
rect 4000 3950 4040 3960
rect 4120 3950 4160 3960
rect 4280 3950 4360 3960
rect 4520 3950 4720 3960
rect 4800 3950 4840 3960
rect 5440 3950 5480 3960
rect 6400 3950 6600 3960
rect 7120 3950 7160 3960
rect 8240 3950 8280 3960
rect 8320 3950 8360 3960
rect 8440 3950 8520 3960
rect 8560 3950 8600 3960
rect 8640 3950 8760 3960
rect 9680 3950 9720 3960
rect 3200 3940 3240 3950
rect 4000 3940 4040 3950
rect 4120 3940 4160 3950
rect 4280 3940 4360 3950
rect 4520 3940 4720 3950
rect 4800 3940 4840 3950
rect 5440 3940 5480 3950
rect 6400 3940 6600 3950
rect 7120 3940 7160 3950
rect 8240 3940 8280 3950
rect 8320 3940 8360 3950
rect 8440 3940 8520 3950
rect 8560 3940 8600 3950
rect 8640 3940 8760 3950
rect 9680 3940 9720 3950
rect 3200 3930 3280 3940
rect 4080 3930 4120 3940
rect 4320 3930 4360 3940
rect 4520 3930 4720 3940
rect 5120 3930 5160 3940
rect 6400 3930 6600 3940
rect 7120 3930 7160 3940
rect 8000 3930 8040 3940
rect 8240 3930 8280 3940
rect 8440 3930 8520 3940
rect 8680 3930 8720 3940
rect 9600 3930 9640 3940
rect 9720 3930 9760 3940
rect 3200 3920 3280 3930
rect 4080 3920 4120 3930
rect 4320 3920 4360 3930
rect 4520 3920 4720 3930
rect 5120 3920 5160 3930
rect 6400 3920 6600 3930
rect 7120 3920 7160 3930
rect 8000 3920 8040 3930
rect 8240 3920 8280 3930
rect 8440 3920 8520 3930
rect 8680 3920 8720 3930
rect 9600 3920 9640 3930
rect 9720 3920 9760 3930
rect 3200 3910 3280 3920
rect 4080 3910 4120 3920
rect 4320 3910 4360 3920
rect 4520 3910 4720 3920
rect 5120 3910 5160 3920
rect 6400 3910 6600 3920
rect 7120 3910 7160 3920
rect 8000 3910 8040 3920
rect 8240 3910 8280 3920
rect 8440 3910 8520 3920
rect 8680 3910 8720 3920
rect 9600 3910 9640 3920
rect 9720 3910 9760 3920
rect 3200 3900 3280 3910
rect 4080 3900 4120 3910
rect 4320 3900 4360 3910
rect 4520 3900 4720 3910
rect 5120 3900 5160 3910
rect 6400 3900 6600 3910
rect 7120 3900 7160 3910
rect 8000 3900 8040 3910
rect 8240 3900 8280 3910
rect 8440 3900 8520 3910
rect 8680 3900 8720 3910
rect 9600 3900 9640 3910
rect 9720 3900 9760 3910
rect 3160 3890 3200 3900
rect 3920 3890 3960 3900
rect 4000 3890 4080 3900
rect 4320 3890 4400 3900
rect 4560 3890 4640 3900
rect 5160 3890 5200 3900
rect 6440 3890 6600 3900
rect 8000 3890 8040 3900
rect 8200 3890 8240 3900
rect 8320 3890 8360 3900
rect 8400 3890 8480 3900
rect 8600 3890 8720 3900
rect 9440 3890 9480 3900
rect 9720 3890 9840 3900
rect 3160 3880 3200 3890
rect 3920 3880 3960 3890
rect 4000 3880 4080 3890
rect 4320 3880 4400 3890
rect 4560 3880 4640 3890
rect 5160 3880 5200 3890
rect 6440 3880 6600 3890
rect 8000 3880 8040 3890
rect 8200 3880 8240 3890
rect 8320 3880 8360 3890
rect 8400 3880 8480 3890
rect 8600 3880 8720 3890
rect 9440 3880 9480 3890
rect 9720 3880 9840 3890
rect 3160 3870 3200 3880
rect 3920 3870 3960 3880
rect 4000 3870 4080 3880
rect 4320 3870 4400 3880
rect 4560 3870 4640 3880
rect 5160 3870 5200 3880
rect 6440 3870 6600 3880
rect 8000 3870 8040 3880
rect 8200 3870 8240 3880
rect 8320 3870 8360 3880
rect 8400 3870 8480 3880
rect 8600 3870 8720 3880
rect 9440 3870 9480 3880
rect 9720 3870 9840 3880
rect 3160 3860 3200 3870
rect 3920 3860 3960 3870
rect 4000 3860 4080 3870
rect 4320 3860 4400 3870
rect 4560 3860 4640 3870
rect 5160 3860 5200 3870
rect 6440 3860 6600 3870
rect 8000 3860 8040 3870
rect 8200 3860 8240 3870
rect 8320 3860 8360 3870
rect 8400 3860 8480 3870
rect 8600 3860 8720 3870
rect 9440 3860 9480 3870
rect 9720 3860 9840 3870
rect 3160 3850 3200 3860
rect 3240 3850 3280 3860
rect 3880 3850 3920 3860
rect 3960 3850 4080 3860
rect 4320 3850 4400 3860
rect 4600 3850 4640 3860
rect 5160 3850 5200 3860
rect 6520 3850 6600 3860
rect 7080 3850 7120 3860
rect 8240 3850 8280 3860
rect 8320 3850 8480 3860
rect 8560 3850 8680 3860
rect 9560 3850 9600 3860
rect 9720 3850 9880 3860
rect 3160 3840 3200 3850
rect 3240 3840 3280 3850
rect 3880 3840 3920 3850
rect 3960 3840 4080 3850
rect 4320 3840 4400 3850
rect 4600 3840 4640 3850
rect 5160 3840 5200 3850
rect 6520 3840 6600 3850
rect 7080 3840 7120 3850
rect 8240 3840 8280 3850
rect 8320 3840 8480 3850
rect 8560 3840 8680 3850
rect 9560 3840 9600 3850
rect 9720 3840 9880 3850
rect 3160 3830 3200 3840
rect 3240 3830 3280 3840
rect 3880 3830 3920 3840
rect 3960 3830 4080 3840
rect 4320 3830 4400 3840
rect 4600 3830 4640 3840
rect 5160 3830 5200 3840
rect 6520 3830 6600 3840
rect 7080 3830 7120 3840
rect 8240 3830 8280 3840
rect 8320 3830 8480 3840
rect 8560 3830 8680 3840
rect 9560 3830 9600 3840
rect 9720 3830 9880 3840
rect 3160 3820 3200 3830
rect 3240 3820 3280 3830
rect 3880 3820 3920 3830
rect 3960 3820 4080 3830
rect 4320 3820 4400 3830
rect 4600 3820 4640 3830
rect 5160 3820 5200 3830
rect 6520 3820 6600 3830
rect 7080 3820 7120 3830
rect 8240 3820 8280 3830
rect 8320 3820 8480 3830
rect 8560 3820 8680 3830
rect 9560 3820 9600 3830
rect 9720 3820 9880 3830
rect 3000 3810 3080 3820
rect 3240 3810 3280 3820
rect 3880 3810 4040 3820
rect 4280 3810 4440 3820
rect 5160 3810 5240 3820
rect 6520 3810 6600 3820
rect 8280 3810 8520 3820
rect 8640 3810 8680 3820
rect 9840 3810 9880 3820
rect 3000 3800 3080 3810
rect 3240 3800 3280 3810
rect 3880 3800 4040 3810
rect 4280 3800 4440 3810
rect 5160 3800 5240 3810
rect 6520 3800 6600 3810
rect 8280 3800 8520 3810
rect 8640 3800 8680 3810
rect 9840 3800 9880 3810
rect 3000 3790 3080 3800
rect 3240 3790 3280 3800
rect 3880 3790 4040 3800
rect 4280 3790 4440 3800
rect 5160 3790 5240 3800
rect 6520 3790 6600 3800
rect 8280 3790 8520 3800
rect 8640 3790 8680 3800
rect 9840 3790 9880 3800
rect 3000 3780 3080 3790
rect 3240 3780 3280 3790
rect 3880 3780 4040 3790
rect 4280 3780 4440 3790
rect 5160 3780 5240 3790
rect 6520 3780 6600 3790
rect 8280 3780 8520 3790
rect 8640 3780 8680 3790
rect 9840 3780 9880 3790
rect 2960 3770 3080 3780
rect 3200 3770 3280 3780
rect 3920 3770 4000 3780
rect 4160 3770 4440 3780
rect 4840 3770 4920 3780
rect 5160 3770 5240 3780
rect 6520 3770 6600 3780
rect 8360 3770 8400 3780
rect 8480 3770 8560 3780
rect 9640 3770 9680 3780
rect 9840 3770 9880 3780
rect 2960 3760 3080 3770
rect 3200 3760 3280 3770
rect 3920 3760 4000 3770
rect 4160 3760 4440 3770
rect 4840 3760 4920 3770
rect 5160 3760 5240 3770
rect 6520 3760 6600 3770
rect 8360 3760 8400 3770
rect 8480 3760 8560 3770
rect 9640 3760 9680 3770
rect 9840 3760 9880 3770
rect 2960 3750 3080 3760
rect 3200 3750 3280 3760
rect 3920 3750 4000 3760
rect 4160 3750 4440 3760
rect 4840 3750 4920 3760
rect 5160 3750 5240 3760
rect 6520 3750 6600 3760
rect 8360 3750 8400 3760
rect 8480 3750 8560 3760
rect 9640 3750 9680 3760
rect 9840 3750 9880 3760
rect 2960 3740 3080 3750
rect 3200 3740 3280 3750
rect 3920 3740 4000 3750
rect 4160 3740 4440 3750
rect 4840 3740 4920 3750
rect 5160 3740 5240 3750
rect 6520 3740 6600 3750
rect 8360 3740 8400 3750
rect 8480 3740 8560 3750
rect 9640 3740 9680 3750
rect 9840 3740 9880 3750
rect 3000 3730 3120 3740
rect 3160 3730 3280 3740
rect 3920 3730 3960 3740
rect 4040 3730 4080 3740
rect 4120 3730 4200 3740
rect 4240 3730 4440 3740
rect 4800 3730 4840 3740
rect 4880 3730 5280 3740
rect 6520 3730 6600 3740
rect 7000 3730 7040 3740
rect 8520 3730 8560 3740
rect 9680 3730 9990 3740
rect 3000 3720 3120 3730
rect 3160 3720 3280 3730
rect 3920 3720 3960 3730
rect 4040 3720 4080 3730
rect 4120 3720 4200 3730
rect 4240 3720 4440 3730
rect 4800 3720 4840 3730
rect 4880 3720 5280 3730
rect 6520 3720 6600 3730
rect 7000 3720 7040 3730
rect 8520 3720 8560 3730
rect 9680 3720 9990 3730
rect 3000 3710 3120 3720
rect 3160 3710 3280 3720
rect 3920 3710 3960 3720
rect 4040 3710 4080 3720
rect 4120 3710 4200 3720
rect 4240 3710 4440 3720
rect 4800 3710 4840 3720
rect 4880 3710 5280 3720
rect 6520 3710 6600 3720
rect 7000 3710 7040 3720
rect 8520 3710 8560 3720
rect 9680 3710 9990 3720
rect 3000 3700 3120 3710
rect 3160 3700 3280 3710
rect 3920 3700 3960 3710
rect 4040 3700 4080 3710
rect 4120 3700 4200 3710
rect 4240 3700 4440 3710
rect 4800 3700 4840 3710
rect 4880 3700 5280 3710
rect 6520 3700 6600 3710
rect 7000 3700 7040 3710
rect 8520 3700 8560 3710
rect 9680 3700 9990 3710
rect 3080 3690 3280 3700
rect 4000 3690 4120 3700
rect 4160 3690 4240 3700
rect 4320 3690 4440 3700
rect 4800 3690 4880 3700
rect 5000 3690 5280 3700
rect 6560 3690 6600 3700
rect 6960 3690 7000 3700
rect 8200 3690 8240 3700
rect 8360 3690 8400 3700
rect 8480 3690 8520 3700
rect 8600 3690 8640 3700
rect 9560 3690 9640 3700
rect 9840 3690 9960 3700
rect 3080 3680 3280 3690
rect 4000 3680 4120 3690
rect 4160 3680 4240 3690
rect 4320 3680 4440 3690
rect 4800 3680 4880 3690
rect 5000 3680 5280 3690
rect 6560 3680 6600 3690
rect 6960 3680 7000 3690
rect 8200 3680 8240 3690
rect 8360 3680 8400 3690
rect 8480 3680 8520 3690
rect 8600 3680 8640 3690
rect 9560 3680 9640 3690
rect 9840 3680 9960 3690
rect 3080 3670 3280 3680
rect 4000 3670 4120 3680
rect 4160 3670 4240 3680
rect 4320 3670 4440 3680
rect 4800 3670 4880 3680
rect 5000 3670 5280 3680
rect 6560 3670 6600 3680
rect 6960 3670 7000 3680
rect 8200 3670 8240 3680
rect 8360 3670 8400 3680
rect 8480 3670 8520 3680
rect 8600 3670 8640 3680
rect 9560 3670 9640 3680
rect 9840 3670 9960 3680
rect 3080 3660 3280 3670
rect 4000 3660 4120 3670
rect 4160 3660 4240 3670
rect 4320 3660 4440 3670
rect 4800 3660 4880 3670
rect 5000 3660 5280 3670
rect 6560 3660 6600 3670
rect 6960 3660 7000 3670
rect 8200 3660 8240 3670
rect 8360 3660 8400 3670
rect 8480 3660 8520 3670
rect 8600 3660 8640 3670
rect 9560 3660 9640 3670
rect 9840 3660 9960 3670
rect 3240 3650 3280 3660
rect 3960 3650 4040 3660
rect 4320 3650 4440 3660
rect 4800 3650 4960 3660
rect 5120 3650 5280 3660
rect 6520 3650 6600 3660
rect 9520 3650 9560 3660
rect 9640 3650 9680 3660
rect 9840 3650 9920 3660
rect 3240 3640 3280 3650
rect 3960 3640 4040 3650
rect 4320 3640 4440 3650
rect 4800 3640 4960 3650
rect 5120 3640 5280 3650
rect 6520 3640 6600 3650
rect 9520 3640 9560 3650
rect 9640 3640 9680 3650
rect 9840 3640 9920 3650
rect 3240 3630 3280 3640
rect 3960 3630 4040 3640
rect 4320 3630 4440 3640
rect 4800 3630 4960 3640
rect 5120 3630 5280 3640
rect 6520 3630 6600 3640
rect 9520 3630 9560 3640
rect 9640 3630 9680 3640
rect 9840 3630 9920 3640
rect 3240 3620 3280 3630
rect 3960 3620 4040 3630
rect 4320 3620 4440 3630
rect 4800 3620 4960 3630
rect 5120 3620 5280 3630
rect 6520 3620 6600 3630
rect 9520 3620 9560 3630
rect 9640 3620 9680 3630
rect 9840 3620 9920 3630
rect 3920 3610 4040 3620
rect 4320 3610 4440 3620
rect 4760 3610 4840 3620
rect 4880 3610 5040 3620
rect 5120 3610 5320 3620
rect 6520 3610 6600 3620
rect 9440 3610 9480 3620
rect 9560 3610 9680 3620
rect 3920 3600 4040 3610
rect 4320 3600 4440 3610
rect 4760 3600 4840 3610
rect 4880 3600 5040 3610
rect 5120 3600 5320 3610
rect 6520 3600 6600 3610
rect 9440 3600 9480 3610
rect 9560 3600 9680 3610
rect 3920 3590 4040 3600
rect 4320 3590 4440 3600
rect 4760 3590 4840 3600
rect 4880 3590 5040 3600
rect 5120 3590 5320 3600
rect 6520 3590 6600 3600
rect 9440 3590 9480 3600
rect 9560 3590 9680 3600
rect 3920 3580 4040 3590
rect 4320 3580 4440 3590
rect 4760 3580 4840 3590
rect 4880 3580 5040 3590
rect 5120 3580 5320 3590
rect 6520 3580 6600 3590
rect 9440 3580 9480 3590
rect 9560 3580 9680 3590
rect 3280 3570 3360 3580
rect 3960 3570 4040 3580
rect 4280 3570 4480 3580
rect 4680 3570 4720 3580
rect 4800 3570 4840 3580
rect 5000 3570 5080 3580
rect 5120 3570 5320 3580
rect 6520 3570 6600 3580
rect 6880 3570 6920 3580
rect 8360 3570 8400 3580
rect 8480 3570 8520 3580
rect 9240 3570 9400 3580
rect 9640 3570 9680 3580
rect 3280 3560 3360 3570
rect 3960 3560 4040 3570
rect 4280 3560 4480 3570
rect 4680 3560 4720 3570
rect 4800 3560 4840 3570
rect 5000 3560 5080 3570
rect 5120 3560 5320 3570
rect 6520 3560 6600 3570
rect 6880 3560 6920 3570
rect 8360 3560 8400 3570
rect 8480 3560 8520 3570
rect 9240 3560 9400 3570
rect 9640 3560 9680 3570
rect 3280 3550 3360 3560
rect 3960 3550 4040 3560
rect 4280 3550 4480 3560
rect 4680 3550 4720 3560
rect 4800 3550 4840 3560
rect 5000 3550 5080 3560
rect 5120 3550 5320 3560
rect 6520 3550 6600 3560
rect 6880 3550 6920 3560
rect 8360 3550 8400 3560
rect 8480 3550 8520 3560
rect 9240 3550 9400 3560
rect 9640 3550 9680 3560
rect 3280 3540 3360 3550
rect 3960 3540 4040 3550
rect 4280 3540 4480 3550
rect 4680 3540 4720 3550
rect 4800 3540 4840 3550
rect 5000 3540 5080 3550
rect 5120 3540 5320 3550
rect 6520 3540 6600 3550
rect 6880 3540 6920 3550
rect 8360 3540 8400 3550
rect 8480 3540 8520 3550
rect 9240 3540 9400 3550
rect 9640 3540 9680 3550
rect 3320 3530 3400 3540
rect 4000 3530 4040 3540
rect 4240 3530 4520 3540
rect 4600 3530 4680 3540
rect 4760 3530 4840 3540
rect 5080 3530 5320 3540
rect 6480 3530 6560 3540
rect 6840 3530 6880 3540
rect 8360 3530 8400 3540
rect 8480 3530 8520 3540
rect 9160 3530 9240 3540
rect 9440 3530 9480 3540
rect 9600 3530 9680 3540
rect 3320 3520 3400 3530
rect 4000 3520 4040 3530
rect 4240 3520 4520 3530
rect 4600 3520 4680 3530
rect 4760 3520 4840 3530
rect 5080 3520 5320 3530
rect 6480 3520 6560 3530
rect 6840 3520 6880 3530
rect 8360 3520 8400 3530
rect 8480 3520 8520 3530
rect 9160 3520 9240 3530
rect 9440 3520 9480 3530
rect 9600 3520 9680 3530
rect 3320 3510 3400 3520
rect 4000 3510 4040 3520
rect 4240 3510 4520 3520
rect 4600 3510 4680 3520
rect 4760 3510 4840 3520
rect 5080 3510 5320 3520
rect 6480 3510 6560 3520
rect 6840 3510 6880 3520
rect 8360 3510 8400 3520
rect 8480 3510 8520 3520
rect 9160 3510 9240 3520
rect 9440 3510 9480 3520
rect 9600 3510 9680 3520
rect 3320 3500 3400 3510
rect 4000 3500 4040 3510
rect 4240 3500 4520 3510
rect 4600 3500 4680 3510
rect 4760 3500 4840 3510
rect 5080 3500 5320 3510
rect 6480 3500 6560 3510
rect 6840 3500 6880 3510
rect 8360 3500 8400 3510
rect 8480 3500 8520 3510
rect 9160 3500 9240 3510
rect 9440 3500 9480 3510
rect 9600 3500 9680 3510
rect 2400 3490 2480 3500
rect 2600 3490 2680 3500
rect 3360 3490 3400 3500
rect 4000 3490 4080 3500
rect 4200 3490 4280 3500
rect 4400 3490 4480 3500
rect 4760 3490 4800 3500
rect 4920 3490 4960 3500
rect 5040 3490 5320 3500
rect 6480 3490 6560 3500
rect 6800 3490 6840 3500
rect 8520 3490 8560 3500
rect 9120 3490 9200 3500
rect 9360 3490 9400 3500
rect 9520 3490 9560 3500
rect 9600 3490 9640 3500
rect 2400 3480 2480 3490
rect 2600 3480 2680 3490
rect 3360 3480 3400 3490
rect 4000 3480 4080 3490
rect 4200 3480 4280 3490
rect 4400 3480 4480 3490
rect 4760 3480 4800 3490
rect 4920 3480 4960 3490
rect 5040 3480 5320 3490
rect 6480 3480 6560 3490
rect 6800 3480 6840 3490
rect 8520 3480 8560 3490
rect 9120 3480 9200 3490
rect 9360 3480 9400 3490
rect 9520 3480 9560 3490
rect 9600 3480 9640 3490
rect 2400 3470 2480 3480
rect 2600 3470 2680 3480
rect 3360 3470 3400 3480
rect 4000 3470 4080 3480
rect 4200 3470 4280 3480
rect 4400 3470 4480 3480
rect 4760 3470 4800 3480
rect 4920 3470 4960 3480
rect 5040 3470 5320 3480
rect 6480 3470 6560 3480
rect 6800 3470 6840 3480
rect 8520 3470 8560 3480
rect 9120 3470 9200 3480
rect 9360 3470 9400 3480
rect 9520 3470 9560 3480
rect 9600 3470 9640 3480
rect 2400 3460 2480 3470
rect 2600 3460 2680 3470
rect 3360 3460 3400 3470
rect 4000 3460 4080 3470
rect 4200 3460 4280 3470
rect 4400 3460 4480 3470
rect 4760 3460 4800 3470
rect 4920 3460 4960 3470
rect 5040 3460 5320 3470
rect 6480 3460 6560 3470
rect 6800 3460 6840 3470
rect 8520 3460 8560 3470
rect 9120 3460 9200 3470
rect 9360 3460 9400 3470
rect 9520 3460 9560 3470
rect 9600 3460 9640 3470
rect 2280 3450 2360 3460
rect 2840 3450 2880 3460
rect 4000 3450 4080 3460
rect 4160 3450 4280 3460
rect 4760 3450 4800 3460
rect 4840 3450 4880 3460
rect 5120 3450 5320 3460
rect 6440 3450 6560 3460
rect 9080 3450 9160 3460
rect 9240 3450 9280 3460
rect 9440 3450 9520 3460
rect 2280 3440 2360 3450
rect 2840 3440 2880 3450
rect 4000 3440 4080 3450
rect 4160 3440 4280 3450
rect 4760 3440 4800 3450
rect 4840 3440 4880 3450
rect 5120 3440 5320 3450
rect 6440 3440 6560 3450
rect 9080 3440 9160 3450
rect 9240 3440 9280 3450
rect 9440 3440 9520 3450
rect 2280 3430 2360 3440
rect 2840 3430 2880 3440
rect 4000 3430 4080 3440
rect 4160 3430 4280 3440
rect 4760 3430 4800 3440
rect 4840 3430 4880 3440
rect 5120 3430 5320 3440
rect 6440 3430 6560 3440
rect 9080 3430 9160 3440
rect 9240 3430 9280 3440
rect 9440 3430 9520 3440
rect 2280 3420 2360 3430
rect 2840 3420 2880 3430
rect 4000 3420 4080 3430
rect 4160 3420 4280 3430
rect 4760 3420 4800 3430
rect 4840 3420 4880 3430
rect 5120 3420 5320 3430
rect 6440 3420 6560 3430
rect 9080 3420 9160 3430
rect 9240 3420 9280 3430
rect 9440 3420 9520 3430
rect 2920 3410 2960 3420
rect 4000 3410 4240 3420
rect 4360 3410 4400 3420
rect 5000 3410 5040 3420
rect 5200 3410 5320 3420
rect 6400 3410 6520 3420
rect 6720 3410 6760 3420
rect 8520 3410 8560 3420
rect 9040 3410 9080 3420
rect 9400 3410 9440 3420
rect 9640 3410 9680 3420
rect 2920 3400 2960 3410
rect 4000 3400 4240 3410
rect 4360 3400 4400 3410
rect 5000 3400 5040 3410
rect 5200 3400 5320 3410
rect 6400 3400 6520 3410
rect 6720 3400 6760 3410
rect 8520 3400 8560 3410
rect 9040 3400 9080 3410
rect 9400 3400 9440 3410
rect 9640 3400 9680 3410
rect 2920 3390 2960 3400
rect 4000 3390 4240 3400
rect 4360 3390 4400 3400
rect 5000 3390 5040 3400
rect 5200 3390 5320 3400
rect 6400 3390 6520 3400
rect 6720 3390 6760 3400
rect 8520 3390 8560 3400
rect 9040 3390 9080 3400
rect 9400 3390 9440 3400
rect 9640 3390 9680 3400
rect 2920 3380 2960 3390
rect 4000 3380 4240 3390
rect 4360 3380 4400 3390
rect 5000 3380 5040 3390
rect 5200 3380 5320 3390
rect 6400 3380 6520 3390
rect 6720 3380 6760 3390
rect 8520 3380 8560 3390
rect 9040 3380 9080 3390
rect 9400 3380 9440 3390
rect 9640 3380 9680 3390
rect 3520 3370 3560 3380
rect 4040 3370 4240 3380
rect 4360 3370 4600 3380
rect 4880 3370 5040 3380
rect 5200 3370 5280 3380
rect 6360 3370 6520 3380
rect 6680 3370 6720 3380
rect 9040 3370 9080 3380
rect 9400 3370 9440 3380
rect 9640 3370 9720 3380
rect 9760 3370 9800 3380
rect 3520 3360 3560 3370
rect 4040 3360 4240 3370
rect 4360 3360 4600 3370
rect 4880 3360 5040 3370
rect 5200 3360 5280 3370
rect 6360 3360 6520 3370
rect 6680 3360 6720 3370
rect 9040 3360 9080 3370
rect 9400 3360 9440 3370
rect 9640 3360 9720 3370
rect 9760 3360 9800 3370
rect 3520 3350 3560 3360
rect 4040 3350 4240 3360
rect 4360 3350 4600 3360
rect 4880 3350 5040 3360
rect 5200 3350 5280 3360
rect 6360 3350 6520 3360
rect 6680 3350 6720 3360
rect 9040 3350 9080 3360
rect 9400 3350 9440 3360
rect 9640 3350 9720 3360
rect 9760 3350 9800 3360
rect 3520 3340 3560 3350
rect 4040 3340 4240 3350
rect 4360 3340 4600 3350
rect 4880 3340 5040 3350
rect 5200 3340 5280 3350
rect 6360 3340 6520 3350
rect 6680 3340 6720 3350
rect 9040 3340 9080 3350
rect 9400 3340 9440 3350
rect 9640 3340 9720 3350
rect 9760 3340 9800 3350
rect 2160 3330 2200 3340
rect 3520 3330 3600 3340
rect 4360 3330 4400 3340
rect 4480 3330 4560 3340
rect 4840 3330 5040 3340
rect 5200 3330 5280 3340
rect 6320 3330 6520 3340
rect 6640 3330 6680 3340
rect 8480 3330 8520 3340
rect 8920 3330 9040 3340
rect 9320 3330 9400 3340
rect 9640 3330 9680 3340
rect 9760 3330 9800 3340
rect 2160 3320 2200 3330
rect 3520 3320 3600 3330
rect 4360 3320 4400 3330
rect 4480 3320 4560 3330
rect 4840 3320 5040 3330
rect 5200 3320 5280 3330
rect 6320 3320 6520 3330
rect 6640 3320 6680 3330
rect 8480 3320 8520 3330
rect 8920 3320 9040 3330
rect 9320 3320 9400 3330
rect 9640 3320 9680 3330
rect 9760 3320 9800 3330
rect 2160 3310 2200 3320
rect 3520 3310 3600 3320
rect 4360 3310 4400 3320
rect 4480 3310 4560 3320
rect 4840 3310 5040 3320
rect 5200 3310 5280 3320
rect 6320 3310 6520 3320
rect 6640 3310 6680 3320
rect 8480 3310 8520 3320
rect 8920 3310 9040 3320
rect 9320 3310 9400 3320
rect 9640 3310 9680 3320
rect 9760 3310 9800 3320
rect 2160 3300 2200 3310
rect 3520 3300 3600 3310
rect 4360 3300 4400 3310
rect 4480 3300 4560 3310
rect 4840 3300 5040 3310
rect 5200 3300 5280 3310
rect 6320 3300 6520 3310
rect 6640 3300 6680 3310
rect 8480 3300 8520 3310
rect 8920 3300 9040 3310
rect 9320 3300 9400 3310
rect 9640 3300 9680 3310
rect 9760 3300 9800 3310
rect 2120 3290 2160 3300
rect 4360 3290 4480 3300
rect 4760 3290 4960 3300
rect 5200 3290 5280 3300
rect 6240 3290 6520 3300
rect 6560 3290 6640 3300
rect 8840 3290 9040 3300
rect 9320 3290 9360 3300
rect 9440 3290 9480 3300
rect 9560 3290 9600 3300
rect 9720 3290 9760 3300
rect 9960 3290 9990 3300
rect 2120 3280 2160 3290
rect 4360 3280 4480 3290
rect 4760 3280 4960 3290
rect 5200 3280 5280 3290
rect 6240 3280 6520 3290
rect 6560 3280 6640 3290
rect 8840 3280 9040 3290
rect 9320 3280 9360 3290
rect 9440 3280 9480 3290
rect 9560 3280 9600 3290
rect 9720 3280 9760 3290
rect 9960 3280 9990 3290
rect 2120 3270 2160 3280
rect 4360 3270 4480 3280
rect 4760 3270 4960 3280
rect 5200 3270 5280 3280
rect 6240 3270 6520 3280
rect 6560 3270 6640 3280
rect 8840 3270 9040 3280
rect 9320 3270 9360 3280
rect 9440 3270 9480 3280
rect 9560 3270 9600 3280
rect 9720 3270 9760 3280
rect 9960 3270 9990 3280
rect 2120 3260 2160 3270
rect 4360 3260 4480 3270
rect 4760 3260 4960 3270
rect 5200 3260 5280 3270
rect 6240 3260 6520 3270
rect 6560 3260 6640 3270
rect 8840 3260 9040 3270
rect 9320 3260 9360 3270
rect 9440 3260 9480 3270
rect 9560 3260 9600 3270
rect 9720 3260 9760 3270
rect 9960 3260 9990 3270
rect 3120 3250 3160 3260
rect 4680 3250 4920 3260
rect 5200 3250 5280 3260
rect 6240 3250 6480 3260
rect 8440 3250 8480 3260
rect 8960 3250 9040 3260
rect 9120 3250 9160 3260
rect 9280 3250 9360 3260
rect 9440 3250 9520 3260
rect 9680 3250 9720 3260
rect 9920 3250 9990 3260
rect 3120 3240 3160 3250
rect 4680 3240 4920 3250
rect 5200 3240 5280 3250
rect 6240 3240 6480 3250
rect 8440 3240 8480 3250
rect 8960 3240 9040 3250
rect 9120 3240 9160 3250
rect 9280 3240 9360 3250
rect 9440 3240 9520 3250
rect 9680 3240 9720 3250
rect 9920 3240 9990 3250
rect 3120 3230 3160 3240
rect 4680 3230 4920 3240
rect 5200 3230 5280 3240
rect 6240 3230 6480 3240
rect 8440 3230 8480 3240
rect 8960 3230 9040 3240
rect 9120 3230 9160 3240
rect 9280 3230 9360 3240
rect 9440 3230 9520 3240
rect 9680 3230 9720 3240
rect 9920 3230 9990 3240
rect 3120 3220 3160 3230
rect 4680 3220 4920 3230
rect 5200 3220 5280 3230
rect 6240 3220 6480 3230
rect 8440 3220 8480 3230
rect 8960 3220 9040 3230
rect 9120 3220 9160 3230
rect 9280 3220 9360 3230
rect 9440 3220 9520 3230
rect 9680 3220 9720 3230
rect 9920 3220 9990 3230
rect 2080 3210 2120 3220
rect 4600 3210 4880 3220
rect 4960 3210 5000 3220
rect 5200 3210 5280 3220
rect 6280 3210 6400 3220
rect 9000 3210 9040 3220
rect 9280 3210 9320 3220
rect 9400 3210 9480 3220
rect 9600 3210 9640 3220
rect 9880 3210 9990 3220
rect 2080 3200 2120 3210
rect 4600 3200 4880 3210
rect 4960 3200 5000 3210
rect 5200 3200 5280 3210
rect 6280 3200 6400 3210
rect 9000 3200 9040 3210
rect 9280 3200 9320 3210
rect 9400 3200 9480 3210
rect 9600 3200 9640 3210
rect 9880 3200 9990 3210
rect 2080 3190 2120 3200
rect 4600 3190 4880 3200
rect 4960 3190 5000 3200
rect 5200 3190 5280 3200
rect 6280 3190 6400 3200
rect 9000 3190 9040 3200
rect 9280 3190 9320 3200
rect 9400 3190 9480 3200
rect 9600 3190 9640 3200
rect 9880 3190 9990 3200
rect 2080 3180 2120 3190
rect 4600 3180 4880 3190
rect 4960 3180 5000 3190
rect 5200 3180 5280 3190
rect 6280 3180 6400 3190
rect 9000 3180 9040 3190
rect 9280 3180 9320 3190
rect 9400 3180 9480 3190
rect 9600 3180 9640 3190
rect 9880 3180 9990 3190
rect 2080 3170 2120 3180
rect 4240 3170 4320 3180
rect 4600 3170 4880 3180
rect 4960 3170 5000 3180
rect 5200 3170 5240 3180
rect 8400 3170 8440 3180
rect 8880 3170 9000 3180
rect 9400 3170 9440 3180
rect 9560 3170 9640 3180
rect 9880 3170 9920 3180
rect 9960 3170 9990 3180
rect 2080 3160 2120 3170
rect 4240 3160 4320 3170
rect 4600 3160 4880 3170
rect 4960 3160 5000 3170
rect 5200 3160 5240 3170
rect 8400 3160 8440 3170
rect 8880 3160 9000 3170
rect 9400 3160 9440 3170
rect 9560 3160 9640 3170
rect 9880 3160 9920 3170
rect 9960 3160 9990 3170
rect 2080 3150 2120 3160
rect 4240 3150 4320 3160
rect 4600 3150 4880 3160
rect 4960 3150 5000 3160
rect 5200 3150 5240 3160
rect 8400 3150 8440 3160
rect 8880 3150 9000 3160
rect 9400 3150 9440 3160
rect 9560 3150 9640 3160
rect 9880 3150 9920 3160
rect 9960 3150 9990 3160
rect 2080 3140 2120 3150
rect 4240 3140 4320 3150
rect 4600 3140 4880 3150
rect 4960 3140 5000 3150
rect 5200 3140 5240 3150
rect 8400 3140 8440 3150
rect 8880 3140 9000 3150
rect 9400 3140 9440 3150
rect 9560 3140 9640 3150
rect 9880 3140 9920 3150
rect 9960 3140 9990 3150
rect 2080 3130 2120 3140
rect 4240 3130 4480 3140
rect 4600 3130 4800 3140
rect 4920 3130 5000 3140
rect 5200 3130 5240 3140
rect 8800 3130 8920 3140
rect 8960 3130 9040 3140
rect 9840 3130 9920 3140
rect 2080 3120 2120 3130
rect 4240 3120 4480 3130
rect 4600 3120 4800 3130
rect 4920 3120 5000 3130
rect 5200 3120 5240 3130
rect 8800 3120 8920 3130
rect 8960 3120 9040 3130
rect 9840 3120 9920 3130
rect 2080 3110 2120 3120
rect 4240 3110 4480 3120
rect 4600 3110 4800 3120
rect 4920 3110 5000 3120
rect 5200 3110 5240 3120
rect 8800 3110 8920 3120
rect 8960 3110 9040 3120
rect 9840 3110 9920 3120
rect 2080 3100 2120 3110
rect 4240 3100 4480 3110
rect 4600 3100 4800 3110
rect 4920 3100 5000 3110
rect 5200 3100 5240 3110
rect 8800 3100 8920 3110
rect 8960 3100 9040 3110
rect 9840 3100 9920 3110
rect 2080 3090 2120 3100
rect 3880 3090 3920 3100
rect 3960 3090 4000 3100
rect 4280 3090 4520 3100
rect 4920 3090 5000 3100
rect 5160 3090 5240 3100
rect 8360 3090 8400 3100
rect 8840 3090 9000 3100
rect 9880 3090 9990 3100
rect 2080 3080 2120 3090
rect 3880 3080 3920 3090
rect 3960 3080 4000 3090
rect 4280 3080 4520 3090
rect 4920 3080 5000 3090
rect 5160 3080 5240 3090
rect 8360 3080 8400 3090
rect 8840 3080 9000 3090
rect 9880 3080 9990 3090
rect 2080 3070 2120 3080
rect 3880 3070 3920 3080
rect 3960 3070 4000 3080
rect 4280 3070 4520 3080
rect 4920 3070 5000 3080
rect 5160 3070 5240 3080
rect 8360 3070 8400 3080
rect 8840 3070 9000 3080
rect 9880 3070 9990 3080
rect 2080 3060 2120 3070
rect 3880 3060 3920 3070
rect 3960 3060 4000 3070
rect 4280 3060 4520 3070
rect 4920 3060 5000 3070
rect 5160 3060 5240 3070
rect 8360 3060 8400 3070
rect 8840 3060 9000 3070
rect 9880 3060 9990 3070
rect 2040 3050 2120 3060
rect 3120 3050 3160 3060
rect 3880 3050 3920 3060
rect 4320 3050 4360 3060
rect 4400 3050 4520 3060
rect 4880 3050 5000 3060
rect 5120 3050 5200 3060
rect 8400 3050 8440 3060
rect 8720 3050 8920 3060
rect 9480 3050 9520 3060
rect 9760 3050 9800 3060
rect 9880 3050 9960 3060
rect 2040 3040 2120 3050
rect 3120 3040 3160 3050
rect 3880 3040 3920 3050
rect 4320 3040 4360 3050
rect 4400 3040 4520 3050
rect 4880 3040 5000 3050
rect 5120 3040 5200 3050
rect 8400 3040 8440 3050
rect 8720 3040 8920 3050
rect 9480 3040 9520 3050
rect 9760 3040 9800 3050
rect 9880 3040 9960 3050
rect 2040 3030 2120 3040
rect 3120 3030 3160 3040
rect 3880 3030 3920 3040
rect 4320 3030 4360 3040
rect 4400 3030 4520 3040
rect 4880 3030 5000 3040
rect 5120 3030 5200 3040
rect 8400 3030 8440 3040
rect 8720 3030 8920 3040
rect 9480 3030 9520 3040
rect 9760 3030 9800 3040
rect 9880 3030 9960 3040
rect 2040 3020 2120 3030
rect 3120 3020 3160 3030
rect 3880 3020 3920 3030
rect 4320 3020 4360 3030
rect 4400 3020 4520 3030
rect 4880 3020 5000 3030
rect 5120 3020 5200 3030
rect 8400 3020 8440 3030
rect 8720 3020 8920 3030
rect 9480 3020 9520 3030
rect 9760 3020 9800 3030
rect 9880 3020 9960 3030
rect 2040 3010 2080 3020
rect 3120 3010 3160 3020
rect 3880 3010 3920 3020
rect 4000 3010 4040 3020
rect 4360 3010 4480 3020
rect 4880 3010 5200 3020
rect 8320 3010 8360 3020
rect 8600 3010 8720 3020
rect 8760 3010 8920 3020
rect 9760 3010 9800 3020
rect 9880 3010 9960 3020
rect 2040 3000 2080 3010
rect 3120 3000 3160 3010
rect 3880 3000 3920 3010
rect 4000 3000 4040 3010
rect 4360 3000 4480 3010
rect 4880 3000 5200 3010
rect 8320 3000 8360 3010
rect 8600 3000 8720 3010
rect 8760 3000 8920 3010
rect 9760 3000 9800 3010
rect 9880 3000 9960 3010
rect 2040 2990 2080 3000
rect 3120 2990 3160 3000
rect 3880 2990 3920 3000
rect 4000 2990 4040 3000
rect 4360 2990 4480 3000
rect 4880 2990 5200 3000
rect 8320 2990 8360 3000
rect 8600 2990 8720 3000
rect 8760 2990 8920 3000
rect 9760 2990 9800 3000
rect 9880 2990 9960 3000
rect 2040 2980 2080 2990
rect 3120 2980 3160 2990
rect 3880 2980 3920 2990
rect 4000 2980 4040 2990
rect 4360 2980 4480 2990
rect 4880 2980 5200 2990
rect 8320 2980 8360 2990
rect 8600 2980 8720 2990
rect 8760 2980 8920 2990
rect 9760 2980 9800 2990
rect 9880 2980 9960 2990
rect 2040 2970 2080 2980
rect 3120 2970 3160 2980
rect 3880 2970 3920 2980
rect 4040 2970 4080 2980
rect 4120 2970 4160 2980
rect 4400 2970 4480 2980
rect 4920 2970 5160 2980
rect 8400 2970 8440 2980
rect 8560 2970 8800 2980
rect 8840 2970 8920 2980
rect 9440 2970 9480 2980
rect 9880 2970 9960 2980
rect 2040 2960 2080 2970
rect 3120 2960 3160 2970
rect 3880 2960 3920 2970
rect 4040 2960 4080 2970
rect 4120 2960 4160 2970
rect 4400 2960 4480 2970
rect 4920 2960 5160 2970
rect 8400 2960 8440 2970
rect 8560 2960 8800 2970
rect 8840 2960 8920 2970
rect 9440 2960 9480 2970
rect 9880 2960 9960 2970
rect 2040 2950 2080 2960
rect 3120 2950 3160 2960
rect 3880 2950 3920 2960
rect 4040 2950 4080 2960
rect 4120 2950 4160 2960
rect 4400 2950 4480 2960
rect 4920 2950 5160 2960
rect 8400 2950 8440 2960
rect 8560 2950 8800 2960
rect 8840 2950 8920 2960
rect 9440 2950 9480 2960
rect 9880 2950 9960 2960
rect 2040 2940 2080 2950
rect 3120 2940 3160 2950
rect 3880 2940 3920 2950
rect 4040 2940 4080 2950
rect 4120 2940 4160 2950
rect 4400 2940 4480 2950
rect 4920 2940 5160 2950
rect 8400 2940 8440 2950
rect 8560 2940 8800 2950
rect 8840 2940 8920 2950
rect 9440 2940 9480 2950
rect 9880 2940 9960 2950
rect 2040 2930 2080 2940
rect 4440 2930 4520 2940
rect 4920 2930 5160 2940
rect 8520 2930 8680 2940
rect 9400 2930 9440 2940
rect 9680 2930 9720 2940
rect 9920 2930 9960 2940
rect 2040 2920 2080 2930
rect 4440 2920 4520 2930
rect 4920 2920 5160 2930
rect 8520 2920 8680 2930
rect 9400 2920 9440 2930
rect 9680 2920 9720 2930
rect 9920 2920 9960 2930
rect 2040 2910 2080 2920
rect 4440 2910 4520 2920
rect 4920 2910 5160 2920
rect 8520 2910 8680 2920
rect 9400 2910 9440 2920
rect 9680 2910 9720 2920
rect 9920 2910 9960 2920
rect 2040 2900 2080 2910
rect 4440 2900 4520 2910
rect 4920 2900 5160 2910
rect 8520 2900 8680 2910
rect 9400 2900 9440 2910
rect 9680 2900 9720 2910
rect 9920 2900 9960 2910
rect 2000 2890 2080 2900
rect 8240 2890 8280 2900
rect 8520 2890 8640 2900
rect 8720 2890 8800 2900
rect 9120 2890 9200 2900
rect 9360 2890 9400 2900
rect 9680 2890 9720 2900
rect 9920 2890 9990 2900
rect 2000 2880 2080 2890
rect 8240 2880 8280 2890
rect 8520 2880 8640 2890
rect 8720 2880 8800 2890
rect 9120 2880 9200 2890
rect 9360 2880 9400 2890
rect 9680 2880 9720 2890
rect 9920 2880 9990 2890
rect 2000 2870 2080 2880
rect 8240 2870 8280 2880
rect 8520 2870 8640 2880
rect 8720 2870 8800 2880
rect 9120 2870 9200 2880
rect 9360 2870 9400 2880
rect 9680 2870 9720 2880
rect 9920 2870 9990 2880
rect 2000 2860 2080 2870
rect 8240 2860 8280 2870
rect 8520 2860 8640 2870
rect 8720 2860 8800 2870
rect 9120 2860 9200 2870
rect 9360 2860 9400 2870
rect 9680 2860 9720 2870
rect 9920 2860 9990 2870
rect 2000 2850 2040 2860
rect 3080 2850 3160 2860
rect 8520 2850 8640 2860
rect 8840 2850 8880 2860
rect 9080 2850 9200 2860
rect 9360 2850 9400 2860
rect 9920 2850 9990 2860
rect 2000 2840 2040 2850
rect 3080 2840 3160 2850
rect 8520 2840 8640 2850
rect 8840 2840 8880 2850
rect 9080 2840 9200 2850
rect 9360 2840 9400 2850
rect 9920 2840 9990 2850
rect 2000 2830 2040 2840
rect 3080 2830 3160 2840
rect 8520 2830 8640 2840
rect 8840 2830 8880 2840
rect 9080 2830 9200 2840
rect 9360 2830 9400 2840
rect 9920 2830 9990 2840
rect 2000 2820 2040 2830
rect 3080 2820 3160 2830
rect 8520 2820 8640 2830
rect 8840 2820 8880 2830
rect 9080 2820 9200 2830
rect 9360 2820 9400 2830
rect 9920 2820 9990 2830
rect 2000 2810 2080 2820
rect 2240 2810 2400 2820
rect 2840 2810 3120 2820
rect 3960 2810 4000 2820
rect 4240 2810 4280 2820
rect 7160 2810 7200 2820
rect 8520 2810 8640 2820
rect 8720 2810 8800 2820
rect 9040 2810 9160 2820
rect 9200 2810 9280 2820
rect 9320 2810 9400 2820
rect 9440 2810 9480 2820
rect 9560 2810 9680 2820
rect 9920 2810 9990 2820
rect 2000 2800 2080 2810
rect 2240 2800 2400 2810
rect 2840 2800 3120 2810
rect 3960 2800 4000 2810
rect 4240 2800 4280 2810
rect 7160 2800 7200 2810
rect 8520 2800 8640 2810
rect 8720 2800 8800 2810
rect 9040 2800 9160 2810
rect 9200 2800 9280 2810
rect 9320 2800 9400 2810
rect 9440 2800 9480 2810
rect 9560 2800 9680 2810
rect 9920 2800 9990 2810
rect 2000 2790 2080 2800
rect 2240 2790 2400 2800
rect 2840 2790 3120 2800
rect 3960 2790 4000 2800
rect 4240 2790 4280 2800
rect 7160 2790 7200 2800
rect 8520 2790 8640 2800
rect 8720 2790 8800 2800
rect 9040 2790 9160 2800
rect 9200 2790 9280 2800
rect 9320 2790 9400 2800
rect 9440 2790 9480 2800
rect 9560 2790 9680 2800
rect 9920 2790 9990 2800
rect 2000 2780 2080 2790
rect 2240 2780 2400 2790
rect 2840 2780 3120 2790
rect 3960 2780 4000 2790
rect 4240 2780 4280 2790
rect 7160 2780 7200 2790
rect 8520 2780 8640 2790
rect 8720 2780 8800 2790
rect 9040 2780 9160 2790
rect 9200 2780 9280 2790
rect 9320 2780 9400 2790
rect 9440 2780 9480 2790
rect 9560 2780 9680 2790
rect 9920 2780 9990 2790
rect 2040 2770 2080 2780
rect 2200 2770 2440 2780
rect 2800 2770 3040 2780
rect 3080 2770 3120 2780
rect 3920 2770 3960 2780
rect 4160 2770 4200 2780
rect 4240 2770 4280 2780
rect 7080 2770 7120 2780
rect 7600 2770 7640 2780
rect 8560 2770 8640 2780
rect 9200 2770 9280 2780
rect 9400 2770 9480 2780
rect 9520 2770 9560 2780
rect 9600 2770 9640 2780
rect 9680 2770 9720 2780
rect 9880 2770 9920 2780
rect 2040 2760 2080 2770
rect 2200 2760 2440 2770
rect 2800 2760 3040 2770
rect 3080 2760 3120 2770
rect 3920 2760 3960 2770
rect 4160 2760 4200 2770
rect 4240 2760 4280 2770
rect 7080 2760 7120 2770
rect 7600 2760 7640 2770
rect 8560 2760 8640 2770
rect 9200 2760 9280 2770
rect 9400 2760 9480 2770
rect 9520 2760 9560 2770
rect 9600 2760 9640 2770
rect 9680 2760 9720 2770
rect 9880 2760 9920 2770
rect 2040 2750 2080 2760
rect 2200 2750 2440 2760
rect 2800 2750 3040 2760
rect 3080 2750 3120 2760
rect 3920 2750 3960 2760
rect 4160 2750 4200 2760
rect 4240 2750 4280 2760
rect 7080 2750 7120 2760
rect 7600 2750 7640 2760
rect 8560 2750 8640 2760
rect 9200 2750 9280 2760
rect 9400 2750 9480 2760
rect 9520 2750 9560 2760
rect 9600 2750 9640 2760
rect 9680 2750 9720 2760
rect 9880 2750 9920 2760
rect 2040 2740 2080 2750
rect 2200 2740 2440 2750
rect 2800 2740 3040 2750
rect 3080 2740 3120 2750
rect 3920 2740 3960 2750
rect 4160 2740 4200 2750
rect 4240 2740 4280 2750
rect 7080 2740 7120 2750
rect 7600 2740 7640 2750
rect 8560 2740 8640 2750
rect 9200 2740 9280 2750
rect 9400 2740 9480 2750
rect 9520 2740 9560 2750
rect 9600 2740 9640 2750
rect 9680 2740 9720 2750
rect 9880 2740 9920 2750
rect 2040 2730 2080 2740
rect 2280 2730 2480 2740
rect 2760 2730 2960 2740
rect 3120 2730 3160 2740
rect 3920 2730 3960 2740
rect 4240 2730 4280 2740
rect 7000 2730 7040 2740
rect 8120 2730 8160 2740
rect 8560 2730 8640 2740
rect 9280 2730 9320 2740
rect 9360 2730 9400 2740
rect 9560 2730 9640 2740
rect 9680 2730 9720 2740
rect 9880 2730 9920 2740
rect 2040 2720 2080 2730
rect 2280 2720 2480 2730
rect 2760 2720 2960 2730
rect 3120 2720 3160 2730
rect 3920 2720 3960 2730
rect 4240 2720 4280 2730
rect 7000 2720 7040 2730
rect 8120 2720 8160 2730
rect 8560 2720 8640 2730
rect 9280 2720 9320 2730
rect 9360 2720 9400 2730
rect 9560 2720 9640 2730
rect 9680 2720 9720 2730
rect 9880 2720 9920 2730
rect 2040 2710 2080 2720
rect 2280 2710 2480 2720
rect 2760 2710 2960 2720
rect 3120 2710 3160 2720
rect 3920 2710 3960 2720
rect 4240 2710 4280 2720
rect 7000 2710 7040 2720
rect 8120 2710 8160 2720
rect 8560 2710 8640 2720
rect 9280 2710 9320 2720
rect 9360 2710 9400 2720
rect 9560 2710 9640 2720
rect 9680 2710 9720 2720
rect 9880 2710 9920 2720
rect 2040 2700 2080 2710
rect 2280 2700 2480 2710
rect 2760 2700 2960 2710
rect 3120 2700 3160 2710
rect 3920 2700 3960 2710
rect 4240 2700 4280 2710
rect 7000 2700 7040 2710
rect 8120 2700 8160 2710
rect 8560 2700 8640 2710
rect 9280 2700 9320 2710
rect 9360 2700 9400 2710
rect 9560 2700 9640 2710
rect 9680 2700 9720 2710
rect 9880 2700 9920 2710
rect 2000 2690 2040 2700
rect 2200 2690 2280 2700
rect 2320 2690 2480 2700
rect 2760 2690 2800 2700
rect 2840 2690 2920 2700
rect 2960 2690 3120 2700
rect 4200 2690 4280 2700
rect 8080 2690 8120 2700
rect 8560 2690 8640 2700
rect 9240 2690 9280 2700
rect 9680 2690 9720 2700
rect 9920 2690 9960 2700
rect 2000 2680 2040 2690
rect 2200 2680 2280 2690
rect 2320 2680 2480 2690
rect 2760 2680 2800 2690
rect 2840 2680 2920 2690
rect 2960 2680 3120 2690
rect 4200 2680 4280 2690
rect 8080 2680 8120 2690
rect 8560 2680 8640 2690
rect 9240 2680 9280 2690
rect 9680 2680 9720 2690
rect 9920 2680 9960 2690
rect 2000 2670 2040 2680
rect 2200 2670 2280 2680
rect 2320 2670 2480 2680
rect 2760 2670 2800 2680
rect 2840 2670 2920 2680
rect 2960 2670 3120 2680
rect 4200 2670 4280 2680
rect 8080 2670 8120 2680
rect 8560 2670 8640 2680
rect 9240 2670 9280 2680
rect 9680 2670 9720 2680
rect 9920 2670 9960 2680
rect 2000 2660 2040 2670
rect 2200 2660 2280 2670
rect 2320 2660 2480 2670
rect 2760 2660 2800 2670
rect 2840 2660 2920 2670
rect 2960 2660 3120 2670
rect 4200 2660 4280 2670
rect 8080 2660 8120 2670
rect 8560 2660 8640 2670
rect 9240 2660 9280 2670
rect 9680 2660 9720 2670
rect 9920 2660 9960 2670
rect 2000 2650 2120 2660
rect 2440 2650 2480 2660
rect 2720 2650 2760 2660
rect 2960 2650 3040 2660
rect 4240 2650 4280 2660
rect 7160 2650 7200 2660
rect 7680 2650 7720 2660
rect 8040 2650 8080 2660
rect 8520 2650 8560 2660
rect 8600 2650 8880 2660
rect 9200 2650 9240 2660
rect 9760 2650 9800 2660
rect 9840 2650 9960 2660
rect 2000 2640 2120 2650
rect 2440 2640 2480 2650
rect 2720 2640 2760 2650
rect 2960 2640 3040 2650
rect 4240 2640 4280 2650
rect 7160 2640 7200 2650
rect 7680 2640 7720 2650
rect 8040 2640 8080 2650
rect 8520 2640 8560 2650
rect 8600 2640 8880 2650
rect 9200 2640 9240 2650
rect 9760 2640 9800 2650
rect 9840 2640 9960 2650
rect 2000 2630 2120 2640
rect 2440 2630 2480 2640
rect 2720 2630 2760 2640
rect 2960 2630 3040 2640
rect 4240 2630 4280 2640
rect 7160 2630 7200 2640
rect 7680 2630 7720 2640
rect 8040 2630 8080 2640
rect 8520 2630 8560 2640
rect 8600 2630 8880 2640
rect 9200 2630 9240 2640
rect 9760 2630 9800 2640
rect 9840 2630 9960 2640
rect 2000 2620 2120 2630
rect 2440 2620 2480 2630
rect 2720 2620 2760 2630
rect 2960 2620 3040 2630
rect 4240 2620 4280 2630
rect 7160 2620 7200 2630
rect 7680 2620 7720 2630
rect 8040 2620 8080 2630
rect 8520 2620 8560 2630
rect 8600 2620 8880 2630
rect 9200 2620 9240 2630
rect 9760 2620 9800 2630
rect 9840 2620 9960 2630
rect 1960 2610 2040 2620
rect 2440 2610 2480 2620
rect 2720 2610 2760 2620
rect 3920 2610 3960 2620
rect 4240 2610 4280 2620
rect 7120 2610 7280 2620
rect 8000 2610 8040 2620
rect 8400 2610 8480 2620
rect 8560 2610 8880 2620
rect 1960 2600 2040 2610
rect 2440 2600 2480 2610
rect 2720 2600 2760 2610
rect 3920 2600 3960 2610
rect 4240 2600 4280 2610
rect 7120 2600 7280 2610
rect 8000 2600 8040 2610
rect 8400 2600 8480 2610
rect 8560 2600 8880 2610
rect 1960 2590 2040 2600
rect 2440 2590 2480 2600
rect 2720 2590 2760 2600
rect 3920 2590 3960 2600
rect 4240 2590 4280 2600
rect 7120 2590 7280 2600
rect 8000 2590 8040 2600
rect 8400 2590 8480 2600
rect 8560 2590 8880 2600
rect 1960 2580 2040 2590
rect 2440 2580 2480 2590
rect 2720 2580 2760 2590
rect 3920 2580 3960 2590
rect 4240 2580 4280 2590
rect 7120 2580 7280 2590
rect 8000 2580 8040 2590
rect 8400 2580 8480 2590
rect 8560 2580 8880 2590
rect 1960 2570 2000 2580
rect 2400 2570 2440 2580
rect 2720 2570 2840 2580
rect 3960 2570 4000 2580
rect 4040 2570 4120 2580
rect 7120 2570 7240 2580
rect 7280 2570 7320 2580
rect 7960 2570 8000 2580
rect 8400 2570 8880 2580
rect 8920 2570 9000 2580
rect 9160 2570 9200 2580
rect 9360 2570 9600 2580
rect 1960 2560 2000 2570
rect 2400 2560 2440 2570
rect 2720 2560 2840 2570
rect 3960 2560 4000 2570
rect 4040 2560 4120 2570
rect 7120 2560 7240 2570
rect 7280 2560 7320 2570
rect 7960 2560 8000 2570
rect 8400 2560 8880 2570
rect 8920 2560 9000 2570
rect 9160 2560 9200 2570
rect 9360 2560 9600 2570
rect 1960 2550 2000 2560
rect 2400 2550 2440 2560
rect 2720 2550 2840 2560
rect 3960 2550 4000 2560
rect 4040 2550 4120 2560
rect 7120 2550 7240 2560
rect 7280 2550 7320 2560
rect 7960 2550 8000 2560
rect 8400 2550 8880 2560
rect 8920 2550 9000 2560
rect 9160 2550 9200 2560
rect 9360 2550 9600 2560
rect 1960 2540 2000 2550
rect 2400 2540 2440 2550
rect 2720 2540 2840 2550
rect 3960 2540 4000 2550
rect 4040 2540 4120 2550
rect 7120 2540 7240 2550
rect 7280 2540 7320 2550
rect 7960 2540 8000 2550
rect 8400 2540 8880 2550
rect 8920 2540 9000 2550
rect 9160 2540 9200 2550
rect 9360 2540 9600 2550
rect 2120 2530 2160 2540
rect 2360 2530 2400 2540
rect 2840 2530 2920 2540
rect 3080 2530 3160 2540
rect 4000 2530 4080 2540
rect 7200 2530 7240 2540
rect 7320 2530 7360 2540
rect 7920 2530 7960 2540
rect 8400 2530 9000 2540
rect 9280 2530 9360 2540
rect 9600 2530 9680 2540
rect 2120 2520 2160 2530
rect 2360 2520 2400 2530
rect 2840 2520 2920 2530
rect 3080 2520 3160 2530
rect 4000 2520 4080 2530
rect 7200 2520 7240 2530
rect 7320 2520 7360 2530
rect 7920 2520 7960 2530
rect 8400 2520 9000 2530
rect 9280 2520 9360 2530
rect 9600 2520 9680 2530
rect 2120 2510 2160 2520
rect 2360 2510 2400 2520
rect 2840 2510 2920 2520
rect 3080 2510 3160 2520
rect 4000 2510 4080 2520
rect 7200 2510 7240 2520
rect 7320 2510 7360 2520
rect 7920 2510 7960 2520
rect 8400 2510 9000 2520
rect 9280 2510 9360 2520
rect 9600 2510 9680 2520
rect 2120 2500 2160 2510
rect 2360 2500 2400 2510
rect 2840 2500 2920 2510
rect 3080 2500 3160 2510
rect 4000 2500 4080 2510
rect 7200 2500 7240 2510
rect 7320 2500 7360 2510
rect 7920 2500 7960 2510
rect 8400 2500 9000 2510
rect 9280 2500 9360 2510
rect 9600 2500 9680 2510
rect 2200 2490 2320 2500
rect 3040 2490 3120 2500
rect 6760 2490 6880 2500
rect 7240 2490 7280 2500
rect 7800 2490 7880 2500
rect 8400 2490 8960 2500
rect 9120 2490 9160 2500
rect 9240 2490 9280 2500
rect 9680 2490 9720 2500
rect 2200 2480 2320 2490
rect 3040 2480 3120 2490
rect 6760 2480 6880 2490
rect 7240 2480 7280 2490
rect 7800 2480 7880 2490
rect 8400 2480 8960 2490
rect 9120 2480 9160 2490
rect 9240 2480 9280 2490
rect 9680 2480 9720 2490
rect 2200 2470 2320 2480
rect 3040 2470 3120 2480
rect 6760 2470 6880 2480
rect 7240 2470 7280 2480
rect 7800 2470 7880 2480
rect 8400 2470 8960 2480
rect 9120 2470 9160 2480
rect 9240 2470 9280 2480
rect 9680 2470 9720 2480
rect 2200 2460 2320 2470
rect 3040 2460 3120 2470
rect 6760 2460 6880 2470
rect 7240 2460 7280 2470
rect 7800 2460 7880 2470
rect 8400 2460 8960 2470
rect 9120 2460 9160 2470
rect 9240 2460 9280 2470
rect 9680 2460 9720 2470
rect 1920 2450 1960 2460
rect 2080 2450 2280 2460
rect 3200 2450 3240 2460
rect 6800 2450 6880 2460
rect 7280 2450 7320 2460
rect 7400 2450 7440 2460
rect 8400 2450 9160 2460
rect 9200 2450 9280 2460
rect 9760 2450 9800 2460
rect 1920 2440 1960 2450
rect 2080 2440 2280 2450
rect 3200 2440 3240 2450
rect 6800 2440 6880 2450
rect 7280 2440 7320 2450
rect 7400 2440 7440 2450
rect 8400 2440 9160 2450
rect 9200 2440 9280 2450
rect 9760 2440 9800 2450
rect 1920 2430 1960 2440
rect 2080 2430 2280 2440
rect 3200 2430 3240 2440
rect 6800 2430 6880 2440
rect 7280 2430 7320 2440
rect 7400 2430 7440 2440
rect 8400 2430 9160 2440
rect 9200 2430 9280 2440
rect 9760 2430 9800 2440
rect 1920 2420 1960 2430
rect 2080 2420 2280 2430
rect 3200 2420 3240 2430
rect 6800 2420 6880 2430
rect 7280 2420 7320 2430
rect 7400 2420 7440 2430
rect 8400 2420 9160 2430
rect 9200 2420 9280 2430
rect 9760 2420 9800 2430
rect 1920 2410 1960 2420
rect 3200 2410 3240 2420
rect 6880 2410 6960 2420
rect 7440 2410 7480 2420
rect 8400 2410 9200 2420
rect 9240 2410 9280 2420
rect 9480 2410 9560 2420
rect 9800 2410 9840 2420
rect 1920 2400 1960 2410
rect 3200 2400 3240 2410
rect 6880 2400 6960 2410
rect 7440 2400 7480 2410
rect 8400 2400 9200 2410
rect 9240 2400 9280 2410
rect 9480 2400 9560 2410
rect 9800 2400 9840 2410
rect 1920 2390 1960 2400
rect 3200 2390 3240 2400
rect 6880 2390 6960 2400
rect 7440 2390 7480 2400
rect 8400 2390 9200 2400
rect 9240 2390 9280 2400
rect 9480 2390 9560 2400
rect 9800 2390 9840 2400
rect 1920 2380 1960 2390
rect 3200 2380 3240 2390
rect 6880 2380 6960 2390
rect 7440 2380 7480 2390
rect 8400 2380 9200 2390
rect 9240 2380 9280 2390
rect 9480 2380 9560 2390
rect 9800 2380 9840 2390
rect 1920 2370 1960 2380
rect 6920 2370 7120 2380
rect 7400 2370 7440 2380
rect 7480 2370 7520 2380
rect 8440 2370 8680 2380
rect 8760 2370 9160 2380
rect 9200 2370 9280 2380
rect 9480 2370 9560 2380
rect 9800 2370 9840 2380
rect 1920 2360 1960 2370
rect 6920 2360 7120 2370
rect 7400 2360 7440 2370
rect 7480 2360 7520 2370
rect 8440 2360 8680 2370
rect 8760 2360 9160 2370
rect 9200 2360 9280 2370
rect 9480 2360 9560 2370
rect 9800 2360 9840 2370
rect 1920 2350 1960 2360
rect 6920 2350 7120 2360
rect 7400 2350 7440 2360
rect 7480 2350 7520 2360
rect 8440 2350 8680 2360
rect 8760 2350 9160 2360
rect 9200 2350 9280 2360
rect 9480 2350 9560 2360
rect 9800 2350 9840 2360
rect 1920 2340 1960 2350
rect 6920 2340 7120 2350
rect 7400 2340 7440 2350
rect 7480 2340 7520 2350
rect 8440 2340 8680 2350
rect 8760 2340 9160 2350
rect 9200 2340 9280 2350
rect 9480 2340 9560 2350
rect 9800 2340 9840 2350
rect 1880 2330 1920 2340
rect 3240 2330 3280 2340
rect 7040 2330 7200 2340
rect 7520 2330 7560 2340
rect 8360 2330 8400 2340
rect 8560 2330 8640 2340
rect 8760 2330 8840 2340
rect 8960 2330 9160 2340
rect 9480 2330 9560 2340
rect 9800 2330 9840 2340
rect 1880 2320 1920 2330
rect 3240 2320 3280 2330
rect 7040 2320 7200 2330
rect 7520 2320 7560 2330
rect 8360 2320 8400 2330
rect 8560 2320 8640 2330
rect 8760 2320 8840 2330
rect 8960 2320 9160 2330
rect 9480 2320 9560 2330
rect 9800 2320 9840 2330
rect 1880 2310 1920 2320
rect 3240 2310 3280 2320
rect 7040 2310 7200 2320
rect 7520 2310 7560 2320
rect 8360 2310 8400 2320
rect 8560 2310 8640 2320
rect 8760 2310 8840 2320
rect 8960 2310 9160 2320
rect 9480 2310 9560 2320
rect 9800 2310 9840 2320
rect 1880 2300 1920 2310
rect 3240 2300 3280 2310
rect 7040 2300 7200 2310
rect 7520 2300 7560 2310
rect 8360 2300 8400 2310
rect 8560 2300 8640 2310
rect 8760 2300 8840 2310
rect 8960 2300 9160 2310
rect 9480 2300 9560 2310
rect 9800 2300 9840 2310
rect 1880 2290 1920 2300
rect 3240 2290 3280 2300
rect 7240 2290 7400 2300
rect 7480 2290 7520 2300
rect 7600 2290 7640 2300
rect 8600 2290 8680 2300
rect 8720 2290 9120 2300
rect 9800 2290 9840 2300
rect 1880 2280 1920 2290
rect 3240 2280 3280 2290
rect 7240 2280 7400 2290
rect 7480 2280 7520 2290
rect 7600 2280 7640 2290
rect 8600 2280 8680 2290
rect 8720 2280 9120 2290
rect 9800 2280 9840 2290
rect 1880 2270 1920 2280
rect 3240 2270 3280 2280
rect 7240 2270 7400 2280
rect 7480 2270 7520 2280
rect 7600 2270 7640 2280
rect 8600 2270 8680 2280
rect 8720 2270 9120 2280
rect 9800 2270 9840 2280
rect 1880 2260 1920 2270
rect 3240 2260 3280 2270
rect 7240 2260 7400 2270
rect 7480 2260 7520 2270
rect 7600 2260 7640 2270
rect 8600 2260 8680 2270
rect 8720 2260 9120 2270
rect 9800 2260 9840 2270
rect 1880 2250 1920 2260
rect 2680 2250 2720 2260
rect 3240 2250 3280 2260
rect 6400 2250 6440 2260
rect 6760 2250 6800 2260
rect 7480 2250 7520 2260
rect 8680 2250 8720 2260
rect 8800 2250 8880 2260
rect 9000 2250 9080 2260
rect 9240 2250 9320 2260
rect 1880 2240 1920 2250
rect 2680 2240 2720 2250
rect 3240 2240 3280 2250
rect 6400 2240 6440 2250
rect 6760 2240 6800 2250
rect 7480 2240 7520 2250
rect 8680 2240 8720 2250
rect 8800 2240 8880 2250
rect 9000 2240 9080 2250
rect 9240 2240 9320 2250
rect 1880 2230 1920 2240
rect 2680 2230 2720 2240
rect 3240 2230 3280 2240
rect 6400 2230 6440 2240
rect 6760 2230 6800 2240
rect 7480 2230 7520 2240
rect 8680 2230 8720 2240
rect 8800 2230 8880 2240
rect 9000 2230 9080 2240
rect 9240 2230 9320 2240
rect 1880 2220 1920 2230
rect 2680 2220 2720 2230
rect 3240 2220 3280 2230
rect 6400 2220 6440 2230
rect 6760 2220 6800 2230
rect 7480 2220 7520 2230
rect 8680 2220 8720 2230
rect 8800 2220 8880 2230
rect 9000 2220 9080 2230
rect 9240 2220 9320 2230
rect 1880 2210 1920 2220
rect 2440 2210 2600 2220
rect 2720 2210 2840 2220
rect 3240 2210 3280 2220
rect 6400 2210 6440 2220
rect 6760 2210 6800 2220
rect 7480 2210 7520 2220
rect 7680 2210 7720 2220
rect 9320 2210 9400 2220
rect 9800 2210 9840 2220
rect 9960 2210 9990 2220
rect 1880 2200 1920 2210
rect 2440 2200 2600 2210
rect 2720 2200 2840 2210
rect 3240 2200 3280 2210
rect 6400 2200 6440 2210
rect 6760 2200 6800 2210
rect 7480 2200 7520 2210
rect 7680 2200 7720 2210
rect 9320 2200 9400 2210
rect 9800 2200 9840 2210
rect 9960 2200 9990 2210
rect 1880 2190 1920 2200
rect 2440 2190 2600 2200
rect 2720 2190 2840 2200
rect 3240 2190 3280 2200
rect 6400 2190 6440 2200
rect 6760 2190 6800 2200
rect 7480 2190 7520 2200
rect 7680 2190 7720 2200
rect 9320 2190 9400 2200
rect 9800 2190 9840 2200
rect 9960 2190 9990 2200
rect 1880 2180 1920 2190
rect 2440 2180 2600 2190
rect 2720 2180 2840 2190
rect 3240 2180 3280 2190
rect 6400 2180 6440 2190
rect 6760 2180 6800 2190
rect 7480 2180 7520 2190
rect 7680 2180 7720 2190
rect 9320 2180 9400 2190
rect 9800 2180 9840 2190
rect 9960 2180 9990 2190
rect 1880 2170 1920 2180
rect 2240 2170 2280 2180
rect 2360 2170 2400 2180
rect 2800 2170 2840 2180
rect 3240 2170 3280 2180
rect 6400 2170 6480 2180
rect 6760 2170 6840 2180
rect 7760 2170 7840 2180
rect 9240 2170 9280 2180
rect 9400 2170 9480 2180
rect 9760 2170 9800 2180
rect 1880 2160 1920 2170
rect 2240 2160 2280 2170
rect 2360 2160 2400 2170
rect 2800 2160 2840 2170
rect 3240 2160 3280 2170
rect 6400 2160 6480 2170
rect 6760 2160 6840 2170
rect 7760 2160 7840 2170
rect 9240 2160 9280 2170
rect 9400 2160 9480 2170
rect 9760 2160 9800 2170
rect 1880 2150 1920 2160
rect 2240 2150 2280 2160
rect 2360 2150 2400 2160
rect 2800 2150 2840 2160
rect 3240 2150 3280 2160
rect 6400 2150 6480 2160
rect 6760 2150 6840 2160
rect 7760 2150 7840 2160
rect 9240 2150 9280 2160
rect 9400 2150 9480 2160
rect 9760 2150 9800 2160
rect 1880 2140 1920 2150
rect 2240 2140 2280 2150
rect 2360 2140 2400 2150
rect 2800 2140 2840 2150
rect 3240 2140 3280 2150
rect 6400 2140 6480 2150
rect 6760 2140 6840 2150
rect 7760 2140 7840 2150
rect 9240 2140 9280 2150
rect 9400 2140 9480 2150
rect 9760 2140 9800 2150
rect 1880 2130 1920 2140
rect 2200 2130 2280 2140
rect 2360 2130 2560 2140
rect 2640 2130 2800 2140
rect 3240 2130 3280 2140
rect 6360 2130 6480 2140
rect 6800 2130 6880 2140
rect 7840 2130 7880 2140
rect 8360 2130 8400 2140
rect 9320 2130 9360 2140
rect 9480 2130 9640 2140
rect 9680 2130 9760 2140
rect 1880 2120 1920 2130
rect 2200 2120 2280 2130
rect 2360 2120 2560 2130
rect 2640 2120 2800 2130
rect 3240 2120 3280 2130
rect 6360 2120 6480 2130
rect 6800 2120 6880 2130
rect 7840 2120 7880 2130
rect 8360 2120 8400 2130
rect 9320 2120 9360 2130
rect 9480 2120 9640 2130
rect 9680 2120 9760 2130
rect 1880 2110 1920 2120
rect 2200 2110 2280 2120
rect 2360 2110 2560 2120
rect 2640 2110 2800 2120
rect 3240 2110 3280 2120
rect 6360 2110 6480 2120
rect 6800 2110 6880 2120
rect 7840 2110 7880 2120
rect 8360 2110 8400 2120
rect 9320 2110 9360 2120
rect 9480 2110 9640 2120
rect 9680 2110 9760 2120
rect 1880 2100 1920 2110
rect 2200 2100 2280 2110
rect 2360 2100 2560 2110
rect 2640 2100 2800 2110
rect 3240 2100 3280 2110
rect 6360 2100 6480 2110
rect 6800 2100 6880 2110
rect 7840 2100 7880 2110
rect 8360 2100 8400 2110
rect 9320 2100 9360 2110
rect 9480 2100 9640 2110
rect 9680 2100 9760 2110
rect 1880 2090 1960 2100
rect 2200 2090 2240 2100
rect 3200 2090 3280 2100
rect 6400 2090 6480 2100
rect 6800 2090 6920 2100
rect 7280 2090 7320 2100
rect 7880 2090 7920 2100
rect 8360 2090 8400 2100
rect 9240 2090 9280 2100
rect 9320 2090 9480 2100
rect 9680 2090 9720 2100
rect 1880 2080 1960 2090
rect 2200 2080 2240 2090
rect 3200 2080 3280 2090
rect 6400 2080 6480 2090
rect 6800 2080 6920 2090
rect 7280 2080 7320 2090
rect 7880 2080 7920 2090
rect 8360 2080 8400 2090
rect 9240 2080 9280 2090
rect 9320 2080 9480 2090
rect 9680 2080 9720 2090
rect 1880 2070 1960 2080
rect 2200 2070 2240 2080
rect 3200 2070 3280 2080
rect 6400 2070 6480 2080
rect 6800 2070 6920 2080
rect 7280 2070 7320 2080
rect 7880 2070 7920 2080
rect 8360 2070 8400 2080
rect 9240 2070 9280 2080
rect 9320 2070 9480 2080
rect 9680 2070 9720 2080
rect 1880 2060 1960 2070
rect 2200 2060 2240 2070
rect 3200 2060 3280 2070
rect 6400 2060 6480 2070
rect 6800 2060 6920 2070
rect 7280 2060 7320 2070
rect 7880 2060 7920 2070
rect 8360 2060 8400 2070
rect 9240 2060 9280 2070
rect 9320 2060 9480 2070
rect 9680 2060 9720 2070
rect 1880 2050 2000 2060
rect 2120 2050 2200 2060
rect 3160 2050 3240 2060
rect 6360 2050 6480 2060
rect 6800 2050 6960 2060
rect 7280 2050 7320 2060
rect 8360 2050 8400 2060
rect 9600 2050 9680 2060
rect 1880 2040 2000 2050
rect 2120 2040 2200 2050
rect 3160 2040 3240 2050
rect 6360 2040 6480 2050
rect 6800 2040 6960 2050
rect 7280 2040 7320 2050
rect 8360 2040 8400 2050
rect 9600 2040 9680 2050
rect 1880 2030 2000 2040
rect 2120 2030 2200 2040
rect 3160 2030 3240 2040
rect 6360 2030 6480 2040
rect 6800 2030 6960 2040
rect 7280 2030 7320 2040
rect 8360 2030 8400 2040
rect 9600 2030 9680 2040
rect 1880 2020 2000 2030
rect 2120 2020 2200 2030
rect 3160 2020 3240 2030
rect 6360 2020 6480 2030
rect 6800 2020 6960 2030
rect 7280 2020 7320 2030
rect 8360 2020 8400 2030
rect 9600 2020 9680 2030
rect 1880 2010 2200 2020
rect 3120 2010 3240 2020
rect 6360 2010 6480 2020
rect 6840 2010 7040 2020
rect 7280 2010 7320 2020
rect 7960 2010 8000 2020
rect 8360 2010 8400 2020
rect 8440 2010 8520 2020
rect 9080 2010 9200 2020
rect 1880 2000 2200 2010
rect 3120 2000 3240 2010
rect 6360 2000 6480 2010
rect 6840 2000 7040 2010
rect 7280 2000 7320 2010
rect 7960 2000 8000 2010
rect 8360 2000 8400 2010
rect 8440 2000 8520 2010
rect 9080 2000 9200 2010
rect 1880 1990 2200 2000
rect 3120 1990 3240 2000
rect 6360 1990 6480 2000
rect 6840 1990 7040 2000
rect 7280 1990 7320 2000
rect 7960 1990 8000 2000
rect 8360 1990 8400 2000
rect 8440 1990 8520 2000
rect 9080 1990 9200 2000
rect 1880 1980 2200 1990
rect 3120 1980 3240 1990
rect 6360 1980 6480 1990
rect 6840 1980 7040 1990
rect 7280 1980 7320 1990
rect 7960 1980 8000 1990
rect 8360 1980 8400 1990
rect 8440 1980 8520 1990
rect 9080 1980 9200 1990
rect 1880 1970 2160 1980
rect 3120 1970 3240 1980
rect 6360 1970 6480 1980
rect 6840 1970 7120 1980
rect 7240 1970 7320 1980
rect 8360 1970 8400 1980
rect 8440 1970 8640 1980
rect 9040 1970 9120 1980
rect 9880 1970 9960 1980
rect 1880 1960 2160 1970
rect 3120 1960 3240 1970
rect 6360 1960 6480 1970
rect 6840 1960 7120 1970
rect 7240 1960 7320 1970
rect 8360 1960 8400 1970
rect 8440 1960 8640 1970
rect 9040 1960 9120 1970
rect 9880 1960 9960 1970
rect 1880 1950 2160 1960
rect 3120 1950 3240 1960
rect 6360 1950 6480 1960
rect 6840 1950 7120 1960
rect 7240 1950 7320 1960
rect 8360 1950 8400 1960
rect 8440 1950 8640 1960
rect 9040 1950 9120 1960
rect 9880 1950 9960 1960
rect 1880 1940 2160 1950
rect 3120 1940 3240 1950
rect 6360 1940 6480 1950
rect 6840 1940 7120 1950
rect 7240 1940 7320 1950
rect 8360 1940 8400 1950
rect 8440 1940 8640 1950
rect 9040 1940 9120 1950
rect 9880 1940 9960 1950
rect 1880 1930 2160 1940
rect 2600 1930 2760 1940
rect 3120 1930 3240 1940
rect 4480 1930 4520 1940
rect 4800 1930 4840 1940
rect 6400 1930 6480 1940
rect 6840 1930 7320 1940
rect 7840 1930 7920 1940
rect 8360 1930 8400 1940
rect 8440 1930 8720 1940
rect 8960 1930 9120 1940
rect 9600 1930 9720 1940
rect 9880 1930 9990 1940
rect 1880 1920 2160 1930
rect 2600 1920 2760 1930
rect 3120 1920 3240 1930
rect 4480 1920 4520 1930
rect 4800 1920 4840 1930
rect 6400 1920 6480 1930
rect 6840 1920 7320 1930
rect 7840 1920 7920 1930
rect 8360 1920 8400 1930
rect 8440 1920 8720 1930
rect 8960 1920 9120 1930
rect 9600 1920 9720 1930
rect 9880 1920 9990 1930
rect 1880 1910 2160 1920
rect 2600 1910 2760 1920
rect 3120 1910 3240 1920
rect 4480 1910 4520 1920
rect 4800 1910 4840 1920
rect 6400 1910 6480 1920
rect 6840 1910 7320 1920
rect 7840 1910 7920 1920
rect 8360 1910 8400 1920
rect 8440 1910 8720 1920
rect 8960 1910 9120 1920
rect 9600 1910 9720 1920
rect 9880 1910 9990 1920
rect 1880 1900 2160 1910
rect 2600 1900 2760 1910
rect 3120 1900 3240 1910
rect 4480 1900 4520 1910
rect 4800 1900 4840 1910
rect 6400 1900 6480 1910
rect 6840 1900 7320 1910
rect 7840 1900 7920 1910
rect 8360 1900 8400 1910
rect 8440 1900 8720 1910
rect 8960 1900 9120 1910
rect 9600 1900 9720 1910
rect 9880 1900 9990 1910
rect 1880 1890 2160 1900
rect 2400 1890 2440 1900
rect 2800 1890 3000 1900
rect 3120 1890 3280 1900
rect 4480 1890 4520 1900
rect 5000 1890 5040 1900
rect 5080 1890 5160 1900
rect 6840 1890 7320 1900
rect 7840 1890 7920 1900
rect 8360 1890 8400 1900
rect 8440 1890 8640 1900
rect 9000 1890 9200 1900
rect 9680 1890 9760 1900
rect 1880 1880 2160 1890
rect 2400 1880 2440 1890
rect 2800 1880 3000 1890
rect 3120 1880 3280 1890
rect 4480 1880 4520 1890
rect 5000 1880 5040 1890
rect 5080 1880 5160 1890
rect 6840 1880 7320 1890
rect 7840 1880 7920 1890
rect 8360 1880 8400 1890
rect 8440 1880 8640 1890
rect 9000 1880 9200 1890
rect 9680 1880 9760 1890
rect 1880 1870 2160 1880
rect 2400 1870 2440 1880
rect 2800 1870 3000 1880
rect 3120 1870 3280 1880
rect 4480 1870 4520 1880
rect 5000 1870 5040 1880
rect 5080 1870 5160 1880
rect 6840 1870 7320 1880
rect 7840 1870 7920 1880
rect 8360 1870 8400 1880
rect 8440 1870 8640 1880
rect 9000 1870 9200 1880
rect 9680 1870 9760 1880
rect 1880 1860 2160 1870
rect 2400 1860 2440 1870
rect 2800 1860 3000 1870
rect 3120 1860 3280 1870
rect 4480 1860 4520 1870
rect 5000 1860 5040 1870
rect 5080 1860 5160 1870
rect 6840 1860 7320 1870
rect 7840 1860 7920 1870
rect 8360 1860 8400 1870
rect 8440 1860 8640 1870
rect 9000 1860 9200 1870
rect 9680 1860 9760 1870
rect 1880 1850 2160 1860
rect 2200 1850 2360 1860
rect 2880 1850 2960 1860
rect 3120 1850 3280 1860
rect 4480 1850 4520 1860
rect 5000 1850 5040 1860
rect 5160 1850 5200 1860
rect 5240 1850 5320 1860
rect 6840 1850 7320 1860
rect 7840 1850 7920 1860
rect 8440 1850 8640 1860
rect 8960 1850 9120 1860
rect 9200 1850 9400 1860
rect 9680 1850 9720 1860
rect 9760 1850 9800 1860
rect 1880 1840 2160 1850
rect 2200 1840 2360 1850
rect 2880 1840 2960 1850
rect 3120 1840 3280 1850
rect 4480 1840 4520 1850
rect 5000 1840 5040 1850
rect 5160 1840 5200 1850
rect 5240 1840 5320 1850
rect 6840 1840 7320 1850
rect 7840 1840 7920 1850
rect 8440 1840 8640 1850
rect 8960 1840 9120 1850
rect 9200 1840 9400 1850
rect 9680 1840 9720 1850
rect 9760 1840 9800 1850
rect 1880 1830 2160 1840
rect 2200 1830 2360 1840
rect 2880 1830 2960 1840
rect 3120 1830 3280 1840
rect 4480 1830 4520 1840
rect 5000 1830 5040 1840
rect 5160 1830 5200 1840
rect 5240 1830 5320 1840
rect 6840 1830 7320 1840
rect 7840 1830 7920 1840
rect 8440 1830 8640 1840
rect 8960 1830 9120 1840
rect 9200 1830 9400 1840
rect 9680 1830 9720 1840
rect 9760 1830 9800 1840
rect 1880 1820 2160 1830
rect 2200 1820 2360 1830
rect 2880 1820 2960 1830
rect 3120 1820 3280 1830
rect 4480 1820 4520 1830
rect 5000 1820 5040 1830
rect 5160 1820 5200 1830
rect 5240 1820 5320 1830
rect 6840 1820 7320 1830
rect 7840 1820 7920 1830
rect 8440 1820 8640 1830
rect 8960 1820 9120 1830
rect 9200 1820 9400 1830
rect 9680 1820 9720 1830
rect 9760 1820 9800 1830
rect 1880 1810 2120 1820
rect 2200 1810 2280 1820
rect 2800 1810 2920 1820
rect 3160 1810 3280 1820
rect 4120 1810 4200 1820
rect 4480 1810 4520 1820
rect 4800 1810 4880 1820
rect 5000 1810 5080 1820
rect 5160 1810 5200 1820
rect 5320 1810 5360 1820
rect 6360 1810 6440 1820
rect 6840 1810 7320 1820
rect 7840 1810 7920 1820
rect 8440 1810 8640 1820
rect 8920 1810 9120 1820
rect 9200 1810 9320 1820
rect 9400 1810 9440 1820
rect 9680 1810 9720 1820
rect 9760 1810 9800 1820
rect 9920 1810 9990 1820
rect 1880 1800 2120 1810
rect 2200 1800 2280 1810
rect 2800 1800 2920 1810
rect 3160 1800 3280 1810
rect 4120 1800 4200 1810
rect 4480 1800 4520 1810
rect 4800 1800 4880 1810
rect 5000 1800 5080 1810
rect 5160 1800 5200 1810
rect 5320 1800 5360 1810
rect 6360 1800 6440 1810
rect 6840 1800 7320 1810
rect 7840 1800 7920 1810
rect 8440 1800 8640 1810
rect 8920 1800 9120 1810
rect 9200 1800 9320 1810
rect 9400 1800 9440 1810
rect 9680 1800 9720 1810
rect 9760 1800 9800 1810
rect 9920 1800 9990 1810
rect 1880 1790 2120 1800
rect 2200 1790 2280 1800
rect 2800 1790 2920 1800
rect 3160 1790 3280 1800
rect 4120 1790 4200 1800
rect 4480 1790 4520 1800
rect 4800 1790 4880 1800
rect 5000 1790 5080 1800
rect 5160 1790 5200 1800
rect 5320 1790 5360 1800
rect 6360 1790 6440 1800
rect 6840 1790 7320 1800
rect 7840 1790 7920 1800
rect 8440 1790 8640 1800
rect 8920 1790 9120 1800
rect 9200 1790 9320 1800
rect 9400 1790 9440 1800
rect 9680 1790 9720 1800
rect 9760 1790 9800 1800
rect 9920 1790 9990 1800
rect 1880 1780 2120 1790
rect 2200 1780 2280 1790
rect 2800 1780 2920 1790
rect 3160 1780 3280 1790
rect 4120 1780 4200 1790
rect 4480 1780 4520 1790
rect 4800 1780 4880 1790
rect 5000 1780 5080 1790
rect 5160 1780 5200 1790
rect 5320 1780 5360 1790
rect 6360 1780 6440 1790
rect 6840 1780 7320 1790
rect 7840 1780 7920 1790
rect 8440 1780 8640 1790
rect 8920 1780 9120 1790
rect 9200 1780 9320 1790
rect 9400 1780 9440 1790
rect 9680 1780 9720 1790
rect 9760 1780 9800 1790
rect 9920 1780 9990 1790
rect 1880 1770 2040 1780
rect 2200 1770 2240 1780
rect 2360 1770 2440 1780
rect 2520 1770 2760 1780
rect 3160 1770 3240 1780
rect 4200 1770 4240 1780
rect 4480 1770 4520 1780
rect 4720 1770 4760 1780
rect 4840 1770 4880 1780
rect 4960 1770 5080 1780
rect 5120 1770 5160 1780
rect 5240 1770 5320 1780
rect 5400 1770 5480 1780
rect 6360 1770 6400 1780
rect 6840 1770 7040 1780
rect 7120 1770 7360 1780
rect 7840 1770 7920 1780
rect 8480 1770 8600 1780
rect 8920 1770 9120 1780
rect 9200 1770 9240 1780
rect 9680 1770 9720 1780
rect 9760 1770 9800 1780
rect 1880 1760 2040 1770
rect 2200 1760 2240 1770
rect 2360 1760 2440 1770
rect 2520 1760 2760 1770
rect 3160 1760 3240 1770
rect 4200 1760 4240 1770
rect 4480 1760 4520 1770
rect 4720 1760 4760 1770
rect 4840 1760 4880 1770
rect 4960 1760 5080 1770
rect 5120 1760 5160 1770
rect 5240 1760 5320 1770
rect 5400 1760 5480 1770
rect 6360 1760 6400 1770
rect 6840 1760 7040 1770
rect 7120 1760 7360 1770
rect 7840 1760 7920 1770
rect 8480 1760 8600 1770
rect 8920 1760 9120 1770
rect 9200 1760 9240 1770
rect 9680 1760 9720 1770
rect 9760 1760 9800 1770
rect 1880 1750 2040 1760
rect 2200 1750 2240 1760
rect 2360 1750 2440 1760
rect 2520 1750 2760 1760
rect 3160 1750 3240 1760
rect 4200 1750 4240 1760
rect 4480 1750 4520 1760
rect 4720 1750 4760 1760
rect 4840 1750 4880 1760
rect 4960 1750 5080 1760
rect 5120 1750 5160 1760
rect 5240 1750 5320 1760
rect 5400 1750 5480 1760
rect 6360 1750 6400 1760
rect 6840 1750 7040 1760
rect 7120 1750 7360 1760
rect 7840 1750 7920 1760
rect 8480 1750 8600 1760
rect 8920 1750 9120 1760
rect 9200 1750 9240 1760
rect 9680 1750 9720 1760
rect 9760 1750 9800 1760
rect 1880 1740 2040 1750
rect 2200 1740 2240 1750
rect 2360 1740 2440 1750
rect 2520 1740 2760 1750
rect 3160 1740 3240 1750
rect 4200 1740 4240 1750
rect 4480 1740 4520 1750
rect 4720 1740 4760 1750
rect 4840 1740 4880 1750
rect 4960 1740 5080 1750
rect 5120 1740 5160 1750
rect 5240 1740 5320 1750
rect 5400 1740 5480 1750
rect 6360 1740 6400 1750
rect 6840 1740 7040 1750
rect 7120 1740 7360 1750
rect 7840 1740 7920 1750
rect 8480 1740 8600 1750
rect 8920 1740 9120 1750
rect 9200 1740 9240 1750
rect 9680 1740 9720 1750
rect 9760 1740 9800 1750
rect 1920 1730 2040 1740
rect 2440 1730 2680 1740
rect 3160 1730 3240 1740
rect 4160 1730 4240 1740
rect 4480 1730 4520 1740
rect 4760 1730 4800 1740
rect 4840 1730 4880 1740
rect 4960 1730 5000 1740
rect 5120 1730 5160 1740
rect 5240 1730 5320 1740
rect 5360 1730 5400 1740
rect 5480 1730 5560 1740
rect 6840 1730 7000 1740
rect 7120 1730 7360 1740
rect 7840 1730 7960 1740
rect 8320 1730 8360 1740
rect 8520 1730 8600 1740
rect 8880 1730 9120 1740
rect 9200 1730 9240 1740
rect 9680 1730 9720 1740
rect 9760 1730 9800 1740
rect 9880 1730 9960 1740
rect 1920 1720 2040 1730
rect 2440 1720 2680 1730
rect 3160 1720 3240 1730
rect 4160 1720 4240 1730
rect 4480 1720 4520 1730
rect 4760 1720 4800 1730
rect 4840 1720 4880 1730
rect 4960 1720 5000 1730
rect 5120 1720 5160 1730
rect 5240 1720 5320 1730
rect 5360 1720 5400 1730
rect 5480 1720 5560 1730
rect 6840 1720 7000 1730
rect 7120 1720 7360 1730
rect 7840 1720 7960 1730
rect 8320 1720 8360 1730
rect 8520 1720 8600 1730
rect 8880 1720 9120 1730
rect 9200 1720 9240 1730
rect 9680 1720 9720 1730
rect 9760 1720 9800 1730
rect 9880 1720 9960 1730
rect 1920 1710 2040 1720
rect 2440 1710 2680 1720
rect 3160 1710 3240 1720
rect 4160 1710 4240 1720
rect 4480 1710 4520 1720
rect 4760 1710 4800 1720
rect 4840 1710 4880 1720
rect 4960 1710 5000 1720
rect 5120 1710 5160 1720
rect 5240 1710 5320 1720
rect 5360 1710 5400 1720
rect 5480 1710 5560 1720
rect 6840 1710 7000 1720
rect 7120 1710 7360 1720
rect 7840 1710 7960 1720
rect 8320 1710 8360 1720
rect 8520 1710 8600 1720
rect 8880 1710 9120 1720
rect 9200 1710 9240 1720
rect 9680 1710 9720 1720
rect 9760 1710 9800 1720
rect 9880 1710 9960 1720
rect 1920 1700 2040 1710
rect 2440 1700 2680 1710
rect 3160 1700 3240 1710
rect 4160 1700 4240 1710
rect 4480 1700 4520 1710
rect 4760 1700 4800 1710
rect 4840 1700 4880 1710
rect 4960 1700 5000 1710
rect 5120 1700 5160 1710
rect 5240 1700 5320 1710
rect 5360 1700 5400 1710
rect 5480 1700 5560 1710
rect 6840 1700 7000 1710
rect 7120 1700 7360 1710
rect 7840 1700 7960 1710
rect 8320 1700 8360 1710
rect 8520 1700 8600 1710
rect 8880 1700 9120 1710
rect 9200 1700 9240 1710
rect 9680 1700 9720 1710
rect 9760 1700 9800 1710
rect 9880 1700 9960 1710
rect 1920 1690 2040 1700
rect 2480 1690 2680 1700
rect 3120 1690 3200 1700
rect 4080 1690 4240 1700
rect 4840 1690 4880 1700
rect 4960 1690 5000 1700
rect 5080 1690 5120 1700
rect 5200 1690 5280 1700
rect 5320 1690 5480 1700
rect 5520 1690 5560 1700
rect 6840 1690 7000 1700
rect 7120 1690 7360 1700
rect 7880 1690 7960 1700
rect 8320 1690 8360 1700
rect 8520 1690 8600 1700
rect 8840 1690 9080 1700
rect 9200 1690 9240 1700
rect 9720 1690 9800 1700
rect 1920 1680 2040 1690
rect 2480 1680 2680 1690
rect 3120 1680 3200 1690
rect 4080 1680 4240 1690
rect 4840 1680 4880 1690
rect 4960 1680 5000 1690
rect 5080 1680 5120 1690
rect 5200 1680 5280 1690
rect 5320 1680 5480 1690
rect 5520 1680 5560 1690
rect 6840 1680 7000 1690
rect 7120 1680 7360 1690
rect 7880 1680 7960 1690
rect 8320 1680 8360 1690
rect 8520 1680 8600 1690
rect 8840 1680 9080 1690
rect 9200 1680 9240 1690
rect 9720 1680 9800 1690
rect 1920 1670 2040 1680
rect 2480 1670 2680 1680
rect 3120 1670 3200 1680
rect 4080 1670 4240 1680
rect 4840 1670 4880 1680
rect 4960 1670 5000 1680
rect 5080 1670 5120 1680
rect 5200 1670 5280 1680
rect 5320 1670 5480 1680
rect 5520 1670 5560 1680
rect 6840 1670 7000 1680
rect 7120 1670 7360 1680
rect 7880 1670 7960 1680
rect 8320 1670 8360 1680
rect 8520 1670 8600 1680
rect 8840 1670 9080 1680
rect 9200 1670 9240 1680
rect 9720 1670 9800 1680
rect 1920 1660 2040 1670
rect 2480 1660 2680 1670
rect 3120 1660 3200 1670
rect 4080 1660 4240 1670
rect 4840 1660 4880 1670
rect 4960 1660 5000 1670
rect 5080 1660 5120 1670
rect 5200 1660 5280 1670
rect 5320 1660 5480 1670
rect 5520 1660 5560 1670
rect 6840 1660 7000 1670
rect 7120 1660 7360 1670
rect 7880 1660 7960 1670
rect 8320 1660 8360 1670
rect 8520 1660 8600 1670
rect 8840 1660 9080 1670
rect 9200 1660 9240 1670
rect 9720 1660 9800 1670
rect 1920 1650 2080 1660
rect 2400 1650 2760 1660
rect 3080 1650 3200 1660
rect 4200 1650 4280 1660
rect 4480 1650 4520 1660
rect 4960 1650 5000 1660
rect 5080 1650 5120 1660
rect 5200 1650 5360 1660
rect 5400 1650 5560 1660
rect 6840 1650 7000 1660
rect 7160 1650 7360 1660
rect 7880 1650 7960 1660
rect 8480 1650 8640 1660
rect 8840 1650 9080 1660
rect 9200 1650 9240 1660
rect 9840 1650 9880 1660
rect 1920 1640 2080 1650
rect 2400 1640 2760 1650
rect 3080 1640 3200 1650
rect 4200 1640 4280 1650
rect 4480 1640 4520 1650
rect 4960 1640 5000 1650
rect 5080 1640 5120 1650
rect 5200 1640 5360 1650
rect 5400 1640 5560 1650
rect 6840 1640 7000 1650
rect 7160 1640 7360 1650
rect 7880 1640 7960 1650
rect 8480 1640 8640 1650
rect 8840 1640 9080 1650
rect 9200 1640 9240 1650
rect 9840 1640 9880 1650
rect 1920 1630 2080 1640
rect 2400 1630 2760 1640
rect 3080 1630 3200 1640
rect 4200 1630 4280 1640
rect 4480 1630 4520 1640
rect 4960 1630 5000 1640
rect 5080 1630 5120 1640
rect 5200 1630 5360 1640
rect 5400 1630 5560 1640
rect 6840 1630 7000 1640
rect 7160 1630 7360 1640
rect 7880 1630 7960 1640
rect 8480 1630 8640 1640
rect 8840 1630 9080 1640
rect 9200 1630 9240 1640
rect 9840 1630 9880 1640
rect 1920 1620 2080 1630
rect 2400 1620 2760 1630
rect 3080 1620 3200 1630
rect 4200 1620 4280 1630
rect 4480 1620 4520 1630
rect 4960 1620 5000 1630
rect 5080 1620 5120 1630
rect 5200 1620 5360 1630
rect 5400 1620 5560 1630
rect 6840 1620 7000 1630
rect 7160 1620 7360 1630
rect 7880 1620 7960 1630
rect 8480 1620 8640 1630
rect 8840 1620 9080 1630
rect 9200 1620 9240 1630
rect 9840 1620 9880 1630
rect 1960 1610 2080 1620
rect 2360 1610 2720 1620
rect 3040 1610 3160 1620
rect 4200 1610 4280 1620
rect 5160 1610 5240 1620
rect 5280 1610 5320 1620
rect 5360 1610 5520 1620
rect 5560 1610 5680 1620
rect 6840 1610 7000 1620
rect 7120 1610 7360 1620
rect 7880 1610 7960 1620
rect 8440 1610 8640 1620
rect 8680 1610 8720 1620
rect 8760 1610 9080 1620
rect 9120 1610 9200 1620
rect 1960 1600 2080 1610
rect 2360 1600 2720 1610
rect 3040 1600 3160 1610
rect 4200 1600 4280 1610
rect 5160 1600 5240 1610
rect 5280 1600 5320 1610
rect 5360 1600 5520 1610
rect 5560 1600 5680 1610
rect 6840 1600 7000 1610
rect 7120 1600 7360 1610
rect 7880 1600 7960 1610
rect 8440 1600 8640 1610
rect 8680 1600 8720 1610
rect 8760 1600 9080 1610
rect 9120 1600 9200 1610
rect 1960 1590 2080 1600
rect 2360 1590 2720 1600
rect 3040 1590 3160 1600
rect 4200 1590 4280 1600
rect 5160 1590 5240 1600
rect 5280 1590 5320 1600
rect 5360 1590 5520 1600
rect 5560 1590 5680 1600
rect 6840 1590 7000 1600
rect 7120 1590 7360 1600
rect 7880 1590 7960 1600
rect 8440 1590 8640 1600
rect 8680 1590 8720 1600
rect 8760 1590 9080 1600
rect 9120 1590 9200 1600
rect 1960 1580 2080 1590
rect 2360 1580 2720 1590
rect 3040 1580 3160 1590
rect 4200 1580 4280 1590
rect 5160 1580 5240 1590
rect 5280 1580 5320 1590
rect 5360 1580 5520 1590
rect 5560 1580 5680 1590
rect 6840 1580 7000 1590
rect 7120 1580 7360 1590
rect 7880 1580 7960 1590
rect 8440 1580 8640 1590
rect 8680 1580 8720 1590
rect 8760 1580 9080 1590
rect 9120 1580 9200 1590
rect 2000 1570 2120 1580
rect 2440 1570 2520 1580
rect 2960 1570 3120 1580
rect 4240 1570 4280 1580
rect 5240 1570 5320 1580
rect 5560 1570 5600 1580
rect 5640 1570 5720 1580
rect 6840 1570 7000 1580
rect 7160 1570 7360 1580
rect 7880 1570 8000 1580
rect 8280 1570 8320 1580
rect 8440 1570 8600 1580
rect 8680 1570 9080 1580
rect 9720 1570 9760 1580
rect 9840 1570 9960 1580
rect 2000 1560 2120 1570
rect 2440 1560 2520 1570
rect 2960 1560 3120 1570
rect 4240 1560 4280 1570
rect 5240 1560 5320 1570
rect 5560 1560 5600 1570
rect 5640 1560 5720 1570
rect 6840 1560 7000 1570
rect 7160 1560 7360 1570
rect 7880 1560 8000 1570
rect 8280 1560 8320 1570
rect 8440 1560 8600 1570
rect 8680 1560 9080 1570
rect 9720 1560 9760 1570
rect 9840 1560 9960 1570
rect 2000 1550 2120 1560
rect 2440 1550 2520 1560
rect 2960 1550 3120 1560
rect 4240 1550 4280 1560
rect 5240 1550 5320 1560
rect 5560 1550 5600 1560
rect 5640 1550 5720 1560
rect 6840 1550 7000 1560
rect 7160 1550 7360 1560
rect 7880 1550 8000 1560
rect 8280 1550 8320 1560
rect 8440 1550 8600 1560
rect 8680 1550 9080 1560
rect 9720 1550 9760 1560
rect 9840 1550 9960 1560
rect 2000 1540 2120 1550
rect 2440 1540 2520 1550
rect 2960 1540 3120 1550
rect 4240 1540 4280 1550
rect 5240 1540 5320 1550
rect 5560 1540 5600 1550
rect 5640 1540 5720 1550
rect 6840 1540 7000 1550
rect 7160 1540 7360 1550
rect 7880 1540 8000 1550
rect 8280 1540 8320 1550
rect 8440 1540 8600 1550
rect 8680 1540 9080 1550
rect 9720 1540 9760 1550
rect 9840 1540 9960 1550
rect 2000 1530 2200 1540
rect 2920 1530 3080 1540
rect 4320 1530 4360 1540
rect 5280 1530 5320 1540
rect 5560 1530 5640 1540
rect 5680 1530 5720 1540
rect 6840 1530 7000 1540
rect 7200 1530 7360 1540
rect 7880 1530 8000 1540
rect 8280 1530 8320 1540
rect 8440 1530 8640 1540
rect 8680 1530 9080 1540
rect 9880 1530 9990 1540
rect 2000 1520 2200 1530
rect 2920 1520 3080 1530
rect 4320 1520 4360 1530
rect 5280 1520 5320 1530
rect 5560 1520 5640 1530
rect 5680 1520 5720 1530
rect 6840 1520 7000 1530
rect 7200 1520 7360 1530
rect 7880 1520 8000 1530
rect 8280 1520 8320 1530
rect 8440 1520 8640 1530
rect 8680 1520 9080 1530
rect 9880 1520 9990 1530
rect 2000 1510 2200 1520
rect 2920 1510 3080 1520
rect 4320 1510 4360 1520
rect 5280 1510 5320 1520
rect 5560 1510 5640 1520
rect 5680 1510 5720 1520
rect 6840 1510 7000 1520
rect 7200 1510 7360 1520
rect 7880 1510 8000 1520
rect 8280 1510 8320 1520
rect 8440 1510 8640 1520
rect 8680 1510 9080 1520
rect 9880 1510 9990 1520
rect 2000 1500 2200 1510
rect 2920 1500 3080 1510
rect 4320 1500 4360 1510
rect 5280 1500 5320 1510
rect 5560 1500 5640 1510
rect 5680 1500 5720 1510
rect 6840 1500 7000 1510
rect 7200 1500 7360 1510
rect 7880 1500 8000 1510
rect 8280 1500 8320 1510
rect 8440 1500 8640 1510
rect 8680 1500 9080 1510
rect 9880 1500 9990 1510
rect 2040 1490 2200 1500
rect 2880 1490 2960 1500
rect 3000 1490 3040 1500
rect 4160 1490 4240 1500
rect 5440 1490 5520 1500
rect 5560 1490 5640 1500
rect 5680 1490 5720 1500
rect 6800 1490 6960 1500
rect 7240 1490 7360 1500
rect 7880 1490 8000 1500
rect 8440 1490 8600 1500
rect 8720 1490 9080 1500
rect 9120 1490 9200 1500
rect 9680 1490 9720 1500
rect 9880 1490 9920 1500
rect 2040 1480 2200 1490
rect 2880 1480 2960 1490
rect 3000 1480 3040 1490
rect 4160 1480 4240 1490
rect 5440 1480 5520 1490
rect 5560 1480 5640 1490
rect 5680 1480 5720 1490
rect 6800 1480 6960 1490
rect 7240 1480 7360 1490
rect 7880 1480 8000 1490
rect 8440 1480 8600 1490
rect 8720 1480 9080 1490
rect 9120 1480 9200 1490
rect 9680 1480 9720 1490
rect 9880 1480 9920 1490
rect 2040 1470 2200 1480
rect 2880 1470 2960 1480
rect 3000 1470 3040 1480
rect 4160 1470 4240 1480
rect 5440 1470 5520 1480
rect 5560 1470 5640 1480
rect 5680 1470 5720 1480
rect 6800 1470 6960 1480
rect 7240 1470 7360 1480
rect 7880 1470 8000 1480
rect 8440 1470 8600 1480
rect 8720 1470 9080 1480
rect 9120 1470 9200 1480
rect 9680 1470 9720 1480
rect 9880 1470 9920 1480
rect 2040 1460 2200 1470
rect 2880 1460 2960 1470
rect 3000 1460 3040 1470
rect 4160 1460 4240 1470
rect 5440 1460 5520 1470
rect 5560 1460 5640 1470
rect 5680 1460 5720 1470
rect 6800 1460 6960 1470
rect 7240 1460 7360 1470
rect 7880 1460 8000 1470
rect 8440 1460 8600 1470
rect 8720 1460 9080 1470
rect 9120 1460 9200 1470
rect 9680 1460 9720 1470
rect 9880 1460 9920 1470
rect 2080 1450 2240 1460
rect 2840 1450 2920 1460
rect 4160 1450 4280 1460
rect 5440 1450 5560 1460
rect 5600 1450 5640 1460
rect 6800 1450 6880 1460
rect 7240 1450 7360 1460
rect 7880 1450 8000 1460
rect 8240 1450 8280 1460
rect 8440 1450 8600 1460
rect 8680 1450 9120 1460
rect 9560 1450 9720 1460
rect 9760 1450 9800 1460
rect 2080 1440 2240 1450
rect 2840 1440 2920 1450
rect 4160 1440 4280 1450
rect 5440 1440 5560 1450
rect 5600 1440 5640 1450
rect 6800 1440 6880 1450
rect 7240 1440 7360 1450
rect 7880 1440 8000 1450
rect 8240 1440 8280 1450
rect 8440 1440 8600 1450
rect 8680 1440 9120 1450
rect 9560 1440 9720 1450
rect 9760 1440 9800 1450
rect 2080 1430 2240 1440
rect 2840 1430 2920 1440
rect 4160 1430 4280 1440
rect 5440 1430 5560 1440
rect 5600 1430 5640 1440
rect 6800 1430 6880 1440
rect 7240 1430 7360 1440
rect 7880 1430 8000 1440
rect 8240 1430 8280 1440
rect 8440 1430 8600 1440
rect 8680 1430 9120 1440
rect 9560 1430 9720 1440
rect 9760 1430 9800 1440
rect 2080 1420 2240 1430
rect 2840 1420 2920 1430
rect 4160 1420 4280 1430
rect 5440 1420 5560 1430
rect 5600 1420 5640 1430
rect 6800 1420 6880 1430
rect 7240 1420 7360 1430
rect 7880 1420 8000 1430
rect 8240 1420 8280 1430
rect 8440 1420 8600 1430
rect 8680 1420 9120 1430
rect 9560 1420 9720 1430
rect 9760 1420 9800 1430
rect 2120 1410 2280 1420
rect 2800 1410 2880 1420
rect 4160 1410 4320 1420
rect 4360 1410 4400 1420
rect 5440 1410 5520 1420
rect 5560 1410 5600 1420
rect 6800 1410 6840 1420
rect 7280 1410 7360 1420
rect 7920 1410 8000 1420
rect 8200 1410 8280 1420
rect 8440 1410 9120 1420
rect 9200 1410 9280 1420
rect 9600 1410 9680 1420
rect 9920 1410 9990 1420
rect 2120 1400 2280 1410
rect 2800 1400 2880 1410
rect 4160 1400 4320 1410
rect 4360 1400 4400 1410
rect 5440 1400 5520 1410
rect 5560 1400 5600 1410
rect 6800 1400 6840 1410
rect 7280 1400 7360 1410
rect 7920 1400 8000 1410
rect 8200 1400 8280 1410
rect 8440 1400 9120 1410
rect 9200 1400 9280 1410
rect 9600 1400 9680 1410
rect 9920 1400 9990 1410
rect 2120 1390 2280 1400
rect 2800 1390 2880 1400
rect 4160 1390 4320 1400
rect 4360 1390 4400 1400
rect 5440 1390 5520 1400
rect 5560 1390 5600 1400
rect 6800 1390 6840 1400
rect 7280 1390 7360 1400
rect 7920 1390 8000 1400
rect 8200 1390 8280 1400
rect 8440 1390 9120 1400
rect 9200 1390 9280 1400
rect 9600 1390 9680 1400
rect 9920 1390 9990 1400
rect 2120 1380 2280 1390
rect 2800 1380 2880 1390
rect 4160 1380 4320 1390
rect 4360 1380 4400 1390
rect 5440 1380 5520 1390
rect 5560 1380 5600 1390
rect 6800 1380 6840 1390
rect 7280 1380 7360 1390
rect 7920 1380 8000 1390
rect 8200 1380 8280 1390
rect 8440 1380 9120 1390
rect 9200 1380 9280 1390
rect 9600 1380 9680 1390
rect 9920 1380 9990 1390
rect 2200 1370 2360 1380
rect 2760 1370 2840 1380
rect 3560 1370 3600 1380
rect 4240 1370 4320 1380
rect 5520 1370 5600 1380
rect 7280 1370 7400 1380
rect 7920 1370 8000 1380
rect 8160 1370 8240 1380
rect 8440 1370 9120 1380
rect 9160 1370 9280 1380
rect 9640 1370 9680 1380
rect 9720 1370 9760 1380
rect 9800 1370 9840 1380
rect 9960 1370 9990 1380
rect 2200 1360 2360 1370
rect 2760 1360 2840 1370
rect 3560 1360 3600 1370
rect 4240 1360 4320 1370
rect 5520 1360 5600 1370
rect 7280 1360 7400 1370
rect 7920 1360 8000 1370
rect 8160 1360 8240 1370
rect 8440 1360 9120 1370
rect 9160 1360 9280 1370
rect 9640 1360 9680 1370
rect 9720 1360 9760 1370
rect 9800 1360 9840 1370
rect 9960 1360 9990 1370
rect 2200 1350 2360 1360
rect 2760 1350 2840 1360
rect 3560 1350 3600 1360
rect 4240 1350 4320 1360
rect 5520 1350 5600 1360
rect 7280 1350 7400 1360
rect 7920 1350 8000 1360
rect 8160 1350 8240 1360
rect 8440 1350 9120 1360
rect 9160 1350 9280 1360
rect 9640 1350 9680 1360
rect 9720 1350 9760 1360
rect 9800 1350 9840 1360
rect 9960 1350 9990 1360
rect 2200 1340 2360 1350
rect 2760 1340 2840 1350
rect 3560 1340 3600 1350
rect 4240 1340 4320 1350
rect 5520 1340 5600 1350
rect 7280 1340 7400 1350
rect 7920 1340 8000 1350
rect 8160 1340 8240 1350
rect 8440 1340 9120 1350
rect 9160 1340 9280 1350
rect 9640 1340 9680 1350
rect 9720 1340 9760 1350
rect 9800 1340 9840 1350
rect 9960 1340 9990 1350
rect 2240 1330 2440 1340
rect 2680 1330 2760 1340
rect 3640 1330 3680 1340
rect 4200 1330 4280 1340
rect 7320 1330 7400 1340
rect 7920 1330 8200 1340
rect 8440 1330 9160 1340
rect 9240 1330 9280 1340
rect 9640 1330 9680 1340
rect 9760 1330 9800 1340
rect 9960 1330 9990 1340
rect 2240 1320 2440 1330
rect 2680 1320 2760 1330
rect 3640 1320 3680 1330
rect 4200 1320 4280 1330
rect 7320 1320 7400 1330
rect 7920 1320 8200 1330
rect 8440 1320 9160 1330
rect 9240 1320 9280 1330
rect 9640 1320 9680 1330
rect 9760 1320 9800 1330
rect 9960 1320 9990 1330
rect 2240 1310 2440 1320
rect 2680 1310 2760 1320
rect 3640 1310 3680 1320
rect 4200 1310 4280 1320
rect 7320 1310 7400 1320
rect 7920 1310 8200 1320
rect 8440 1310 9160 1320
rect 9240 1310 9280 1320
rect 9640 1310 9680 1320
rect 9760 1310 9800 1320
rect 9960 1310 9990 1320
rect 2240 1300 2440 1310
rect 2680 1300 2760 1310
rect 3640 1300 3680 1310
rect 4200 1300 4280 1310
rect 7320 1300 7400 1310
rect 7920 1300 8200 1310
rect 8440 1300 9160 1310
rect 9240 1300 9280 1310
rect 9640 1300 9680 1310
rect 9760 1300 9800 1310
rect 9960 1300 9990 1310
rect 2440 1290 2680 1300
rect 4200 1290 4240 1300
rect 4400 1290 4440 1300
rect 7280 1290 7400 1300
rect 7920 1290 8160 1300
rect 8440 1290 9080 1300
rect 9120 1290 9160 1300
rect 9280 1290 9320 1300
rect 9640 1290 9760 1300
rect 9960 1290 9990 1300
rect 2440 1280 2680 1290
rect 4200 1280 4240 1290
rect 4400 1280 4440 1290
rect 7280 1280 7400 1290
rect 7920 1280 8160 1290
rect 8440 1280 9080 1290
rect 9120 1280 9160 1290
rect 9280 1280 9320 1290
rect 9640 1280 9760 1290
rect 9960 1280 9990 1290
rect 2440 1270 2680 1280
rect 4200 1270 4240 1280
rect 4400 1270 4440 1280
rect 7280 1270 7400 1280
rect 7920 1270 8160 1280
rect 8440 1270 9080 1280
rect 9120 1270 9160 1280
rect 9280 1270 9320 1280
rect 9640 1270 9760 1280
rect 9960 1270 9990 1280
rect 2440 1260 2680 1270
rect 4200 1260 4240 1270
rect 4400 1260 4440 1270
rect 7280 1260 7400 1270
rect 7920 1260 8160 1270
rect 8440 1260 9080 1270
rect 9120 1260 9160 1270
rect 9280 1260 9320 1270
rect 9640 1260 9760 1270
rect 9960 1260 9990 1270
rect 3520 1250 3680 1260
rect 5200 1250 5440 1260
rect 7320 1250 7400 1260
rect 7960 1250 8200 1260
rect 8440 1250 8960 1260
rect 9000 1250 9080 1260
rect 9120 1250 9160 1260
rect 9280 1250 9320 1260
rect 9600 1250 9640 1260
rect 9720 1250 9760 1260
rect 9800 1250 9840 1260
rect 9920 1250 9960 1260
rect 3520 1240 3680 1250
rect 5200 1240 5440 1250
rect 7320 1240 7400 1250
rect 7960 1240 8200 1250
rect 8440 1240 8960 1250
rect 9000 1240 9080 1250
rect 9120 1240 9160 1250
rect 9280 1240 9320 1250
rect 9600 1240 9640 1250
rect 9720 1240 9760 1250
rect 9800 1240 9840 1250
rect 9920 1240 9960 1250
rect 3520 1230 3680 1240
rect 5200 1230 5440 1240
rect 7320 1230 7400 1240
rect 7960 1230 8200 1240
rect 8440 1230 8960 1240
rect 9000 1230 9080 1240
rect 9120 1230 9160 1240
rect 9280 1230 9320 1240
rect 9600 1230 9640 1240
rect 9720 1230 9760 1240
rect 9800 1230 9840 1240
rect 9920 1230 9960 1240
rect 3520 1220 3680 1230
rect 5200 1220 5440 1230
rect 7320 1220 7400 1230
rect 7960 1220 8200 1230
rect 8440 1220 8960 1230
rect 9000 1220 9080 1230
rect 9120 1220 9160 1230
rect 9280 1220 9320 1230
rect 9600 1220 9640 1230
rect 9720 1220 9760 1230
rect 9800 1220 9840 1230
rect 9920 1220 9960 1230
rect 3680 1210 3720 1220
rect 3800 1210 3840 1220
rect 4200 1210 4240 1220
rect 5000 1210 5080 1220
rect 5120 1210 5160 1220
rect 5200 1210 5240 1220
rect 5320 1210 5360 1220
rect 6720 1210 6800 1220
rect 7320 1210 7400 1220
rect 7960 1210 8200 1220
rect 8400 1210 8840 1220
rect 9000 1210 9040 1220
rect 9120 1210 9160 1220
rect 9280 1210 9360 1220
rect 9520 1210 9560 1220
rect 9640 1210 9720 1220
rect 9800 1210 9840 1220
rect 9920 1210 9990 1220
rect 3680 1200 3720 1210
rect 3800 1200 3840 1210
rect 4200 1200 4240 1210
rect 5000 1200 5080 1210
rect 5120 1200 5160 1210
rect 5200 1200 5240 1210
rect 5320 1200 5360 1210
rect 6720 1200 6800 1210
rect 7320 1200 7400 1210
rect 7960 1200 8200 1210
rect 8400 1200 8840 1210
rect 9000 1200 9040 1210
rect 9120 1200 9160 1210
rect 9280 1200 9360 1210
rect 9520 1200 9560 1210
rect 9640 1200 9720 1210
rect 9800 1200 9840 1210
rect 9920 1200 9990 1210
rect 3680 1190 3720 1200
rect 3800 1190 3840 1200
rect 4200 1190 4240 1200
rect 5000 1190 5080 1200
rect 5120 1190 5160 1200
rect 5200 1190 5240 1200
rect 5320 1190 5360 1200
rect 6720 1190 6800 1200
rect 7320 1190 7400 1200
rect 7960 1190 8200 1200
rect 8400 1190 8840 1200
rect 9000 1190 9040 1200
rect 9120 1190 9160 1200
rect 9280 1190 9360 1200
rect 9520 1190 9560 1200
rect 9640 1190 9720 1200
rect 9800 1190 9840 1200
rect 9920 1190 9990 1200
rect 3680 1180 3720 1190
rect 3800 1180 3840 1190
rect 4200 1180 4240 1190
rect 5000 1180 5080 1190
rect 5120 1180 5160 1190
rect 5200 1180 5240 1190
rect 5320 1180 5360 1190
rect 6720 1180 6800 1190
rect 7320 1180 7400 1190
rect 7960 1180 8200 1190
rect 8400 1180 8840 1190
rect 9000 1180 9040 1190
rect 9120 1180 9160 1190
rect 9280 1180 9360 1190
rect 9520 1180 9560 1190
rect 9640 1180 9720 1190
rect 9800 1180 9840 1190
rect 9920 1180 9990 1190
rect 800 1170 840 1180
rect 3720 1170 3760 1180
rect 4200 1170 4240 1180
rect 4440 1170 4480 1180
rect 4760 1170 4840 1180
rect 6680 1170 6720 1180
rect 6760 1170 6800 1180
rect 7320 1170 7400 1180
rect 7960 1170 8160 1180
rect 8360 1170 8720 1180
rect 9120 1170 9160 1180
rect 9280 1170 9400 1180
rect 9520 1170 9560 1180
rect 9680 1170 9720 1180
rect 9800 1170 9840 1180
rect 800 1160 840 1170
rect 3720 1160 3760 1170
rect 4200 1160 4240 1170
rect 4440 1160 4480 1170
rect 4760 1160 4840 1170
rect 6680 1160 6720 1170
rect 6760 1160 6800 1170
rect 7320 1160 7400 1170
rect 7960 1160 8160 1170
rect 8360 1160 8720 1170
rect 9120 1160 9160 1170
rect 9280 1160 9400 1170
rect 9520 1160 9560 1170
rect 9680 1160 9720 1170
rect 9800 1160 9840 1170
rect 800 1150 840 1160
rect 3720 1150 3760 1160
rect 4200 1150 4240 1160
rect 4440 1150 4480 1160
rect 4760 1150 4840 1160
rect 6680 1150 6720 1160
rect 6760 1150 6800 1160
rect 7320 1150 7400 1160
rect 7960 1150 8160 1160
rect 8360 1150 8720 1160
rect 9120 1150 9160 1160
rect 9280 1150 9400 1160
rect 9520 1150 9560 1160
rect 9680 1150 9720 1160
rect 9800 1150 9840 1160
rect 800 1140 840 1150
rect 3720 1140 3760 1150
rect 4200 1140 4240 1150
rect 4440 1140 4480 1150
rect 4760 1140 4840 1150
rect 6680 1140 6720 1150
rect 6760 1140 6800 1150
rect 7320 1140 7400 1150
rect 7960 1140 8160 1150
rect 8360 1140 8720 1150
rect 9120 1140 9160 1150
rect 9280 1140 9400 1150
rect 9520 1140 9560 1150
rect 9680 1140 9720 1150
rect 9800 1140 9840 1150
rect 760 1130 840 1140
rect 3720 1130 3760 1140
rect 3920 1130 3960 1140
rect 4440 1130 4480 1140
rect 6600 1130 6640 1140
rect 6760 1130 6800 1140
rect 7320 1130 7400 1140
rect 7960 1130 8160 1140
rect 8360 1130 8680 1140
rect 9120 1130 9160 1140
rect 9280 1130 9400 1140
rect 9520 1130 9560 1140
rect 9600 1130 9640 1140
rect 9840 1130 9960 1140
rect 760 1120 840 1130
rect 3720 1120 3760 1130
rect 3920 1120 3960 1130
rect 4440 1120 4480 1130
rect 6600 1120 6640 1130
rect 6760 1120 6800 1130
rect 7320 1120 7400 1130
rect 7960 1120 8160 1130
rect 8360 1120 8680 1130
rect 9120 1120 9160 1130
rect 9280 1120 9400 1130
rect 9520 1120 9560 1130
rect 9600 1120 9640 1130
rect 9840 1120 9960 1130
rect 760 1110 840 1120
rect 3720 1110 3760 1120
rect 3920 1110 3960 1120
rect 4440 1110 4480 1120
rect 6600 1110 6640 1120
rect 6760 1110 6800 1120
rect 7320 1110 7400 1120
rect 7960 1110 8160 1120
rect 8360 1110 8680 1120
rect 9120 1110 9160 1120
rect 9280 1110 9400 1120
rect 9520 1110 9560 1120
rect 9600 1110 9640 1120
rect 9840 1110 9960 1120
rect 760 1100 840 1110
rect 3720 1100 3760 1110
rect 3920 1100 3960 1110
rect 4440 1100 4480 1110
rect 6600 1100 6640 1110
rect 6760 1100 6800 1110
rect 7320 1100 7400 1110
rect 7960 1100 8160 1110
rect 8360 1100 8680 1110
rect 9120 1100 9160 1110
rect 9280 1100 9400 1110
rect 9520 1100 9560 1110
rect 9600 1100 9640 1110
rect 9840 1100 9960 1110
rect 760 1090 840 1100
rect 1520 1090 1640 1100
rect 3680 1090 3840 1100
rect 3960 1090 4000 1100
rect 6520 1090 6560 1100
rect 7320 1090 7400 1100
rect 7960 1090 8160 1100
rect 8360 1090 8680 1100
rect 9120 1090 9440 1100
rect 9520 1090 9600 1100
rect 9840 1090 9990 1100
rect 760 1080 840 1090
rect 1520 1080 1640 1090
rect 3680 1080 3840 1090
rect 3960 1080 4000 1090
rect 6520 1080 6560 1090
rect 7320 1080 7400 1090
rect 7960 1080 8160 1090
rect 8360 1080 8680 1090
rect 9120 1080 9440 1090
rect 9520 1080 9600 1090
rect 9840 1080 9990 1090
rect 760 1070 840 1080
rect 1520 1070 1640 1080
rect 3680 1070 3840 1080
rect 3960 1070 4000 1080
rect 6520 1070 6560 1080
rect 7320 1070 7400 1080
rect 7960 1070 8160 1080
rect 8360 1070 8680 1080
rect 9120 1070 9440 1080
rect 9520 1070 9600 1080
rect 9840 1070 9990 1080
rect 760 1060 840 1070
rect 1520 1060 1640 1070
rect 3680 1060 3840 1070
rect 3960 1060 4000 1070
rect 6520 1060 6560 1070
rect 7320 1060 7400 1070
rect 7960 1060 8160 1070
rect 8360 1060 8680 1070
rect 9120 1060 9440 1070
rect 9520 1060 9600 1070
rect 9840 1060 9990 1070
rect 760 1050 800 1060
rect 1480 1050 1520 1060
rect 2080 1050 2200 1060
rect 3720 1050 3760 1060
rect 3840 1050 3880 1060
rect 4040 1050 4080 1060
rect 4200 1050 4240 1060
rect 4520 1050 4600 1060
rect 6480 1050 6560 1060
rect 6840 1050 6880 1060
rect 7320 1050 7400 1060
rect 7960 1050 8160 1060
rect 8360 1050 8560 1060
rect 9120 1050 9160 1060
rect 9240 1050 9320 1060
rect 9360 1050 9440 1060
rect 9720 1050 9760 1060
rect 9840 1050 9990 1060
rect 760 1040 800 1050
rect 1480 1040 1520 1050
rect 2080 1040 2200 1050
rect 3720 1040 3760 1050
rect 3840 1040 3880 1050
rect 4040 1040 4080 1050
rect 4200 1040 4240 1050
rect 4520 1040 4600 1050
rect 6480 1040 6560 1050
rect 6840 1040 6880 1050
rect 7320 1040 7400 1050
rect 7960 1040 8160 1050
rect 8360 1040 8560 1050
rect 9120 1040 9160 1050
rect 9240 1040 9320 1050
rect 9360 1040 9440 1050
rect 9720 1040 9760 1050
rect 9840 1040 9990 1050
rect 760 1030 800 1040
rect 1480 1030 1520 1040
rect 2080 1030 2200 1040
rect 3720 1030 3760 1040
rect 3840 1030 3880 1040
rect 4040 1030 4080 1040
rect 4200 1030 4240 1040
rect 4520 1030 4600 1040
rect 6480 1030 6560 1040
rect 6840 1030 6880 1040
rect 7320 1030 7400 1040
rect 7960 1030 8160 1040
rect 8360 1030 8560 1040
rect 9120 1030 9160 1040
rect 9240 1030 9320 1040
rect 9360 1030 9440 1040
rect 9720 1030 9760 1040
rect 9840 1030 9990 1040
rect 760 1020 800 1030
rect 1480 1020 1520 1030
rect 2080 1020 2200 1030
rect 3720 1020 3760 1030
rect 3840 1020 3880 1030
rect 4040 1020 4080 1030
rect 4200 1020 4240 1030
rect 4520 1020 4600 1030
rect 6480 1020 6560 1030
rect 6840 1020 6880 1030
rect 7320 1020 7400 1030
rect 7960 1020 8160 1030
rect 8360 1020 8560 1030
rect 9120 1020 9160 1030
rect 9240 1020 9320 1030
rect 9360 1020 9440 1030
rect 9720 1020 9760 1030
rect 9840 1020 9990 1030
rect 720 1010 800 1020
rect 1440 1010 1480 1020
rect 2040 1010 2280 1020
rect 2680 1010 2720 1020
rect 3840 1010 3880 1020
rect 4200 1010 4240 1020
rect 4680 1010 4720 1020
rect 6440 1010 6520 1020
rect 6840 1010 6880 1020
rect 7320 1010 7400 1020
rect 7960 1010 8120 1020
rect 8360 1010 8560 1020
rect 9120 1010 9160 1020
rect 9480 1010 9560 1020
rect 9720 1010 9760 1020
rect 9800 1010 9840 1020
rect 9920 1010 9960 1020
rect 720 1000 800 1010
rect 1440 1000 1480 1010
rect 2040 1000 2280 1010
rect 2680 1000 2720 1010
rect 3840 1000 3880 1010
rect 4200 1000 4240 1010
rect 4680 1000 4720 1010
rect 6440 1000 6520 1010
rect 6840 1000 6880 1010
rect 7320 1000 7400 1010
rect 7960 1000 8120 1010
rect 8360 1000 8560 1010
rect 9120 1000 9160 1010
rect 9480 1000 9560 1010
rect 9720 1000 9760 1010
rect 9800 1000 9840 1010
rect 9920 1000 9960 1010
rect 720 990 800 1000
rect 1440 990 1480 1000
rect 2040 990 2280 1000
rect 2680 990 2720 1000
rect 3840 990 3880 1000
rect 4200 990 4240 1000
rect 4680 990 4720 1000
rect 6440 990 6520 1000
rect 6840 990 6880 1000
rect 7320 990 7400 1000
rect 7960 990 8120 1000
rect 8360 990 8560 1000
rect 9120 990 9160 1000
rect 9480 990 9560 1000
rect 9720 990 9760 1000
rect 9800 990 9840 1000
rect 9920 990 9960 1000
rect 720 980 800 990
rect 1440 980 1480 990
rect 2040 980 2280 990
rect 2680 980 2720 990
rect 3840 980 3880 990
rect 4200 980 4240 990
rect 4680 980 4720 990
rect 6440 980 6520 990
rect 6840 980 6880 990
rect 7320 980 7400 990
rect 7960 980 8120 990
rect 8360 980 8560 990
rect 9120 980 9160 990
rect 9480 980 9560 990
rect 9720 980 9760 990
rect 9800 980 9840 990
rect 9920 980 9960 990
rect 720 970 800 980
rect 1400 970 1440 980
rect 2040 970 2720 980
rect 3800 970 3880 980
rect 4760 970 4800 980
rect 6480 970 6560 980
rect 6800 970 6880 980
rect 7320 970 7400 980
rect 7960 970 8120 980
rect 8360 970 8560 980
rect 9160 970 9240 980
rect 720 960 800 970
rect 1400 960 1440 970
rect 2040 960 2720 970
rect 3800 960 3880 970
rect 4760 960 4800 970
rect 6480 960 6560 970
rect 6800 960 6880 970
rect 7320 960 7400 970
rect 7960 960 8120 970
rect 8360 960 8560 970
rect 9160 960 9240 970
rect 720 950 800 960
rect 1400 950 1440 960
rect 2040 950 2720 960
rect 3800 950 3880 960
rect 4760 950 4800 960
rect 6480 950 6560 960
rect 6800 950 6880 960
rect 7320 950 7400 960
rect 7960 950 8120 960
rect 8360 950 8560 960
rect 9160 950 9240 960
rect 720 940 800 950
rect 1400 940 1440 950
rect 2040 940 2720 950
rect 3800 940 3880 950
rect 4760 940 4800 950
rect 6480 940 6560 950
rect 6800 940 6880 950
rect 7320 940 7400 950
rect 7960 940 8120 950
rect 8360 940 8560 950
rect 9160 940 9240 950
rect 720 930 760 940
rect 1360 930 1400 940
rect 2040 930 2720 940
rect 3800 930 3880 940
rect 4800 930 4840 940
rect 5360 930 5480 940
rect 5520 930 5560 940
rect 6480 930 6560 940
rect 6800 930 6880 940
rect 7320 930 7400 940
rect 7960 930 8120 940
rect 8400 930 8600 940
rect 9160 930 9200 940
rect 9440 930 9520 940
rect 720 920 760 930
rect 1360 920 1400 930
rect 2040 920 2720 930
rect 3800 920 3880 930
rect 4800 920 4840 930
rect 5360 920 5480 930
rect 5520 920 5560 930
rect 6480 920 6560 930
rect 6800 920 6880 930
rect 7320 920 7400 930
rect 7960 920 8120 930
rect 8400 920 8600 930
rect 9160 920 9200 930
rect 9440 920 9520 930
rect 720 910 760 920
rect 1360 910 1400 920
rect 2040 910 2720 920
rect 3800 910 3880 920
rect 4800 910 4840 920
rect 5360 910 5480 920
rect 5520 910 5560 920
rect 6480 910 6560 920
rect 6800 910 6880 920
rect 7320 910 7400 920
rect 7960 910 8120 920
rect 8400 910 8600 920
rect 9160 910 9200 920
rect 9440 910 9520 920
rect 720 900 760 910
rect 1360 900 1400 910
rect 2040 900 2720 910
rect 3800 900 3880 910
rect 4800 900 4840 910
rect 5360 900 5480 910
rect 5520 900 5560 910
rect 6480 900 6560 910
rect 6800 900 6880 910
rect 7320 900 7400 910
rect 7960 900 8120 910
rect 8400 900 8600 910
rect 9160 900 9200 910
rect 9440 900 9520 910
rect 680 890 760 900
rect 1280 890 1360 900
rect 2040 890 2680 900
rect 3840 890 4040 900
rect 4840 890 4880 900
rect 5360 890 5400 900
rect 6480 890 6560 900
rect 6800 890 6880 900
rect 7280 890 7400 900
rect 8000 890 8120 900
rect 8440 890 8640 900
rect 9160 890 9200 900
rect 9520 890 9560 900
rect 680 880 760 890
rect 1280 880 1360 890
rect 2040 880 2680 890
rect 3840 880 4040 890
rect 4840 880 4880 890
rect 5360 880 5400 890
rect 6480 880 6560 890
rect 6800 880 6880 890
rect 7280 880 7400 890
rect 8000 880 8120 890
rect 8440 880 8640 890
rect 9160 880 9200 890
rect 9520 880 9560 890
rect 680 870 760 880
rect 1280 870 1360 880
rect 2040 870 2680 880
rect 3840 870 4040 880
rect 4840 870 4880 880
rect 5360 870 5400 880
rect 6480 870 6560 880
rect 6800 870 6880 880
rect 7280 870 7400 880
rect 8000 870 8120 880
rect 8440 870 8640 880
rect 9160 870 9200 880
rect 9520 870 9560 880
rect 680 860 760 870
rect 1280 860 1360 870
rect 2040 860 2680 870
rect 3840 860 4040 870
rect 4840 860 4880 870
rect 5360 860 5400 870
rect 6480 860 6560 870
rect 6800 860 6880 870
rect 7280 860 7400 870
rect 8000 860 8120 870
rect 8440 860 8640 870
rect 9160 860 9200 870
rect 9520 860 9560 870
rect 680 850 760 860
rect 1240 850 1320 860
rect 2040 850 2440 860
rect 2480 850 2520 860
rect 2560 850 2640 860
rect 3880 850 4040 860
rect 4240 850 4280 860
rect 6480 850 6560 860
rect 6840 850 6880 860
rect 7280 850 7360 860
rect 8000 850 8120 860
rect 8480 850 8640 860
rect 9160 850 9200 860
rect 9440 850 9480 860
rect 680 840 760 850
rect 1240 840 1320 850
rect 2040 840 2440 850
rect 2480 840 2520 850
rect 2560 840 2640 850
rect 3880 840 4040 850
rect 4240 840 4280 850
rect 6480 840 6560 850
rect 6840 840 6880 850
rect 7280 840 7360 850
rect 8000 840 8120 850
rect 8480 840 8640 850
rect 9160 840 9200 850
rect 9440 840 9480 850
rect 680 830 760 840
rect 1240 830 1320 840
rect 2040 830 2440 840
rect 2480 830 2520 840
rect 2560 830 2640 840
rect 3880 830 4040 840
rect 4240 830 4280 840
rect 6480 830 6560 840
rect 6840 830 6880 840
rect 7280 830 7360 840
rect 8000 830 8120 840
rect 8480 830 8640 840
rect 9160 830 9200 840
rect 9440 830 9480 840
rect 680 820 760 830
rect 1240 820 1320 830
rect 2040 820 2440 830
rect 2480 820 2520 830
rect 2560 820 2640 830
rect 3880 820 4040 830
rect 4240 820 4280 830
rect 6480 820 6560 830
rect 6840 820 6880 830
rect 7280 820 7360 830
rect 8000 820 8120 830
rect 8480 820 8640 830
rect 9160 820 9200 830
rect 9440 820 9480 830
rect 680 810 760 820
rect 1200 810 1280 820
rect 2040 810 2360 820
rect 2440 810 2480 820
rect 4000 810 4040 820
rect 4280 810 4360 820
rect 4880 810 4920 820
rect 6520 810 6600 820
rect 6840 810 6880 820
rect 7280 810 7360 820
rect 8000 810 8120 820
rect 9360 810 9400 820
rect 680 800 760 810
rect 1200 800 1280 810
rect 2040 800 2360 810
rect 2440 800 2480 810
rect 4000 800 4040 810
rect 4280 800 4360 810
rect 4880 800 4920 810
rect 6520 800 6600 810
rect 6840 800 6880 810
rect 7280 800 7360 810
rect 8000 800 8120 810
rect 9360 800 9400 810
rect 680 790 760 800
rect 1200 790 1280 800
rect 2040 790 2360 800
rect 2440 790 2480 800
rect 4000 790 4040 800
rect 4280 790 4360 800
rect 4880 790 4920 800
rect 6520 790 6600 800
rect 6840 790 6880 800
rect 7280 790 7360 800
rect 8000 790 8120 800
rect 9360 790 9400 800
rect 680 780 760 790
rect 1200 780 1280 790
rect 2040 780 2360 790
rect 2440 780 2480 790
rect 4000 780 4040 790
rect 4280 780 4360 790
rect 4880 780 4920 790
rect 6520 780 6600 790
rect 6840 780 6880 790
rect 7280 780 7360 790
rect 8000 780 8120 790
rect 9360 780 9400 790
rect 640 770 720 780
rect 1160 770 1240 780
rect 2080 770 2320 780
rect 2480 770 2520 780
rect 3560 770 3720 780
rect 3760 770 3800 780
rect 3840 770 3880 780
rect 4000 770 4040 780
rect 4320 770 4360 780
rect 6520 770 6600 780
rect 6840 770 6880 780
rect 7280 770 7360 780
rect 8000 770 8120 780
rect 9200 770 9240 780
rect 640 760 720 770
rect 1160 760 1240 770
rect 2080 760 2320 770
rect 2480 760 2520 770
rect 3560 760 3720 770
rect 3760 760 3800 770
rect 3840 760 3880 770
rect 4000 760 4040 770
rect 4320 760 4360 770
rect 6520 760 6600 770
rect 6840 760 6880 770
rect 7280 760 7360 770
rect 8000 760 8120 770
rect 9200 760 9240 770
rect 640 750 720 760
rect 1160 750 1240 760
rect 2080 750 2320 760
rect 2480 750 2520 760
rect 3560 750 3720 760
rect 3760 750 3800 760
rect 3840 750 3880 760
rect 4000 750 4040 760
rect 4320 750 4360 760
rect 6520 750 6600 760
rect 6840 750 6880 760
rect 7280 750 7360 760
rect 8000 750 8120 760
rect 9200 750 9240 760
rect 640 740 720 750
rect 1160 740 1240 750
rect 2080 740 2320 750
rect 2480 740 2520 750
rect 3560 740 3720 750
rect 3760 740 3800 750
rect 3840 740 3880 750
rect 4000 740 4040 750
rect 4320 740 4360 750
rect 6520 740 6600 750
rect 6840 740 6880 750
rect 7280 740 7360 750
rect 8000 740 8120 750
rect 9200 740 9240 750
rect 640 730 720 740
rect 1080 730 1200 740
rect 2080 730 2240 740
rect 2400 730 2440 740
rect 3400 730 3480 740
rect 4040 730 4200 740
rect 4720 730 4800 740
rect 6560 730 6600 740
rect 6880 730 6920 740
rect 7280 730 7360 740
rect 8000 730 8120 740
rect 9200 730 9240 740
rect 9320 730 9400 740
rect 640 720 720 730
rect 1080 720 1200 730
rect 2080 720 2240 730
rect 2400 720 2440 730
rect 3400 720 3480 730
rect 4040 720 4200 730
rect 4720 720 4800 730
rect 6560 720 6600 730
rect 6880 720 6920 730
rect 7280 720 7360 730
rect 8000 720 8120 730
rect 9200 720 9240 730
rect 9320 720 9400 730
rect 640 710 720 720
rect 1080 710 1200 720
rect 2080 710 2240 720
rect 2400 710 2440 720
rect 3400 710 3480 720
rect 4040 710 4200 720
rect 4720 710 4800 720
rect 6560 710 6600 720
rect 6880 710 6920 720
rect 7280 710 7360 720
rect 8000 710 8120 720
rect 9200 710 9240 720
rect 9320 710 9400 720
rect 640 700 720 710
rect 1080 700 1200 710
rect 2080 700 2240 710
rect 2400 700 2440 710
rect 3400 700 3480 710
rect 4040 700 4200 710
rect 4720 700 4800 710
rect 6560 700 6600 710
rect 6880 700 6920 710
rect 7280 700 7360 710
rect 8000 700 8120 710
rect 9200 700 9240 710
rect 9320 700 9400 710
rect 640 690 680 700
rect 1040 690 1200 700
rect 2120 690 2240 700
rect 2320 690 2360 700
rect 3320 690 3360 700
rect 4040 690 4120 700
rect 4160 690 4200 700
rect 4800 690 4840 700
rect 6560 690 6640 700
rect 6840 690 6920 700
rect 7240 690 7360 700
rect 8040 690 8120 700
rect 9200 690 9240 700
rect 640 680 680 690
rect 1040 680 1200 690
rect 2120 680 2240 690
rect 2320 680 2360 690
rect 3320 680 3360 690
rect 4040 680 4120 690
rect 4160 680 4200 690
rect 4800 680 4840 690
rect 6560 680 6640 690
rect 6840 680 6920 690
rect 7240 680 7360 690
rect 8040 680 8120 690
rect 9200 680 9240 690
rect 640 670 680 680
rect 1040 670 1200 680
rect 2120 670 2240 680
rect 2320 670 2360 680
rect 3320 670 3360 680
rect 4040 670 4120 680
rect 4160 670 4200 680
rect 4800 670 4840 680
rect 6560 670 6640 680
rect 6840 670 6920 680
rect 7240 670 7360 680
rect 8040 670 8120 680
rect 9200 670 9240 680
rect 640 660 680 670
rect 1040 660 1200 670
rect 2120 660 2240 670
rect 2320 660 2360 670
rect 3320 660 3360 670
rect 4040 660 4120 670
rect 4160 660 4200 670
rect 4800 660 4840 670
rect 6560 660 6640 670
rect 6840 660 6920 670
rect 7240 660 7360 670
rect 8040 660 8120 670
rect 9200 660 9240 670
rect 720 650 760 660
rect 1000 650 1160 660
rect 2120 650 2280 660
rect 4080 650 4120 660
rect 4680 650 4720 660
rect 4800 650 4840 660
rect 6600 650 6680 660
rect 6840 650 6960 660
rect 7240 650 7320 660
rect 8040 650 8120 660
rect 9160 650 9240 660
rect 9280 650 9360 660
rect 9600 650 9720 660
rect 720 640 760 650
rect 1000 640 1160 650
rect 2120 640 2280 650
rect 4080 640 4120 650
rect 4680 640 4720 650
rect 4800 640 4840 650
rect 6600 640 6680 650
rect 6840 640 6960 650
rect 7240 640 7320 650
rect 8040 640 8120 650
rect 9160 640 9240 650
rect 9280 640 9360 650
rect 9600 640 9720 650
rect 720 630 760 640
rect 1000 630 1160 640
rect 2120 630 2280 640
rect 4080 630 4120 640
rect 4680 630 4720 640
rect 4800 630 4840 640
rect 6600 630 6680 640
rect 6840 630 6960 640
rect 7240 630 7320 640
rect 8040 630 8120 640
rect 9160 630 9240 640
rect 9280 630 9360 640
rect 9600 630 9720 640
rect 720 620 760 630
rect 1000 620 1160 630
rect 2120 620 2280 630
rect 4080 620 4120 630
rect 4680 620 4720 630
rect 4800 620 4840 630
rect 6600 620 6680 630
rect 6840 620 6960 630
rect 7240 620 7320 630
rect 8040 620 8120 630
rect 9160 620 9240 630
rect 9280 620 9360 630
rect 9600 620 9720 630
rect 440 610 480 620
rect 560 610 640 620
rect 720 610 760 620
rect 920 610 1080 620
rect 2160 610 2200 620
rect 3120 610 3200 620
rect 4040 610 4080 620
rect 4520 610 4560 620
rect 4680 610 4720 620
rect 4760 610 4800 620
rect 4920 610 4960 620
rect 6600 610 6720 620
rect 6920 610 7000 620
rect 7200 610 7320 620
rect 9160 610 9280 620
rect 440 600 480 610
rect 560 600 640 610
rect 720 600 760 610
rect 920 600 1080 610
rect 2160 600 2200 610
rect 3120 600 3200 610
rect 4040 600 4080 610
rect 4520 600 4560 610
rect 4680 600 4720 610
rect 4760 600 4800 610
rect 4920 600 4960 610
rect 6600 600 6720 610
rect 6920 600 7000 610
rect 7200 600 7320 610
rect 9160 600 9280 610
rect 440 590 480 600
rect 560 590 640 600
rect 720 590 760 600
rect 920 590 1080 600
rect 2160 590 2200 600
rect 3120 590 3200 600
rect 4040 590 4080 600
rect 4520 590 4560 600
rect 4680 590 4720 600
rect 4760 590 4800 600
rect 4920 590 4960 600
rect 6600 590 6720 600
rect 6920 590 7000 600
rect 7200 590 7320 600
rect 9160 590 9280 600
rect 440 580 480 590
rect 560 580 640 590
rect 720 580 760 590
rect 920 580 1080 590
rect 2160 580 2200 590
rect 3120 580 3200 590
rect 4040 580 4080 590
rect 4520 580 4560 590
rect 4680 580 4720 590
rect 4760 580 4800 590
rect 4920 580 4960 590
rect 6600 580 6720 590
rect 6920 580 7000 590
rect 7200 580 7320 590
rect 9160 580 9280 590
rect 600 570 640 580
rect 920 570 1040 580
rect 1280 570 1440 580
rect 3000 570 3120 580
rect 4360 570 4480 580
rect 4640 570 4680 580
rect 4760 570 4800 580
rect 4840 570 4880 580
rect 4920 570 4960 580
rect 6640 570 6720 580
rect 6920 570 7040 580
rect 7160 570 7320 580
rect 9200 570 9240 580
rect 9280 570 9320 580
rect 600 560 640 570
rect 920 560 1040 570
rect 1280 560 1440 570
rect 3000 560 3120 570
rect 4360 560 4480 570
rect 4640 560 4680 570
rect 4760 560 4800 570
rect 4840 560 4880 570
rect 4920 560 4960 570
rect 6640 560 6720 570
rect 6920 560 7040 570
rect 7160 560 7320 570
rect 9200 560 9240 570
rect 9280 560 9320 570
rect 600 550 640 560
rect 920 550 1040 560
rect 1280 550 1440 560
rect 3000 550 3120 560
rect 4360 550 4480 560
rect 4640 550 4680 560
rect 4760 550 4800 560
rect 4840 550 4880 560
rect 4920 550 4960 560
rect 6640 550 6720 560
rect 6920 550 7040 560
rect 7160 550 7320 560
rect 9200 550 9240 560
rect 9280 550 9320 560
rect 600 540 640 550
rect 920 540 1040 550
rect 1280 540 1440 550
rect 3000 540 3120 550
rect 4360 540 4480 550
rect 4640 540 4680 550
rect 4760 540 4800 550
rect 4840 540 4880 550
rect 4920 540 4960 550
rect 6640 540 6720 550
rect 6920 540 7040 550
rect 7160 540 7320 550
rect 9200 540 9240 550
rect 9280 540 9320 550
rect 520 530 640 540
rect 960 530 1040 540
rect 1240 530 1280 540
rect 2960 530 3000 540
rect 4240 530 4360 540
rect 4560 530 4640 540
rect 4760 530 4800 540
rect 6640 530 6760 540
rect 6880 530 7080 540
rect 7120 530 7280 540
rect 9200 530 9240 540
rect 9920 530 9990 540
rect 520 520 640 530
rect 960 520 1040 530
rect 1240 520 1280 530
rect 2960 520 3000 530
rect 4240 520 4360 530
rect 4560 520 4640 530
rect 4760 520 4800 530
rect 6640 520 6760 530
rect 6880 520 7080 530
rect 7120 520 7280 530
rect 9200 520 9240 530
rect 9920 520 9990 530
rect 520 510 640 520
rect 960 510 1040 520
rect 1240 510 1280 520
rect 2960 510 3000 520
rect 4240 510 4360 520
rect 4560 510 4640 520
rect 4760 510 4800 520
rect 6640 510 6760 520
rect 6880 510 7080 520
rect 7120 510 7280 520
rect 9200 510 9240 520
rect 9920 510 9990 520
rect 520 500 640 510
rect 960 500 1040 510
rect 1240 500 1280 510
rect 2960 500 3000 510
rect 4240 500 4360 510
rect 4560 500 4640 510
rect 4760 500 4800 510
rect 6640 500 6760 510
rect 6880 500 7080 510
rect 7120 500 7280 510
rect 9200 500 9240 510
rect 9920 500 9990 510
rect 160 490 320 500
rect 360 490 400 500
rect 440 490 520 500
rect 1160 490 1200 500
rect 2800 490 2880 500
rect 4200 490 4240 500
rect 4760 490 4800 500
rect 4880 490 4920 500
rect 6680 490 6760 500
rect 6880 490 7280 500
rect 9160 490 9200 500
rect 9880 490 9960 500
rect 160 480 320 490
rect 360 480 400 490
rect 440 480 520 490
rect 1160 480 1200 490
rect 2800 480 2880 490
rect 4200 480 4240 490
rect 4760 480 4800 490
rect 4880 480 4920 490
rect 6680 480 6760 490
rect 6880 480 7280 490
rect 9160 480 9200 490
rect 9880 480 9960 490
rect 160 470 320 480
rect 360 470 400 480
rect 440 470 520 480
rect 1160 470 1200 480
rect 2800 470 2880 480
rect 4200 470 4240 480
rect 4760 470 4800 480
rect 4880 470 4920 480
rect 6680 470 6760 480
rect 6880 470 7280 480
rect 9160 470 9200 480
rect 9880 470 9960 480
rect 160 460 320 470
rect 360 460 400 470
rect 440 460 520 470
rect 1160 460 1200 470
rect 2800 460 2880 470
rect 4200 460 4240 470
rect 4760 460 4800 470
rect 4880 460 4920 470
rect 6680 460 6760 470
rect 6880 460 7280 470
rect 9160 460 9200 470
rect 9880 460 9960 470
rect 280 450 360 460
rect 440 450 480 460
rect 1120 450 1160 460
rect 1960 450 2040 460
rect 2240 450 2280 460
rect 2640 450 2720 460
rect 4160 450 4200 460
rect 4880 450 4920 460
rect 6720 450 7240 460
rect 9120 450 9160 460
rect 9200 450 9240 460
rect 9280 450 9360 460
rect 280 440 360 450
rect 440 440 480 450
rect 1120 440 1160 450
rect 1960 440 2040 450
rect 2240 440 2280 450
rect 2640 440 2720 450
rect 4160 440 4200 450
rect 4880 440 4920 450
rect 6720 440 7240 450
rect 9120 440 9160 450
rect 9200 440 9240 450
rect 9280 440 9360 450
rect 280 430 360 440
rect 440 430 480 440
rect 1120 430 1160 440
rect 1960 430 2040 440
rect 2240 430 2280 440
rect 2640 430 2720 440
rect 4160 430 4200 440
rect 4880 430 4920 440
rect 6720 430 7240 440
rect 9120 430 9160 440
rect 9200 430 9240 440
rect 9280 430 9360 440
rect 280 420 360 430
rect 440 420 480 430
rect 1120 420 1160 430
rect 1960 420 2040 430
rect 2240 420 2280 430
rect 2640 420 2720 430
rect 4160 420 4200 430
rect 4880 420 4920 430
rect 6720 420 7240 430
rect 9120 420 9160 430
rect 9200 420 9240 430
rect 9280 420 9360 430
rect 280 410 400 420
rect 440 410 480 420
rect 1080 410 1120 420
rect 4160 410 4200 420
rect 4720 410 4760 420
rect 6720 410 7240 420
rect 9120 410 9160 420
rect 9280 410 9320 420
rect 9360 410 9400 420
rect 280 400 400 410
rect 440 400 480 410
rect 1080 400 1120 410
rect 4160 400 4200 410
rect 4720 400 4760 410
rect 6720 400 7240 410
rect 9120 400 9160 410
rect 9280 400 9320 410
rect 9360 400 9400 410
rect 280 390 400 400
rect 440 390 480 400
rect 1080 390 1120 400
rect 4160 390 4200 400
rect 4720 390 4760 400
rect 6720 390 7240 400
rect 9120 390 9160 400
rect 9280 390 9320 400
rect 9360 390 9400 400
rect 280 380 400 390
rect 440 380 480 390
rect 1080 380 1120 390
rect 4160 380 4200 390
rect 4720 380 4760 390
rect 6720 380 7240 390
rect 9120 380 9160 390
rect 9280 380 9320 390
rect 9360 380 9400 390
rect 40 370 80 380
rect 280 370 400 380
rect 4120 370 4200 380
rect 4320 370 4360 380
rect 4720 370 4760 380
rect 4920 370 4960 380
rect 6760 370 7200 380
rect 9160 370 9200 380
rect 9400 370 9440 380
rect 40 360 80 370
rect 280 360 400 370
rect 4120 360 4200 370
rect 4320 360 4360 370
rect 4720 360 4760 370
rect 4920 360 4960 370
rect 6760 360 7200 370
rect 9160 360 9200 370
rect 9400 360 9440 370
rect 40 350 80 360
rect 280 350 400 360
rect 4120 350 4200 360
rect 4320 350 4360 360
rect 4720 350 4760 360
rect 4920 350 4960 360
rect 6760 350 7200 360
rect 9160 350 9200 360
rect 9400 350 9440 360
rect 40 340 80 350
rect 280 340 400 350
rect 4120 340 4200 350
rect 4320 340 4360 350
rect 4720 340 4760 350
rect 4920 340 4960 350
rect 6760 340 7200 350
rect 9160 340 9200 350
rect 9400 340 9440 350
rect 80 330 120 340
rect 240 330 400 340
rect 480 330 720 340
rect 4080 330 4200 340
rect 4240 330 4400 340
rect 4760 330 4960 340
rect 6840 330 7160 340
rect 9080 330 9120 340
rect 9200 330 9240 340
rect 9400 330 9440 340
rect 80 320 120 330
rect 240 320 400 330
rect 480 320 720 330
rect 4080 320 4200 330
rect 4240 320 4400 330
rect 4760 320 4960 330
rect 6840 320 7160 330
rect 9080 320 9120 330
rect 9200 320 9240 330
rect 9400 320 9440 330
rect 80 310 120 320
rect 240 310 400 320
rect 480 310 720 320
rect 4080 310 4200 320
rect 4240 310 4400 320
rect 4760 310 4960 320
rect 6840 310 7160 320
rect 9080 310 9120 320
rect 9200 310 9240 320
rect 9400 310 9440 320
rect 80 300 120 310
rect 240 300 400 310
rect 480 300 720 310
rect 4080 300 4200 310
rect 4240 300 4400 310
rect 4760 300 4960 310
rect 6840 300 7160 310
rect 9080 300 9120 310
rect 9200 300 9240 310
rect 9400 300 9440 310
rect 40 290 400 300
rect 440 290 520 300
rect 560 290 640 300
rect 680 290 840 300
rect 4080 290 4120 300
rect 4200 290 4520 300
rect 4680 290 5000 300
rect 6920 290 7040 300
rect 9040 290 9080 300
rect 9400 290 9480 300
rect 40 280 400 290
rect 440 280 520 290
rect 560 280 640 290
rect 680 280 840 290
rect 4080 280 4120 290
rect 4200 280 4520 290
rect 4680 280 5000 290
rect 6920 280 7040 290
rect 9040 280 9080 290
rect 9400 280 9480 290
rect 40 270 400 280
rect 440 270 520 280
rect 560 270 640 280
rect 680 270 840 280
rect 4080 270 4120 280
rect 4200 270 4520 280
rect 4680 270 5000 280
rect 6920 270 7040 280
rect 9040 270 9080 280
rect 9400 270 9480 280
rect 40 260 400 270
rect 440 260 520 270
rect 560 260 640 270
rect 680 260 840 270
rect 4080 260 4120 270
rect 4200 260 4520 270
rect 4680 260 5000 270
rect 6920 260 7040 270
rect 9040 260 9080 270
rect 9400 260 9480 270
rect 0 250 120 260
rect 200 250 400 260
rect 440 250 640 260
rect 680 250 880 260
rect 1000 250 1040 260
rect 4080 250 4120 260
rect 4160 250 4560 260
rect 4640 250 4960 260
rect 8880 250 8960 260
rect 9040 250 9080 260
rect 9160 250 9200 260
rect 9320 250 9480 260
rect 9800 250 9840 260
rect 0 240 120 250
rect 200 240 400 250
rect 440 240 640 250
rect 680 240 880 250
rect 1000 240 1040 250
rect 4080 240 4120 250
rect 4160 240 4560 250
rect 4640 240 4960 250
rect 8880 240 8960 250
rect 9040 240 9080 250
rect 9160 240 9200 250
rect 9320 240 9480 250
rect 9800 240 9840 250
rect 0 230 120 240
rect 200 230 400 240
rect 440 230 640 240
rect 680 230 880 240
rect 1000 230 1040 240
rect 4080 230 4120 240
rect 4160 230 4560 240
rect 4640 230 4960 240
rect 8880 230 8960 240
rect 9040 230 9080 240
rect 9160 230 9200 240
rect 9320 230 9480 240
rect 9800 230 9840 240
rect 0 220 120 230
rect 200 220 400 230
rect 440 220 640 230
rect 680 220 880 230
rect 1000 220 1040 230
rect 4080 220 4120 230
rect 4160 220 4560 230
rect 4640 220 4960 230
rect 8880 220 8960 230
rect 9040 220 9080 230
rect 9160 220 9200 230
rect 9320 220 9480 230
rect 9800 220 9840 230
rect 0 210 80 220
rect 240 210 360 220
rect 440 210 600 220
rect 680 210 880 220
rect 1000 210 1040 220
rect 4120 210 4160 220
rect 4240 210 4320 220
rect 4400 210 4560 220
rect 4600 210 4920 220
rect 8880 210 8920 220
rect 9000 210 9040 220
rect 9120 210 9160 220
rect 9280 210 9360 220
rect 9720 210 9800 220
rect 9840 210 9990 220
rect 0 200 80 210
rect 240 200 360 210
rect 440 200 600 210
rect 680 200 880 210
rect 1000 200 1040 210
rect 4120 200 4160 210
rect 4240 200 4320 210
rect 4400 200 4560 210
rect 4600 200 4920 210
rect 8880 200 8920 210
rect 9000 200 9040 210
rect 9120 200 9160 210
rect 9280 200 9360 210
rect 9720 200 9800 210
rect 9840 200 9990 210
rect 0 190 80 200
rect 240 190 360 200
rect 440 190 600 200
rect 680 190 880 200
rect 1000 190 1040 200
rect 4120 190 4160 200
rect 4240 190 4320 200
rect 4400 190 4560 200
rect 4600 190 4920 200
rect 8880 190 8920 200
rect 9000 190 9040 200
rect 9120 190 9160 200
rect 9280 190 9360 200
rect 9720 190 9800 200
rect 9840 190 9990 200
rect 0 180 80 190
rect 240 180 360 190
rect 440 180 600 190
rect 680 180 880 190
rect 1000 180 1040 190
rect 4120 180 4160 190
rect 4240 180 4320 190
rect 4400 180 4560 190
rect 4600 180 4920 190
rect 8880 180 8920 190
rect 9000 180 9040 190
rect 9120 180 9160 190
rect 9280 180 9360 190
rect 9720 180 9800 190
rect 9840 180 9990 190
rect 0 170 120 180
rect 240 170 280 180
rect 720 170 800 180
rect 1000 170 1040 180
rect 4160 170 4200 180
rect 4560 170 4840 180
rect 4920 170 4960 180
rect 8840 170 8880 180
rect 9000 170 9040 180
rect 9120 170 9160 180
rect 9320 170 9360 180
rect 9720 170 9760 180
rect 0 160 120 170
rect 240 160 280 170
rect 720 160 800 170
rect 1000 160 1040 170
rect 4160 160 4200 170
rect 4560 160 4840 170
rect 4920 160 4960 170
rect 8840 160 8880 170
rect 9000 160 9040 170
rect 9120 160 9160 170
rect 9320 160 9360 170
rect 9720 160 9760 170
rect 0 150 120 160
rect 240 150 280 160
rect 720 150 800 160
rect 1000 150 1040 160
rect 4160 150 4200 160
rect 4560 150 4840 160
rect 4920 150 4960 160
rect 8840 150 8880 160
rect 9000 150 9040 160
rect 9120 150 9160 160
rect 9320 150 9360 160
rect 9720 150 9760 160
rect 0 140 120 150
rect 240 140 280 150
rect 720 140 800 150
rect 1000 140 1040 150
rect 4160 140 4200 150
rect 4560 140 4840 150
rect 4920 140 4960 150
rect 8840 140 8880 150
rect 9000 140 9040 150
rect 9120 140 9160 150
rect 9320 140 9360 150
rect 9720 140 9760 150
rect 0 130 120 140
rect 1000 130 1040 140
rect 4200 130 4240 140
rect 4560 130 4600 140
rect 4640 130 4680 140
rect 4720 130 4800 140
rect 5000 130 5040 140
rect 9080 130 9160 140
rect 9360 130 9400 140
rect 0 120 120 130
rect 1000 120 1040 130
rect 4200 120 4240 130
rect 4560 120 4600 130
rect 4640 120 4680 130
rect 4720 120 4800 130
rect 5000 120 5040 130
rect 9080 120 9160 130
rect 9360 120 9400 130
rect 0 110 120 120
rect 1000 110 1040 120
rect 4200 110 4240 120
rect 4560 110 4600 120
rect 4640 110 4680 120
rect 4720 110 4800 120
rect 5000 110 5040 120
rect 9080 110 9160 120
rect 9360 110 9400 120
rect 0 100 120 110
rect 1000 100 1040 110
rect 4200 100 4240 110
rect 4560 100 4600 110
rect 4640 100 4680 110
rect 4720 100 4800 110
rect 5000 100 5040 110
rect 9080 100 9160 110
rect 9360 100 9400 110
rect 0 90 120 100
rect 1000 90 1040 100
rect 4240 90 4280 100
rect 4920 90 4960 100
rect 8760 90 8800 100
rect 8920 90 8960 100
rect 9120 90 9160 100
rect 9440 90 9480 100
rect 9560 90 9600 100
rect 9680 90 9760 100
rect 9920 90 9960 100
rect 0 80 120 90
rect 1000 80 1040 90
rect 4240 80 4280 90
rect 4920 80 4960 90
rect 8760 80 8800 90
rect 8920 80 8960 90
rect 9120 80 9160 90
rect 9440 80 9480 90
rect 9560 80 9600 90
rect 9680 80 9760 90
rect 9920 80 9960 90
rect 0 70 120 80
rect 1000 70 1040 80
rect 4240 70 4280 80
rect 4920 70 4960 80
rect 8760 70 8800 80
rect 8920 70 8960 80
rect 9120 70 9160 80
rect 9440 70 9480 80
rect 9560 70 9600 80
rect 9680 70 9760 80
rect 9920 70 9960 80
rect 0 60 120 70
rect 1000 60 1040 70
rect 4240 60 4280 70
rect 4920 60 4960 70
rect 8760 60 8800 70
rect 8920 60 8960 70
rect 9120 60 9160 70
rect 9440 60 9480 70
rect 9560 60 9600 70
rect 9680 60 9760 70
rect 9920 60 9960 70
rect 40 50 120 60
rect 1000 50 1040 60
rect 4320 50 4360 60
rect 4920 50 4960 60
rect 9000 50 9040 60
rect 9080 50 9120 60
rect 9480 50 9760 60
rect 9920 50 9990 60
rect 40 40 120 50
rect 1000 40 1040 50
rect 4320 40 4360 50
rect 4920 40 4960 50
rect 9000 40 9040 50
rect 9080 40 9120 50
rect 9480 40 9760 50
rect 9920 40 9990 50
rect 40 30 120 40
rect 1000 30 1040 40
rect 4320 30 4360 40
rect 4920 30 4960 40
rect 9000 30 9040 40
rect 9080 30 9120 40
rect 9480 30 9760 40
rect 9920 30 9990 40
rect 40 20 120 30
rect 1000 20 1040 30
rect 4320 20 4360 30
rect 4920 20 4960 30
rect 9000 20 9040 30
rect 9080 20 9120 30
rect 9480 20 9760 30
rect 9920 20 9990 30
rect 0 10 80 20
rect 1000 10 1040 20
rect 4920 10 4960 20
rect 5040 10 5080 20
rect 8600 10 8680 20
rect 8880 10 8920 20
rect 9080 10 9120 20
rect 9160 10 9200 20
rect 9480 10 9800 20
rect 9920 10 9960 20
rect 0 0 80 10
rect 1000 0 1040 10
rect 4920 0 4960 10
rect 5040 0 5080 10
rect 8600 0 8680 10
rect 8880 0 8920 10
rect 9080 0 9120 10
rect 9160 0 9200 10
rect 9480 0 9800 10
rect 9920 0 9960 10
<< metal4 >>
rect 0 7490 2120 7500
rect 3360 7490 3560 7500
rect 3840 7490 9520 7500
rect 0 7480 2120 7490
rect 3360 7480 3560 7490
rect 3840 7480 9520 7490
rect 0 7470 2120 7480
rect 3360 7470 3560 7480
rect 3840 7470 9520 7480
rect 0 7460 2120 7470
rect 3360 7460 3560 7470
rect 3840 7460 9520 7470
rect 0 7450 2080 7460
rect 3320 7450 3560 7460
rect 3680 7450 3800 7460
rect 3840 7450 9560 7460
rect 0 7440 2080 7450
rect 3320 7440 3560 7450
rect 3680 7440 3800 7450
rect 3840 7440 9560 7450
rect 0 7430 2080 7440
rect 3320 7430 3560 7440
rect 3680 7430 3800 7440
rect 3840 7430 9560 7440
rect 0 7420 2080 7430
rect 3320 7420 3560 7430
rect 3680 7420 3800 7430
rect 3840 7420 9560 7430
rect 0 7410 2080 7420
rect 3360 7410 3600 7420
rect 3640 7410 3800 7420
rect 3880 7410 9560 7420
rect 0 7400 2080 7410
rect 3360 7400 3600 7410
rect 3640 7400 3800 7410
rect 3880 7400 9560 7410
rect 0 7390 2080 7400
rect 3360 7390 3600 7400
rect 3640 7390 3800 7400
rect 3880 7390 9560 7400
rect 0 7380 2080 7390
rect 3360 7380 3600 7390
rect 3640 7380 3800 7390
rect 3880 7380 9560 7390
rect 0 7370 2040 7380
rect 3360 7370 3840 7380
rect 3880 7370 9560 7380
rect 0 7360 2040 7370
rect 3360 7360 3840 7370
rect 3880 7360 9560 7370
rect 0 7350 2040 7360
rect 3360 7350 3840 7360
rect 3880 7350 9560 7360
rect 0 7340 2040 7350
rect 3360 7340 3840 7350
rect 3880 7340 9560 7350
rect 0 7330 2000 7340
rect 3360 7330 9560 7340
rect 0 7320 2000 7330
rect 3360 7320 9560 7330
rect 0 7310 2000 7320
rect 3360 7310 9560 7320
rect 0 7300 2000 7310
rect 3360 7300 9560 7310
rect 0 7290 2000 7300
rect 3440 7290 3840 7300
rect 3920 7290 9560 7300
rect 0 7280 2000 7290
rect 3440 7280 3840 7290
rect 3920 7280 9560 7290
rect 0 7270 2000 7280
rect 3440 7270 3840 7280
rect 3920 7270 9560 7280
rect 0 7260 2000 7270
rect 3440 7260 3840 7270
rect 3920 7260 9560 7270
rect 0 7250 1960 7260
rect 3440 7250 3800 7260
rect 3920 7250 9560 7260
rect 0 7240 1960 7250
rect 3440 7240 3800 7250
rect 3920 7240 9560 7250
rect 0 7230 1960 7240
rect 3440 7230 3800 7240
rect 3920 7230 9560 7240
rect 0 7220 1960 7230
rect 3440 7220 3800 7230
rect 3920 7220 9560 7230
rect 0 7210 1920 7220
rect 3440 7210 3800 7220
rect 3920 7210 9560 7220
rect 0 7200 1920 7210
rect 3440 7200 3800 7210
rect 3920 7200 9560 7210
rect 0 7190 1920 7200
rect 3440 7190 3800 7200
rect 3920 7190 9560 7200
rect 0 7180 1920 7190
rect 3440 7180 3800 7190
rect 3920 7180 9560 7190
rect 0 7170 1920 7180
rect 3400 7170 3720 7180
rect 3760 7170 3800 7180
rect 3960 7170 9560 7180
rect 0 7160 1920 7170
rect 3400 7160 3720 7170
rect 3760 7160 3800 7170
rect 3960 7160 9560 7170
rect 0 7150 1920 7160
rect 3400 7150 3720 7160
rect 3760 7150 3800 7160
rect 3960 7150 9560 7160
rect 0 7140 1920 7150
rect 3400 7140 3720 7150
rect 3760 7140 3800 7150
rect 3960 7140 9560 7150
rect 0 7130 1920 7140
rect 3480 7130 3520 7140
rect 3560 7130 3640 7140
rect 3960 7130 9560 7140
rect 0 7120 1920 7130
rect 3480 7120 3520 7130
rect 3560 7120 3640 7130
rect 3960 7120 9560 7130
rect 0 7110 1920 7120
rect 3480 7110 3520 7120
rect 3560 7110 3640 7120
rect 3960 7110 9560 7120
rect 0 7100 1920 7110
rect 3480 7100 3520 7110
rect 3560 7100 3640 7110
rect 3960 7100 9560 7110
rect 0 7090 1880 7100
rect 3960 7090 9560 7100
rect 0 7080 1880 7090
rect 3960 7080 9560 7090
rect 0 7070 1880 7080
rect 3960 7070 9560 7080
rect 0 7060 1880 7070
rect 3960 7060 9560 7070
rect 0 7050 1880 7060
rect 3560 7050 3640 7060
rect 3960 7050 9560 7060
rect 0 7040 1880 7050
rect 3560 7040 3640 7050
rect 3960 7040 9560 7050
rect 0 7030 1880 7040
rect 3560 7030 3640 7040
rect 3960 7030 9560 7040
rect 0 7020 1880 7030
rect 3560 7020 3640 7030
rect 3960 7020 9560 7030
rect 0 7010 1880 7020
rect 3760 7010 3800 7020
rect 4000 7010 9560 7020
rect 0 7000 1880 7010
rect 3760 7000 3800 7010
rect 4000 7000 9560 7010
rect 0 6990 1880 7000
rect 3760 6990 3800 7000
rect 4000 6990 9560 7000
rect 0 6980 1880 6990
rect 3760 6980 3800 6990
rect 4000 6980 9560 6990
rect 0 6970 1920 6980
rect 3760 6970 3800 6980
rect 4000 6970 9600 6980
rect 0 6960 1920 6970
rect 3760 6960 3800 6970
rect 4000 6960 9600 6970
rect 0 6950 1920 6960
rect 3760 6950 3800 6960
rect 4000 6950 9600 6960
rect 0 6940 1920 6950
rect 3760 6940 3800 6950
rect 4000 6940 9600 6950
rect 0 6930 1880 6940
rect 4000 6930 9600 6940
rect 0 6920 1880 6930
rect 4000 6920 9600 6930
rect 0 6910 1880 6920
rect 4000 6910 9600 6920
rect 0 6900 1880 6910
rect 4000 6900 9600 6910
rect 0 6890 1880 6900
rect 3400 6890 3480 6900
rect 4000 6890 9600 6900
rect 0 6880 1880 6890
rect 3400 6880 3480 6890
rect 4000 6880 9600 6890
rect 0 6870 1880 6880
rect 3400 6870 3480 6880
rect 4000 6870 9600 6880
rect 0 6860 1880 6870
rect 3400 6860 3480 6870
rect 4000 6860 9600 6870
rect 0 6850 1880 6860
rect 3440 6850 3560 6860
rect 3960 6850 9600 6860
rect 0 6840 1880 6850
rect 3440 6840 3560 6850
rect 3960 6840 9600 6850
rect 0 6830 1880 6840
rect 3440 6830 3560 6840
rect 3960 6830 9600 6840
rect 0 6820 1880 6830
rect 3440 6820 3560 6830
rect 3960 6820 9600 6830
rect 0 6810 1840 6820
rect 3280 6810 3640 6820
rect 3960 6810 9600 6820
rect 0 6800 1840 6810
rect 3280 6800 3640 6810
rect 3960 6800 9600 6810
rect 0 6790 1840 6800
rect 3280 6790 3640 6800
rect 3960 6790 9600 6800
rect 0 6780 1840 6790
rect 3280 6780 3640 6790
rect 3960 6780 9600 6790
rect 0 6770 1840 6780
rect 3400 6770 3680 6780
rect 3960 6770 9560 6780
rect 0 6760 1840 6770
rect 3400 6760 3680 6770
rect 3960 6760 9560 6770
rect 0 6750 1840 6760
rect 3400 6750 3680 6760
rect 3960 6750 9560 6760
rect 0 6740 1840 6750
rect 3400 6740 3680 6750
rect 3960 6740 9560 6750
rect 0 6730 1840 6740
rect 3400 6730 3760 6740
rect 3960 6730 9520 6740
rect 0 6720 1840 6730
rect 3400 6720 3760 6730
rect 3960 6720 9520 6730
rect 0 6710 1840 6720
rect 3400 6710 3760 6720
rect 3960 6710 9520 6720
rect 0 6700 1840 6710
rect 3400 6700 3760 6710
rect 3960 6700 9520 6710
rect 0 6690 1800 6700
rect 2280 6690 2480 6700
rect 3520 6690 3800 6700
rect 3960 6690 9520 6700
rect 0 6680 1800 6690
rect 2280 6680 2480 6690
rect 3520 6680 3800 6690
rect 3960 6680 9520 6690
rect 0 6670 1800 6680
rect 2280 6670 2480 6680
rect 3520 6670 3800 6680
rect 3960 6670 9520 6680
rect 0 6660 1800 6670
rect 2280 6660 2480 6670
rect 3520 6660 3800 6670
rect 3960 6660 9520 6670
rect 0 6650 1760 6660
rect 2240 6650 2520 6660
rect 3640 6650 3840 6660
rect 4000 6650 9480 6660
rect 9560 6650 9600 6660
rect 9880 6650 9990 6660
rect 0 6640 1760 6650
rect 2240 6640 2520 6650
rect 3640 6640 3840 6650
rect 4000 6640 9480 6650
rect 9560 6640 9600 6650
rect 9880 6640 9990 6650
rect 0 6630 1760 6640
rect 2240 6630 2520 6640
rect 3640 6630 3840 6640
rect 4000 6630 9480 6640
rect 9560 6630 9600 6640
rect 9880 6630 9990 6640
rect 0 6620 1760 6630
rect 2240 6620 2520 6630
rect 3640 6620 3840 6630
rect 4000 6620 9480 6630
rect 9560 6620 9600 6630
rect 9880 6620 9990 6630
rect 0 6610 1560 6620
rect 1680 6610 1760 6620
rect 2240 6610 2560 6620
rect 3720 6610 3880 6620
rect 4000 6610 9480 6620
rect 9760 6610 9990 6620
rect 0 6600 1560 6610
rect 1680 6600 1760 6610
rect 2240 6600 2560 6610
rect 3720 6600 3880 6610
rect 4000 6600 9480 6610
rect 9760 6600 9990 6610
rect 0 6590 1560 6600
rect 1680 6590 1760 6600
rect 2240 6590 2560 6600
rect 3720 6590 3880 6600
rect 4000 6590 9480 6600
rect 9760 6590 9990 6600
rect 0 6580 1560 6590
rect 1680 6580 1760 6590
rect 2240 6580 2560 6590
rect 3720 6580 3880 6590
rect 4000 6580 9480 6590
rect 9760 6580 9990 6590
rect 0 6570 1360 6580
rect 1400 6570 1480 6580
rect 2080 6570 2560 6580
rect 3800 6570 3920 6580
rect 4000 6570 6000 6580
rect 6480 6570 6560 6580
rect 6600 6570 9480 6580
rect 9520 6570 9990 6580
rect 0 6560 1360 6570
rect 1400 6560 1480 6570
rect 2080 6560 2560 6570
rect 3800 6560 3920 6570
rect 4000 6560 6000 6570
rect 6480 6560 6560 6570
rect 6600 6560 9480 6570
rect 9520 6560 9990 6570
rect 0 6550 1360 6560
rect 1400 6550 1480 6560
rect 2080 6550 2560 6560
rect 3800 6550 3920 6560
rect 4000 6550 6000 6560
rect 6480 6550 6560 6560
rect 6600 6550 9480 6560
rect 9520 6550 9990 6560
rect 0 6540 1360 6550
rect 1400 6540 1480 6550
rect 2080 6540 2560 6550
rect 3800 6540 3920 6550
rect 4000 6540 6000 6550
rect 6480 6540 6560 6550
rect 6600 6540 9480 6550
rect 9520 6540 9990 6550
rect 0 6530 1320 6540
rect 2080 6530 2240 6540
rect 2280 6530 2520 6540
rect 3880 6530 3960 6540
rect 4040 6530 5840 6540
rect 5880 6530 5960 6540
rect 6680 6530 9920 6540
rect 0 6520 1320 6530
rect 2080 6520 2240 6530
rect 2280 6520 2520 6530
rect 3880 6520 3960 6530
rect 4040 6520 5840 6530
rect 5880 6520 5960 6530
rect 6680 6520 9920 6530
rect 0 6510 1320 6520
rect 2080 6510 2240 6520
rect 2280 6510 2520 6520
rect 3880 6510 3960 6520
rect 4040 6510 5840 6520
rect 5880 6510 5960 6520
rect 6680 6510 9920 6520
rect 0 6500 1320 6510
rect 2080 6500 2240 6510
rect 2280 6500 2520 6510
rect 3880 6500 3960 6510
rect 4040 6500 5840 6510
rect 5880 6500 5960 6510
rect 6680 6500 9920 6510
rect 0 6490 1240 6500
rect 2160 6490 2240 6500
rect 2280 6490 2400 6500
rect 3920 6490 3960 6500
rect 4040 6490 5800 6500
rect 5880 6490 5960 6500
rect 6720 6490 9800 6500
rect 0 6480 1240 6490
rect 2160 6480 2240 6490
rect 2280 6480 2400 6490
rect 3920 6480 3960 6490
rect 4040 6480 5800 6490
rect 5880 6480 5960 6490
rect 6720 6480 9800 6490
rect 0 6470 1240 6480
rect 2160 6470 2240 6480
rect 2280 6470 2400 6480
rect 3920 6470 3960 6480
rect 4040 6470 5800 6480
rect 5880 6470 5960 6480
rect 6720 6470 9800 6480
rect 0 6460 1240 6470
rect 2160 6460 2240 6470
rect 2280 6460 2400 6470
rect 3920 6460 3960 6470
rect 4040 6460 5800 6470
rect 5880 6460 5960 6470
rect 6720 6460 9800 6470
rect 0 6450 1240 6460
rect 2160 6450 2280 6460
rect 2320 6450 2360 6460
rect 4000 6450 5720 6460
rect 6800 6450 9680 6460
rect 0 6440 1240 6450
rect 2160 6440 2280 6450
rect 2320 6440 2360 6450
rect 4000 6440 5720 6450
rect 6800 6440 9680 6450
rect 0 6430 1240 6440
rect 2160 6430 2280 6440
rect 2320 6430 2360 6440
rect 4000 6430 5720 6440
rect 6800 6430 9680 6440
rect 0 6420 1240 6430
rect 2160 6420 2280 6430
rect 2320 6420 2360 6430
rect 4000 6420 5720 6430
rect 6800 6420 9680 6430
rect 0 6410 1200 6420
rect 1640 6410 1720 6420
rect 2120 6410 2360 6420
rect 4040 6410 5680 6420
rect 6840 6410 9640 6420
rect 0 6400 1200 6410
rect 1640 6400 1720 6410
rect 2120 6400 2360 6410
rect 4040 6400 5680 6410
rect 6840 6400 9640 6410
rect 0 6390 1200 6400
rect 1640 6390 1720 6400
rect 2120 6390 2360 6400
rect 4040 6390 5680 6400
rect 6840 6390 9640 6400
rect 0 6380 1200 6390
rect 1640 6380 1720 6390
rect 2120 6380 2360 6390
rect 4040 6380 5680 6390
rect 6840 6380 9640 6390
rect 0 6370 1240 6380
rect 1280 6370 1400 6380
rect 1880 6370 1960 6380
rect 2040 6370 2400 6380
rect 4120 6370 5640 6380
rect 6280 6370 6320 6380
rect 6840 6370 9600 6380
rect 0 6360 1240 6370
rect 1280 6360 1400 6370
rect 1880 6360 1960 6370
rect 2040 6360 2400 6370
rect 4120 6360 5640 6370
rect 6280 6360 6320 6370
rect 6840 6360 9600 6370
rect 0 6350 1240 6360
rect 1280 6350 1400 6360
rect 1880 6350 1960 6360
rect 2040 6350 2400 6360
rect 4120 6350 5640 6360
rect 6280 6350 6320 6360
rect 6840 6350 9600 6360
rect 0 6340 1240 6350
rect 1280 6340 1400 6350
rect 1880 6340 1960 6350
rect 2040 6340 2400 6350
rect 4120 6340 5640 6350
rect 6280 6340 6320 6350
rect 6840 6340 9600 6350
rect 0 6330 1200 6340
rect 1320 6330 1400 6340
rect 1880 6330 2400 6340
rect 4160 6330 5400 6340
rect 5840 6330 6400 6340
rect 6840 6330 9320 6340
rect 9520 6330 9640 6340
rect 0 6320 1200 6330
rect 1320 6320 1400 6330
rect 1880 6320 2400 6330
rect 4160 6320 5400 6330
rect 5840 6320 6400 6330
rect 6840 6320 9320 6330
rect 9520 6320 9640 6330
rect 0 6310 1200 6320
rect 1320 6310 1400 6320
rect 1880 6310 2400 6320
rect 4160 6310 5400 6320
rect 5840 6310 6400 6320
rect 6840 6310 9320 6320
rect 9520 6310 9640 6320
rect 0 6300 1200 6310
rect 1320 6300 1400 6310
rect 1880 6300 2400 6310
rect 4160 6300 5400 6310
rect 5840 6300 6400 6310
rect 6840 6300 9320 6310
rect 9520 6300 9640 6310
rect 0 6290 1200 6300
rect 1320 6290 1400 6300
rect 1840 6290 2400 6300
rect 4200 6290 5360 6300
rect 5720 6290 6440 6300
rect 6840 6290 9280 6300
rect 9320 6290 9400 6300
rect 9440 6290 9480 6300
rect 9520 6290 9640 6300
rect 0 6280 1200 6290
rect 1320 6280 1400 6290
rect 1840 6280 2400 6290
rect 4200 6280 5360 6290
rect 5720 6280 6440 6290
rect 6840 6280 9280 6290
rect 9320 6280 9400 6290
rect 9440 6280 9480 6290
rect 9520 6280 9640 6290
rect 0 6270 1200 6280
rect 1320 6270 1400 6280
rect 1840 6270 2400 6280
rect 4200 6270 5360 6280
rect 5720 6270 6440 6280
rect 6840 6270 9280 6280
rect 9320 6270 9400 6280
rect 9440 6270 9480 6280
rect 9520 6270 9640 6280
rect 0 6260 1200 6270
rect 1320 6260 1400 6270
rect 1840 6260 2400 6270
rect 4200 6260 5360 6270
rect 5720 6260 6440 6270
rect 6840 6260 9280 6270
rect 9320 6260 9400 6270
rect 9440 6260 9480 6270
rect 9520 6260 9640 6270
rect 0 6250 1200 6260
rect 1800 6250 2400 6260
rect 4240 6250 5320 6260
rect 5640 6250 6520 6260
rect 6880 6250 9240 6260
rect 9320 6250 9400 6260
rect 9840 6250 9920 6260
rect 9960 6250 9990 6260
rect 0 6240 1200 6250
rect 1800 6240 2400 6250
rect 4240 6240 5320 6250
rect 5640 6240 6520 6250
rect 6880 6240 9240 6250
rect 9320 6240 9400 6250
rect 9840 6240 9920 6250
rect 9960 6240 9990 6250
rect 0 6230 1200 6240
rect 1800 6230 2400 6240
rect 4240 6230 5320 6240
rect 5640 6230 6520 6240
rect 6880 6230 9240 6240
rect 9320 6230 9400 6240
rect 9840 6230 9920 6240
rect 9960 6230 9990 6240
rect 0 6220 1200 6230
rect 1800 6220 2400 6230
rect 4240 6220 5320 6230
rect 5640 6220 6520 6230
rect 6880 6220 9240 6230
rect 9320 6220 9400 6230
rect 9840 6220 9920 6230
rect 9960 6220 9990 6230
rect 0 6210 1160 6220
rect 1800 6210 2400 6220
rect 4240 6210 5280 6220
rect 5560 6210 6560 6220
rect 6920 6210 9240 6220
rect 9640 6210 9680 6220
rect 9840 6210 9990 6220
rect 0 6200 1160 6210
rect 1800 6200 2400 6210
rect 4240 6200 5280 6210
rect 5560 6200 6560 6210
rect 6920 6200 9240 6210
rect 9640 6200 9680 6210
rect 9840 6200 9990 6210
rect 0 6190 1160 6200
rect 1800 6190 2400 6200
rect 4240 6190 5280 6200
rect 5560 6190 6560 6200
rect 6920 6190 9240 6200
rect 9640 6190 9680 6200
rect 9840 6190 9990 6200
rect 0 6180 1160 6190
rect 1800 6180 2400 6190
rect 4240 6180 5280 6190
rect 5560 6180 6560 6190
rect 6920 6180 9240 6190
rect 9640 6180 9680 6190
rect 9840 6180 9990 6190
rect 0 6170 1200 6180
rect 1800 6170 2400 6180
rect 4280 6170 5240 6180
rect 5480 6170 6640 6180
rect 6960 6170 9200 6180
rect 9840 6170 9990 6180
rect 0 6160 1200 6170
rect 1800 6160 2400 6170
rect 4280 6160 5240 6170
rect 5480 6160 6640 6170
rect 6960 6160 9200 6170
rect 9840 6160 9990 6170
rect 0 6150 1200 6160
rect 1800 6150 2400 6160
rect 4280 6150 5240 6160
rect 5480 6150 6640 6160
rect 6960 6150 9200 6160
rect 9840 6150 9990 6160
rect 0 6140 1200 6150
rect 1800 6140 2400 6150
rect 4280 6140 5240 6150
rect 5480 6140 6640 6150
rect 6960 6140 9200 6150
rect 9840 6140 9990 6150
rect 0 6130 1120 6140
rect 1160 6130 1200 6140
rect 1680 6130 1720 6140
rect 1800 6130 2440 6140
rect 4320 6130 5240 6140
rect 5440 6130 6640 6140
rect 7000 6130 9120 6140
rect 9960 6130 9990 6140
rect 0 6120 1120 6130
rect 1160 6120 1200 6130
rect 1680 6120 1720 6130
rect 1800 6120 2440 6130
rect 4320 6120 5240 6130
rect 5440 6120 6640 6130
rect 7000 6120 9120 6130
rect 9960 6120 9990 6130
rect 0 6110 1120 6120
rect 1160 6110 1200 6120
rect 1680 6110 1720 6120
rect 1800 6110 2440 6120
rect 4320 6110 5240 6120
rect 5440 6110 6640 6120
rect 7000 6110 9120 6120
rect 9960 6110 9990 6120
rect 0 6100 1120 6110
rect 1160 6100 1200 6110
rect 1680 6100 1720 6110
rect 1800 6100 2440 6110
rect 4320 6100 5240 6110
rect 5440 6100 6640 6110
rect 7000 6100 9120 6110
rect 9960 6100 9990 6110
rect 0 6090 1120 6100
rect 1800 6090 2440 6100
rect 3880 6090 3960 6100
rect 4320 6090 5200 6100
rect 5400 6090 6680 6100
rect 7000 6090 9000 6100
rect 9360 6090 9480 6100
rect 9960 6090 9990 6100
rect 0 6080 1120 6090
rect 1800 6080 2440 6090
rect 3880 6080 3960 6090
rect 4320 6080 5200 6090
rect 5400 6080 6680 6090
rect 7000 6080 9000 6090
rect 9360 6080 9480 6090
rect 9960 6080 9990 6090
rect 0 6070 1120 6080
rect 1800 6070 2440 6080
rect 3880 6070 3960 6080
rect 4320 6070 5200 6080
rect 5400 6070 6680 6080
rect 7000 6070 9000 6080
rect 9360 6070 9480 6080
rect 9960 6070 9990 6080
rect 0 6060 1120 6070
rect 1800 6060 2440 6070
rect 3880 6060 3960 6070
rect 4320 6060 5200 6070
rect 5400 6060 6680 6070
rect 7000 6060 9000 6070
rect 9360 6060 9480 6070
rect 9960 6060 9990 6070
rect 0 6050 800 6060
rect 960 6050 1040 6060
rect 1760 6050 2440 6060
rect 3800 6050 4000 6060
rect 4360 6050 5200 6060
rect 5400 6050 6720 6060
rect 7000 6050 8840 6060
rect 9240 6050 9280 6060
rect 9360 6050 9400 6060
rect 9440 6050 9480 6060
rect 9880 6050 9990 6060
rect 0 6040 800 6050
rect 960 6040 1040 6050
rect 1760 6040 2440 6050
rect 3800 6040 4000 6050
rect 4360 6040 5200 6050
rect 5400 6040 6720 6050
rect 7000 6040 8840 6050
rect 9240 6040 9280 6050
rect 9360 6040 9400 6050
rect 9440 6040 9480 6050
rect 9880 6040 9990 6050
rect 0 6030 800 6040
rect 960 6030 1040 6040
rect 1760 6030 2440 6040
rect 3800 6030 4000 6040
rect 4360 6030 5200 6040
rect 5400 6030 6720 6040
rect 7000 6030 8840 6040
rect 9240 6030 9280 6040
rect 9360 6030 9400 6040
rect 9440 6030 9480 6040
rect 9880 6030 9990 6040
rect 0 6020 800 6030
rect 960 6020 1040 6030
rect 1760 6020 2440 6030
rect 3800 6020 4000 6030
rect 4360 6020 5200 6030
rect 5400 6020 6720 6030
rect 7000 6020 8840 6030
rect 9240 6020 9280 6030
rect 9360 6020 9400 6030
rect 9440 6020 9480 6030
rect 9880 6020 9990 6030
rect 0 6010 760 6020
rect 1040 6010 1080 6020
rect 1800 6010 2480 6020
rect 3800 6010 4040 6020
rect 4360 6010 5160 6020
rect 5400 6010 6720 6020
rect 7000 6010 8720 6020
rect 9200 6010 9240 6020
rect 9360 6010 9440 6020
rect 9960 6010 9990 6020
rect 0 6000 760 6010
rect 1040 6000 1080 6010
rect 1800 6000 2480 6010
rect 3800 6000 4040 6010
rect 4360 6000 5160 6010
rect 5400 6000 6720 6010
rect 7000 6000 8720 6010
rect 9200 6000 9240 6010
rect 9360 6000 9440 6010
rect 9960 6000 9990 6010
rect 0 5990 760 6000
rect 1040 5990 1080 6000
rect 1800 5990 2480 6000
rect 3800 5990 4040 6000
rect 4360 5990 5160 6000
rect 5400 5990 6720 6000
rect 7000 5990 8720 6000
rect 9200 5990 9240 6000
rect 9360 5990 9440 6000
rect 9960 5990 9990 6000
rect 0 5980 760 5990
rect 1040 5980 1080 5990
rect 1800 5980 2480 5990
rect 3800 5980 4040 5990
rect 4360 5980 5160 5990
rect 5400 5980 6720 5990
rect 7000 5980 8720 5990
rect 9200 5980 9240 5990
rect 9360 5980 9440 5990
rect 9960 5980 9990 5990
rect 0 5970 720 5980
rect 1800 5970 2480 5980
rect 3800 5970 4080 5980
rect 4360 5970 5160 5980
rect 5360 5970 6720 5980
rect 7000 5970 8600 5980
rect 9040 5970 9120 5980
rect 9200 5970 9280 5980
rect 9360 5970 9400 5980
rect 9440 5970 9480 5980
rect 9960 5970 9990 5980
rect 0 5960 720 5970
rect 1800 5960 2480 5970
rect 3800 5960 4080 5970
rect 4360 5960 5160 5970
rect 5360 5960 6720 5970
rect 7000 5960 8600 5970
rect 9040 5960 9120 5970
rect 9200 5960 9280 5970
rect 9360 5960 9400 5970
rect 9440 5960 9480 5970
rect 9960 5960 9990 5970
rect 0 5950 720 5960
rect 1800 5950 2480 5960
rect 3800 5950 4080 5960
rect 4360 5950 5160 5960
rect 5360 5950 6720 5960
rect 7000 5950 8600 5960
rect 9040 5950 9120 5960
rect 9200 5950 9280 5960
rect 9360 5950 9400 5960
rect 9440 5950 9480 5960
rect 9960 5950 9990 5960
rect 0 5940 720 5950
rect 1800 5940 2480 5950
rect 3800 5940 4080 5950
rect 4360 5940 5160 5950
rect 5360 5940 6720 5950
rect 7000 5940 8600 5950
rect 9040 5940 9120 5950
rect 9200 5940 9280 5950
rect 9360 5940 9400 5950
rect 9440 5940 9480 5950
rect 9960 5940 9990 5950
rect 0 5930 680 5940
rect 840 5930 920 5940
rect 1760 5930 2440 5940
rect 3760 5930 3880 5940
rect 3920 5930 4160 5940
rect 4360 5930 5120 5940
rect 5360 5930 6760 5940
rect 7000 5930 8480 5940
rect 8840 5930 8920 5940
rect 9000 5930 9160 5940
rect 9200 5930 9240 5940
rect 9920 5930 9990 5940
rect 0 5920 680 5930
rect 840 5920 920 5930
rect 1760 5920 2440 5930
rect 3760 5920 3880 5930
rect 3920 5920 4160 5930
rect 4360 5920 5120 5930
rect 5360 5920 6760 5930
rect 7000 5920 8480 5930
rect 8840 5920 8920 5930
rect 9000 5920 9160 5930
rect 9200 5920 9240 5930
rect 9920 5920 9990 5930
rect 0 5910 680 5920
rect 840 5910 920 5920
rect 1760 5910 2440 5920
rect 3760 5910 3880 5920
rect 3920 5910 4160 5920
rect 4360 5910 5120 5920
rect 5360 5910 6760 5920
rect 7000 5910 8480 5920
rect 8840 5910 8920 5920
rect 9000 5910 9160 5920
rect 9200 5910 9240 5920
rect 9920 5910 9990 5920
rect 0 5900 680 5910
rect 840 5900 920 5910
rect 1760 5900 2440 5910
rect 3760 5900 3880 5910
rect 3920 5900 4160 5910
rect 4360 5900 5120 5910
rect 5360 5900 6760 5910
rect 7000 5900 8480 5910
rect 8840 5900 8920 5910
rect 9000 5900 9160 5910
rect 9200 5900 9240 5910
rect 9920 5900 9990 5910
rect 0 5890 640 5900
rect 840 5890 920 5900
rect 1880 5890 2320 5900
rect 3760 5890 5120 5900
rect 5360 5890 6760 5900
rect 7000 5890 8320 5900
rect 8800 5890 8840 5900
rect 8920 5890 8960 5900
rect 9000 5890 9160 5900
rect 9240 5890 9320 5900
rect 9920 5890 9990 5900
rect 0 5880 640 5890
rect 840 5880 920 5890
rect 1880 5880 2320 5890
rect 3760 5880 5120 5890
rect 5360 5880 6760 5890
rect 7000 5880 8320 5890
rect 8800 5880 8840 5890
rect 8920 5880 8960 5890
rect 9000 5880 9160 5890
rect 9240 5880 9320 5890
rect 9920 5880 9990 5890
rect 0 5870 640 5880
rect 840 5870 920 5880
rect 1880 5870 2320 5880
rect 3760 5870 5120 5880
rect 5360 5870 6760 5880
rect 7000 5870 8320 5880
rect 8800 5870 8840 5880
rect 8920 5870 8960 5880
rect 9000 5870 9160 5880
rect 9240 5870 9320 5880
rect 9920 5870 9990 5880
rect 0 5860 640 5870
rect 840 5860 920 5870
rect 1880 5860 2320 5870
rect 3760 5860 5120 5870
rect 5360 5860 6760 5870
rect 7000 5860 8320 5870
rect 8800 5860 8840 5870
rect 8920 5860 8960 5870
rect 9000 5860 9160 5870
rect 9240 5860 9320 5870
rect 9920 5860 9990 5870
rect 0 5850 560 5860
rect 1880 5850 2280 5860
rect 3880 5850 3920 5860
rect 3960 5850 5080 5860
rect 5360 5850 6760 5860
rect 7000 5850 8200 5860
rect 8680 5850 8720 5860
rect 8800 5850 8840 5860
rect 8920 5850 8960 5860
rect 9000 5850 9080 5860
rect 9120 5850 9160 5860
rect 9920 5850 9990 5860
rect 0 5840 560 5850
rect 1880 5840 2280 5850
rect 3880 5840 3920 5850
rect 3960 5840 5080 5850
rect 5360 5840 6760 5850
rect 7000 5840 8200 5850
rect 8680 5840 8720 5850
rect 8800 5840 8840 5850
rect 8920 5840 8960 5850
rect 9000 5840 9080 5850
rect 9120 5840 9160 5850
rect 9920 5840 9990 5850
rect 0 5830 560 5840
rect 1880 5830 2280 5840
rect 3880 5830 3920 5840
rect 3960 5830 5080 5840
rect 5360 5830 6760 5840
rect 7000 5830 8200 5840
rect 8680 5830 8720 5840
rect 8800 5830 8840 5840
rect 8920 5830 8960 5840
rect 9000 5830 9080 5840
rect 9120 5830 9160 5840
rect 9920 5830 9990 5840
rect 0 5820 560 5830
rect 1880 5820 2280 5830
rect 3880 5820 3920 5830
rect 3960 5820 5080 5830
rect 5360 5820 6760 5830
rect 7000 5820 8200 5830
rect 8680 5820 8720 5830
rect 8800 5820 8840 5830
rect 8920 5820 8960 5830
rect 9000 5820 9080 5830
rect 9120 5820 9160 5830
rect 9920 5820 9990 5830
rect 0 5810 560 5820
rect 760 5810 800 5820
rect 1920 5810 2240 5820
rect 2400 5810 2480 5820
rect 3120 5810 3160 5820
rect 3920 5810 5080 5820
rect 5360 5810 6800 5820
rect 7000 5810 8080 5820
rect 8680 5810 8720 5820
rect 8920 5810 8960 5820
rect 9960 5810 9990 5820
rect 0 5800 560 5810
rect 760 5800 800 5810
rect 1920 5800 2240 5810
rect 2400 5800 2480 5810
rect 3120 5800 3160 5810
rect 3920 5800 5080 5810
rect 5360 5800 6800 5810
rect 7000 5800 8080 5810
rect 8680 5800 8720 5810
rect 8920 5800 8960 5810
rect 9960 5800 9990 5810
rect 0 5790 560 5800
rect 760 5790 800 5800
rect 1920 5790 2240 5800
rect 2400 5790 2480 5800
rect 3120 5790 3160 5800
rect 3920 5790 5080 5800
rect 5360 5790 6800 5800
rect 7000 5790 8080 5800
rect 8680 5790 8720 5800
rect 8920 5790 8960 5800
rect 9960 5790 9990 5800
rect 0 5780 560 5790
rect 760 5780 800 5790
rect 1920 5780 2240 5790
rect 2400 5780 2480 5790
rect 3120 5780 3160 5790
rect 3920 5780 5080 5790
rect 5360 5780 6800 5790
rect 7000 5780 8080 5790
rect 8680 5780 8720 5790
rect 8920 5780 8960 5790
rect 9960 5780 9990 5790
rect 0 5770 560 5780
rect 720 5770 760 5780
rect 1960 5770 2200 5780
rect 3040 5770 3200 5780
rect 3920 5770 3960 5780
rect 4000 5770 5080 5780
rect 5320 5770 6800 5780
rect 7000 5770 7920 5780
rect 8840 5770 8920 5780
rect 9960 5770 9990 5780
rect 0 5760 560 5770
rect 720 5760 760 5770
rect 1960 5760 2200 5770
rect 3040 5760 3200 5770
rect 3920 5760 3960 5770
rect 4000 5760 5080 5770
rect 5320 5760 6800 5770
rect 7000 5760 7920 5770
rect 8840 5760 8920 5770
rect 9960 5760 9990 5770
rect 0 5750 560 5760
rect 720 5750 760 5760
rect 1960 5750 2200 5760
rect 3040 5750 3200 5760
rect 3920 5750 3960 5760
rect 4000 5750 5080 5760
rect 5320 5750 6800 5760
rect 7000 5750 7920 5760
rect 8840 5750 8920 5760
rect 9960 5750 9990 5760
rect 0 5740 560 5750
rect 720 5740 760 5750
rect 1960 5740 2200 5750
rect 3040 5740 3200 5750
rect 3920 5740 3960 5750
rect 4000 5740 5080 5750
rect 5320 5740 6800 5750
rect 7000 5740 7920 5750
rect 8840 5740 8920 5750
rect 9960 5740 9990 5750
rect 0 5730 600 5740
rect 680 5730 720 5740
rect 1960 5730 2200 5740
rect 3040 5730 3200 5740
rect 4000 5730 5080 5740
rect 5320 5730 6800 5740
rect 7000 5730 7760 5740
rect 8240 5730 8280 5740
rect 8400 5730 8440 5740
rect 9960 5730 9990 5740
rect 0 5720 600 5730
rect 680 5720 720 5730
rect 1960 5720 2200 5730
rect 3040 5720 3200 5730
rect 4000 5720 5080 5730
rect 5320 5720 6800 5730
rect 7000 5720 7760 5730
rect 8240 5720 8280 5730
rect 8400 5720 8440 5730
rect 9960 5720 9990 5730
rect 0 5710 600 5720
rect 680 5710 720 5720
rect 1960 5710 2200 5720
rect 3040 5710 3200 5720
rect 4000 5710 5080 5720
rect 5320 5710 6800 5720
rect 7000 5710 7760 5720
rect 8240 5710 8280 5720
rect 8400 5710 8440 5720
rect 9960 5710 9990 5720
rect 0 5700 600 5710
rect 680 5700 720 5710
rect 1960 5700 2200 5710
rect 3040 5700 3200 5710
rect 4000 5700 5080 5710
rect 5320 5700 6800 5710
rect 7000 5700 7760 5710
rect 8240 5700 8280 5710
rect 8400 5700 8440 5710
rect 9960 5700 9990 5710
rect 0 5690 800 5700
rect 1960 5690 2160 5700
rect 2840 5690 2920 5700
rect 3000 5690 3160 5700
rect 4000 5690 5080 5700
rect 5320 5690 6840 5700
rect 7000 5690 7680 5700
rect 8400 5690 8440 5700
rect 0 5680 800 5690
rect 1960 5680 2160 5690
rect 2840 5680 2920 5690
rect 3000 5680 3160 5690
rect 4000 5680 5080 5690
rect 5320 5680 6840 5690
rect 7000 5680 7680 5690
rect 8400 5680 8440 5690
rect 0 5670 800 5680
rect 1960 5670 2160 5680
rect 2840 5670 2920 5680
rect 3000 5670 3160 5680
rect 4000 5670 5080 5680
rect 5320 5670 6840 5680
rect 7000 5670 7680 5680
rect 8400 5670 8440 5680
rect 0 5660 800 5670
rect 1960 5660 2160 5670
rect 2840 5660 2920 5670
rect 3000 5660 3160 5670
rect 4000 5660 5080 5670
rect 5320 5660 6840 5670
rect 7000 5660 7680 5670
rect 8400 5660 8440 5670
rect 0 5650 520 5660
rect 640 5650 760 5660
rect 2000 5650 2160 5660
rect 2360 5650 2400 5660
rect 2840 5650 3160 5660
rect 3880 5650 3920 5660
rect 3960 5650 5080 5660
rect 5280 5650 5600 5660
rect 5800 5650 6840 5660
rect 7000 5650 7520 5660
rect 8040 5650 8080 5660
rect 8120 5650 8160 5660
rect 8440 5650 8520 5660
rect 0 5640 520 5650
rect 640 5640 760 5650
rect 2000 5640 2160 5650
rect 2360 5640 2400 5650
rect 2840 5640 3160 5650
rect 3880 5640 3920 5650
rect 3960 5640 5080 5650
rect 5280 5640 5600 5650
rect 5800 5640 6840 5650
rect 7000 5640 7520 5650
rect 8040 5640 8080 5650
rect 8120 5640 8160 5650
rect 8440 5640 8520 5650
rect 0 5630 520 5640
rect 640 5630 760 5640
rect 2000 5630 2160 5640
rect 2360 5630 2400 5640
rect 2840 5630 3160 5640
rect 3880 5630 3920 5640
rect 3960 5630 5080 5640
rect 5280 5630 5600 5640
rect 5800 5630 6840 5640
rect 7000 5630 7520 5640
rect 8040 5630 8080 5640
rect 8120 5630 8160 5640
rect 8440 5630 8520 5640
rect 0 5620 520 5630
rect 640 5620 760 5630
rect 2000 5620 2160 5630
rect 2360 5620 2400 5630
rect 2840 5620 3160 5630
rect 3880 5620 3920 5630
rect 3960 5620 5080 5630
rect 5280 5620 5600 5630
rect 5800 5620 6840 5630
rect 7000 5620 7520 5630
rect 8040 5620 8080 5630
rect 8120 5620 8160 5630
rect 8440 5620 8520 5630
rect 0 5610 520 5620
rect 2040 5610 2080 5620
rect 2360 5610 2400 5620
rect 2920 5610 3160 5620
rect 3800 5610 5080 5620
rect 5280 5610 5480 5620
rect 6080 5610 6160 5620
rect 6560 5610 6840 5620
rect 7000 5610 7400 5620
rect 7800 5610 7920 5620
rect 8040 5610 8160 5620
rect 8280 5610 8360 5620
rect 0 5600 520 5610
rect 2040 5600 2080 5610
rect 2360 5600 2400 5610
rect 2920 5600 3160 5610
rect 3800 5600 5080 5610
rect 5280 5600 5480 5610
rect 6080 5600 6160 5610
rect 6560 5600 6840 5610
rect 7000 5600 7400 5610
rect 7800 5600 7920 5610
rect 8040 5600 8160 5610
rect 8280 5600 8360 5610
rect 0 5590 520 5600
rect 2040 5590 2080 5600
rect 2360 5590 2400 5600
rect 2920 5590 3160 5600
rect 3800 5590 5080 5600
rect 5280 5590 5480 5600
rect 6080 5590 6160 5600
rect 6560 5590 6840 5600
rect 7000 5590 7400 5600
rect 7800 5590 7920 5600
rect 8040 5590 8160 5600
rect 8280 5590 8360 5600
rect 0 5580 520 5590
rect 2040 5580 2080 5590
rect 2360 5580 2400 5590
rect 2920 5580 3160 5590
rect 3800 5580 5080 5590
rect 5280 5580 5480 5590
rect 6080 5580 6160 5590
rect 6560 5580 6840 5590
rect 7000 5580 7400 5590
rect 7800 5580 7920 5590
rect 8040 5580 8160 5590
rect 8280 5580 8360 5590
rect 0 5570 520 5580
rect 3000 5570 3160 5580
rect 3800 5570 5080 5580
rect 5280 5570 5440 5580
rect 6640 5570 6880 5580
rect 6960 5570 7280 5580
rect 7320 5570 7360 5580
rect 7680 5570 7720 5580
rect 7800 5570 7840 5580
rect 7880 5570 7920 5580
rect 8040 5570 8080 5580
rect 8960 5570 9000 5580
rect 0 5560 520 5570
rect 3000 5560 3160 5570
rect 3800 5560 5080 5570
rect 5280 5560 5440 5570
rect 6640 5560 6880 5570
rect 6960 5560 7280 5570
rect 7320 5560 7360 5570
rect 7680 5560 7720 5570
rect 7800 5560 7840 5570
rect 7880 5560 7920 5570
rect 8040 5560 8080 5570
rect 8960 5560 9000 5570
rect 0 5550 520 5560
rect 3000 5550 3160 5560
rect 3800 5550 5080 5560
rect 5280 5550 5440 5560
rect 6640 5550 6880 5560
rect 6960 5550 7280 5560
rect 7320 5550 7360 5560
rect 7680 5550 7720 5560
rect 7800 5550 7840 5560
rect 7880 5550 7920 5560
rect 8040 5550 8080 5560
rect 8960 5550 9000 5560
rect 0 5540 520 5550
rect 3000 5540 3160 5550
rect 3800 5540 5080 5550
rect 5280 5540 5440 5550
rect 6640 5540 6880 5550
rect 6960 5540 7280 5550
rect 7320 5540 7360 5550
rect 7680 5540 7720 5550
rect 7800 5540 7840 5550
rect 7880 5540 7920 5550
rect 8040 5540 8080 5550
rect 8960 5540 9000 5550
rect 0 5530 440 5540
rect 3040 5530 3160 5540
rect 3760 5530 5080 5540
rect 5280 5530 5400 5540
rect 6040 5530 6120 5540
rect 6720 5530 6880 5540
rect 6960 5530 7280 5540
rect 7520 5530 7600 5540
rect 7800 5530 7840 5540
rect 7880 5530 7920 5540
rect 8760 5530 8800 5540
rect 8880 5530 8920 5540
rect 8960 5530 9000 5540
rect 0 5520 440 5530
rect 3040 5520 3160 5530
rect 3760 5520 5080 5530
rect 5280 5520 5400 5530
rect 6040 5520 6120 5530
rect 6720 5520 6880 5530
rect 6960 5520 7280 5530
rect 7520 5520 7600 5530
rect 7800 5520 7840 5530
rect 7880 5520 7920 5530
rect 8760 5520 8800 5530
rect 8880 5520 8920 5530
rect 8960 5520 9000 5530
rect 0 5510 440 5520
rect 3040 5510 3160 5520
rect 3760 5510 5080 5520
rect 5280 5510 5400 5520
rect 6040 5510 6120 5520
rect 6720 5510 6880 5520
rect 6960 5510 7280 5520
rect 7520 5510 7600 5520
rect 7800 5510 7840 5520
rect 7880 5510 7920 5520
rect 8760 5510 8800 5520
rect 8880 5510 8920 5520
rect 8960 5510 9000 5520
rect 0 5500 440 5510
rect 3040 5500 3160 5510
rect 3760 5500 5080 5510
rect 5280 5500 5400 5510
rect 6040 5500 6120 5510
rect 6720 5500 6880 5510
rect 6960 5500 7280 5510
rect 7520 5500 7600 5510
rect 7800 5500 7840 5510
rect 7880 5500 7920 5510
rect 8760 5500 8800 5510
rect 8880 5500 8920 5510
rect 8960 5500 9000 5510
rect 0 5490 400 5500
rect 3080 5490 3120 5500
rect 3680 5490 5080 5500
rect 5280 5490 5400 5500
rect 6000 5490 6120 5500
rect 6720 5490 6880 5500
rect 6960 5490 7240 5500
rect 7520 5490 7560 5500
rect 7680 5490 7720 5500
rect 7800 5490 7840 5500
rect 7880 5490 7920 5500
rect 8760 5490 8840 5500
rect 8880 5490 8920 5500
rect 8960 5490 9000 5500
rect 9080 5490 9120 5500
rect 0 5480 400 5490
rect 3080 5480 3120 5490
rect 3680 5480 5080 5490
rect 5280 5480 5400 5490
rect 6000 5480 6120 5490
rect 6720 5480 6880 5490
rect 6960 5480 7240 5490
rect 7520 5480 7560 5490
rect 7680 5480 7720 5490
rect 7800 5480 7840 5490
rect 7880 5480 7920 5490
rect 8760 5480 8840 5490
rect 8880 5480 8920 5490
rect 8960 5480 9000 5490
rect 9080 5480 9120 5490
rect 0 5470 400 5480
rect 3080 5470 3120 5480
rect 3680 5470 5080 5480
rect 5280 5470 5400 5480
rect 6000 5470 6120 5480
rect 6720 5470 6880 5480
rect 6960 5470 7240 5480
rect 7520 5470 7560 5480
rect 7680 5470 7720 5480
rect 7800 5470 7840 5480
rect 7880 5470 7920 5480
rect 8760 5470 8840 5480
rect 8880 5470 8920 5480
rect 8960 5470 9000 5480
rect 9080 5470 9120 5480
rect 0 5460 400 5470
rect 3080 5460 3120 5470
rect 3680 5460 5080 5470
rect 5280 5460 5400 5470
rect 6000 5460 6120 5470
rect 6720 5460 6880 5470
rect 6960 5460 7240 5470
rect 7520 5460 7560 5470
rect 7680 5460 7720 5470
rect 7800 5460 7840 5470
rect 7880 5460 7920 5470
rect 8760 5460 8840 5470
rect 8880 5460 8920 5470
rect 8960 5460 9000 5470
rect 9080 5460 9120 5470
rect 0 5450 440 5460
rect 520 5450 560 5460
rect 3600 5450 5080 5460
rect 5240 5450 5400 5460
rect 6000 5450 6120 5460
rect 6720 5450 6880 5460
rect 6960 5450 7200 5460
rect 7520 5450 7600 5460
rect 7680 5450 7720 5460
rect 7840 5450 7880 5460
rect 8520 5450 8560 5460
rect 8800 5450 8920 5460
rect 9080 5450 9120 5460
rect 0 5440 440 5450
rect 520 5440 560 5450
rect 3600 5440 5080 5450
rect 5240 5440 5400 5450
rect 6000 5440 6120 5450
rect 6720 5440 6880 5450
rect 6960 5440 7200 5450
rect 7520 5440 7600 5450
rect 7680 5440 7720 5450
rect 7840 5440 7880 5450
rect 8520 5440 8560 5450
rect 8800 5440 8920 5450
rect 9080 5440 9120 5450
rect 0 5430 440 5440
rect 520 5430 560 5440
rect 3600 5430 5080 5440
rect 5240 5430 5400 5440
rect 6000 5430 6120 5440
rect 6720 5430 6880 5440
rect 6960 5430 7200 5440
rect 7520 5430 7600 5440
rect 7680 5430 7720 5440
rect 7840 5430 7880 5440
rect 8520 5430 8560 5440
rect 8800 5430 8920 5440
rect 9080 5430 9120 5440
rect 0 5420 440 5430
rect 520 5420 560 5430
rect 3600 5420 5080 5430
rect 5240 5420 5400 5430
rect 6000 5420 6120 5430
rect 6720 5420 6880 5430
rect 6960 5420 7200 5430
rect 7520 5420 7600 5430
rect 7680 5420 7720 5430
rect 7840 5420 7880 5430
rect 8520 5420 8560 5430
rect 8800 5420 8920 5430
rect 9080 5420 9120 5430
rect 0 5410 400 5420
rect 520 5410 560 5420
rect 3600 5410 5080 5420
rect 5240 5410 5400 5420
rect 5960 5410 6120 5420
rect 6720 5410 6880 5420
rect 6960 5410 7240 5420
rect 7520 5410 7560 5420
rect 7600 5410 7640 5420
rect 8360 5410 8400 5420
rect 8440 5410 8480 5420
rect 8520 5410 8600 5420
rect 8640 5410 8680 5420
rect 8720 5410 8760 5420
rect 8800 5410 8840 5420
rect 8880 5410 8920 5420
rect 0 5400 400 5410
rect 520 5400 560 5410
rect 3600 5400 5080 5410
rect 5240 5400 5400 5410
rect 5960 5400 6120 5410
rect 6720 5400 6880 5410
rect 6960 5400 7240 5410
rect 7520 5400 7560 5410
rect 7600 5400 7640 5410
rect 8360 5400 8400 5410
rect 8440 5400 8480 5410
rect 8520 5400 8600 5410
rect 8640 5400 8680 5410
rect 8720 5400 8760 5410
rect 8800 5400 8840 5410
rect 8880 5400 8920 5410
rect 0 5390 400 5400
rect 520 5390 560 5400
rect 3600 5390 5080 5400
rect 5240 5390 5400 5400
rect 5960 5390 6120 5400
rect 6720 5390 6880 5400
rect 6960 5390 7240 5400
rect 7520 5390 7560 5400
rect 7600 5390 7640 5400
rect 8360 5390 8400 5400
rect 8440 5390 8480 5400
rect 8520 5390 8600 5400
rect 8640 5390 8680 5400
rect 8720 5390 8760 5400
rect 8800 5390 8840 5400
rect 8880 5390 8920 5400
rect 0 5380 400 5390
rect 520 5380 560 5390
rect 3600 5380 5080 5390
rect 5240 5380 5400 5390
rect 5960 5380 6120 5390
rect 6720 5380 6880 5390
rect 6960 5380 7240 5390
rect 7520 5380 7560 5390
rect 7600 5380 7640 5390
rect 8360 5380 8400 5390
rect 8440 5380 8480 5390
rect 8520 5380 8600 5390
rect 8640 5380 8680 5390
rect 8720 5380 8760 5390
rect 8800 5380 8840 5390
rect 8880 5380 8920 5390
rect 0 5370 280 5380
rect 3560 5370 5080 5380
rect 5240 5370 5360 5380
rect 5960 5370 6160 5380
rect 6760 5370 6920 5380
rect 6960 5370 7240 5380
rect 8240 5370 8280 5380
rect 8360 5370 8400 5380
rect 8440 5370 8480 5380
rect 8600 5370 8680 5380
rect 8720 5370 8760 5380
rect 8800 5370 8840 5380
rect 9520 5370 9560 5380
rect 0 5360 280 5370
rect 3560 5360 5080 5370
rect 5240 5360 5360 5370
rect 5960 5360 6160 5370
rect 6760 5360 6920 5370
rect 6960 5360 7240 5370
rect 8240 5360 8280 5370
rect 8360 5360 8400 5370
rect 8440 5360 8480 5370
rect 8600 5360 8680 5370
rect 8720 5360 8760 5370
rect 8800 5360 8840 5370
rect 9520 5360 9560 5370
rect 0 5350 280 5360
rect 3560 5350 5080 5360
rect 5240 5350 5360 5360
rect 5960 5350 6160 5360
rect 6760 5350 6920 5360
rect 6960 5350 7240 5360
rect 8240 5350 8280 5360
rect 8360 5350 8400 5360
rect 8440 5350 8480 5360
rect 8600 5350 8680 5360
rect 8720 5350 8760 5360
rect 8800 5350 8840 5360
rect 9520 5350 9560 5360
rect 0 5340 280 5350
rect 3560 5340 5080 5350
rect 5240 5340 5360 5350
rect 5960 5340 6160 5350
rect 6760 5340 6920 5350
rect 6960 5340 7240 5350
rect 8240 5340 8280 5350
rect 8360 5340 8400 5350
rect 8440 5340 8480 5350
rect 8600 5340 8680 5350
rect 8720 5340 8760 5350
rect 8800 5340 8840 5350
rect 9520 5340 9560 5350
rect 0 5330 240 5340
rect 3560 5330 5080 5340
rect 5240 5330 5640 5340
rect 5920 5330 6160 5340
rect 6800 5330 7240 5340
rect 8120 5330 8160 5340
rect 8240 5330 8280 5340
rect 8360 5330 8480 5340
rect 8640 5330 8680 5340
rect 9520 5330 9600 5340
rect 0 5320 240 5330
rect 3560 5320 5080 5330
rect 5240 5320 5640 5330
rect 5920 5320 6160 5330
rect 6800 5320 7240 5330
rect 8120 5320 8160 5330
rect 8240 5320 8280 5330
rect 8360 5320 8480 5330
rect 8640 5320 8680 5330
rect 9520 5320 9600 5330
rect 0 5310 240 5320
rect 3560 5310 5080 5320
rect 5240 5310 5640 5320
rect 5920 5310 6160 5320
rect 6800 5310 7240 5320
rect 8120 5310 8160 5320
rect 8240 5310 8280 5320
rect 8360 5310 8480 5320
rect 8640 5310 8680 5320
rect 9520 5310 9600 5320
rect 0 5300 240 5310
rect 3560 5300 5080 5310
rect 5240 5300 5640 5310
rect 5920 5300 6160 5310
rect 6800 5300 7240 5310
rect 8120 5300 8160 5310
rect 8240 5300 8280 5310
rect 8360 5300 8480 5310
rect 8640 5300 8680 5310
rect 9520 5300 9600 5310
rect 0 5290 200 5300
rect 3560 5290 5080 5300
rect 5240 5290 5560 5300
rect 5920 5290 6160 5300
rect 6800 5290 7240 5300
rect 8000 5290 8160 5300
rect 8240 5290 8320 5300
rect 9120 5290 9160 5300
rect 0 5280 200 5290
rect 3560 5280 5080 5290
rect 5240 5280 5560 5290
rect 5920 5280 6160 5290
rect 6800 5280 7240 5290
rect 8000 5280 8160 5290
rect 8240 5280 8320 5290
rect 9120 5280 9160 5290
rect 0 5270 200 5280
rect 3560 5270 5080 5280
rect 5240 5270 5560 5280
rect 5920 5270 6160 5280
rect 6800 5270 7240 5280
rect 8000 5270 8160 5280
rect 8240 5270 8320 5280
rect 9120 5270 9160 5280
rect 0 5260 200 5270
rect 3560 5260 5080 5270
rect 5240 5260 5560 5270
rect 5920 5260 6160 5270
rect 6800 5260 7240 5270
rect 8000 5260 8160 5270
rect 8240 5260 8320 5270
rect 9120 5260 9160 5270
rect 0 5250 160 5260
rect 3520 5250 5040 5260
rect 5240 5250 5560 5260
rect 5800 5250 6200 5260
rect 6600 5250 7240 5260
rect 8040 5250 8160 5260
rect 8240 5250 8320 5260
rect 9040 5250 9120 5260
rect 9760 5250 9800 5260
rect 9880 5250 9920 5260
rect 0 5240 160 5250
rect 3520 5240 5040 5250
rect 5240 5240 5560 5250
rect 5800 5240 6200 5250
rect 6600 5240 7240 5250
rect 8040 5240 8160 5250
rect 8240 5240 8320 5250
rect 9040 5240 9120 5250
rect 9760 5240 9800 5250
rect 9880 5240 9920 5250
rect 0 5230 160 5240
rect 3520 5230 5040 5240
rect 5240 5230 5560 5240
rect 5800 5230 6200 5240
rect 6600 5230 7240 5240
rect 8040 5230 8160 5240
rect 8240 5230 8320 5240
rect 9040 5230 9120 5240
rect 9760 5230 9800 5240
rect 9880 5230 9920 5240
rect 0 5220 160 5230
rect 3520 5220 5040 5230
rect 5240 5220 5560 5230
rect 5800 5220 6200 5230
rect 6600 5220 7240 5230
rect 8040 5220 8160 5230
rect 8240 5220 8320 5230
rect 9040 5220 9120 5230
rect 9760 5220 9800 5230
rect 9880 5220 9920 5230
rect 0 5210 80 5220
rect 2560 5210 2640 5220
rect 3520 5210 5040 5220
rect 5240 5210 6200 5220
rect 6280 5210 6360 5220
rect 6560 5210 7200 5220
rect 8040 5210 8080 5220
rect 8120 5210 8160 5220
rect 8840 5210 8880 5220
rect 8960 5210 9000 5220
rect 9120 5210 9160 5220
rect 9720 5210 9760 5220
rect 9800 5210 9840 5220
rect 0 5200 80 5210
rect 2560 5200 2640 5210
rect 3520 5200 5040 5210
rect 5240 5200 6200 5210
rect 6280 5200 6360 5210
rect 6560 5200 7200 5210
rect 8040 5200 8080 5210
rect 8120 5200 8160 5210
rect 8840 5200 8880 5210
rect 8960 5200 9000 5210
rect 9120 5200 9160 5210
rect 9720 5200 9760 5210
rect 9800 5200 9840 5210
rect 0 5190 80 5200
rect 2560 5190 2640 5200
rect 3520 5190 5040 5200
rect 5240 5190 6200 5200
rect 6280 5190 6360 5200
rect 6560 5190 7200 5200
rect 8040 5190 8080 5200
rect 8120 5190 8160 5200
rect 8840 5190 8880 5200
rect 8960 5190 9000 5200
rect 9120 5190 9160 5200
rect 9720 5190 9760 5200
rect 9800 5190 9840 5200
rect 0 5180 80 5190
rect 2560 5180 2640 5190
rect 3520 5180 5040 5190
rect 5240 5180 6200 5190
rect 6280 5180 6360 5190
rect 6560 5180 7200 5190
rect 8040 5180 8080 5190
rect 8120 5180 8160 5190
rect 8840 5180 8880 5190
rect 8960 5180 9000 5190
rect 9120 5180 9160 5190
rect 9720 5180 9760 5190
rect 9800 5180 9840 5190
rect 0 5170 40 5180
rect 2560 5170 2680 5180
rect 3480 5170 5080 5180
rect 5240 5170 7280 5180
rect 8040 5170 8080 5180
rect 8640 5170 8680 5180
rect 8760 5170 8800 5180
rect 8840 5170 8880 5180
rect 8960 5170 9040 5180
rect 9520 5170 9560 5180
rect 9720 5170 9760 5180
rect 0 5160 40 5170
rect 2560 5160 2680 5170
rect 3480 5160 5080 5170
rect 5240 5160 7280 5170
rect 8040 5160 8080 5170
rect 8640 5160 8680 5170
rect 8760 5160 8800 5170
rect 8840 5160 8880 5170
rect 8960 5160 9040 5170
rect 9520 5160 9560 5170
rect 9720 5160 9760 5170
rect 0 5150 40 5160
rect 2560 5150 2680 5160
rect 3480 5150 5080 5160
rect 5240 5150 7280 5160
rect 8040 5150 8080 5160
rect 8640 5150 8680 5160
rect 8760 5150 8800 5160
rect 8840 5150 8880 5160
rect 8960 5150 9040 5160
rect 9520 5150 9560 5160
rect 9720 5150 9760 5160
rect 0 5140 40 5150
rect 2560 5140 2680 5150
rect 3480 5140 5080 5150
rect 5240 5140 7280 5150
rect 8040 5140 8080 5150
rect 8640 5140 8680 5150
rect 8760 5140 8800 5150
rect 8840 5140 8880 5150
rect 8960 5140 9040 5150
rect 9520 5140 9560 5150
rect 9720 5140 9760 5150
rect 2560 5130 2640 5140
rect 3440 5130 5120 5140
rect 5240 5130 7280 5140
rect 9520 5130 9560 5140
rect 9600 5130 9640 5140
rect 9800 5130 9840 5140
rect 2560 5120 2640 5130
rect 3440 5120 5120 5130
rect 5240 5120 7280 5130
rect 9520 5120 9560 5130
rect 9600 5120 9640 5130
rect 9800 5120 9840 5130
rect 2560 5110 2640 5120
rect 3440 5110 5120 5120
rect 5240 5110 7280 5120
rect 9520 5110 9560 5120
rect 9600 5110 9640 5120
rect 9800 5110 9840 5120
rect 2560 5100 2640 5110
rect 3440 5100 5120 5110
rect 5240 5100 7280 5110
rect 9520 5100 9560 5110
rect 9600 5100 9640 5110
rect 9800 5100 9840 5110
rect 3440 5090 5120 5100
rect 5240 5090 7280 5100
rect 8320 5090 8360 5100
rect 9280 5090 9320 5100
rect 9400 5090 9440 5100
rect 9600 5090 9640 5100
rect 3440 5080 5120 5090
rect 5240 5080 7280 5090
rect 8320 5080 8360 5090
rect 9280 5080 9320 5090
rect 9400 5080 9440 5090
rect 9600 5080 9640 5090
rect 3440 5070 5120 5080
rect 5240 5070 7280 5080
rect 8320 5070 8360 5080
rect 9280 5070 9320 5080
rect 9400 5070 9440 5080
rect 9600 5070 9640 5080
rect 3440 5060 5120 5070
rect 5240 5060 7280 5070
rect 8320 5060 8360 5070
rect 9280 5060 9320 5070
rect 9400 5060 9440 5070
rect 9600 5060 9640 5070
rect 3400 5050 5160 5060
rect 5240 5050 5680 5060
rect 5800 5050 7280 5060
rect 8160 5050 8240 5060
rect 8280 5050 8320 5060
rect 8360 5050 8400 5060
rect 8440 5050 8480 5060
rect 9280 5050 9320 5060
rect 3400 5040 5160 5050
rect 5240 5040 5680 5050
rect 5800 5040 7280 5050
rect 8160 5040 8240 5050
rect 8280 5040 8320 5050
rect 8360 5040 8400 5050
rect 8440 5040 8480 5050
rect 9280 5040 9320 5050
rect 3400 5030 5160 5040
rect 5240 5030 5680 5040
rect 5800 5030 7280 5040
rect 8160 5030 8240 5040
rect 8280 5030 8320 5040
rect 8360 5030 8400 5040
rect 8440 5030 8480 5040
rect 9280 5030 9320 5040
rect 3400 5020 5160 5030
rect 5240 5020 5680 5030
rect 5800 5020 7280 5030
rect 8160 5020 8240 5030
rect 8280 5020 8320 5030
rect 8360 5020 8400 5030
rect 8440 5020 8480 5030
rect 9280 5020 9320 5030
rect 3400 5010 5160 5020
rect 5240 5010 5600 5020
rect 5800 5010 6320 5020
rect 6440 5010 7280 5020
rect 8080 5010 8120 5020
rect 8240 5010 8280 5020
rect 8320 5010 8360 5020
rect 8440 5010 8520 5020
rect 8880 5010 8920 5020
rect 8960 5010 9000 5020
rect 9040 5010 9080 5020
rect 3400 5000 5160 5010
rect 5240 5000 5600 5010
rect 5800 5000 6320 5010
rect 6440 5000 7280 5010
rect 8080 5000 8120 5010
rect 8240 5000 8280 5010
rect 8320 5000 8360 5010
rect 8440 5000 8520 5010
rect 8880 5000 8920 5010
rect 8960 5000 9000 5010
rect 9040 5000 9080 5010
rect 3400 4990 5160 5000
rect 5240 4990 5600 5000
rect 5800 4990 6320 5000
rect 6440 4990 7280 5000
rect 8080 4990 8120 5000
rect 8240 4990 8280 5000
rect 8320 4990 8360 5000
rect 8440 4990 8520 5000
rect 8880 4990 8920 5000
rect 8960 4990 9000 5000
rect 9040 4990 9080 5000
rect 3400 4980 5160 4990
rect 5240 4980 5600 4990
rect 5800 4980 6320 4990
rect 6440 4980 7280 4990
rect 8080 4980 8120 4990
rect 8240 4980 8280 4990
rect 8320 4980 8360 4990
rect 8440 4980 8520 4990
rect 8880 4980 8920 4990
rect 8960 4980 9000 4990
rect 9040 4980 9080 4990
rect 3400 4970 4000 4980
rect 4080 4970 4200 4980
rect 4440 4970 4640 4980
rect 4720 4970 5200 4980
rect 5240 4970 5520 4980
rect 5880 4970 5920 4980
rect 5960 4970 6040 4980
rect 6200 4970 6280 4980
rect 6560 4970 7320 4980
rect 8000 4970 8120 4980
rect 8160 4970 8200 4980
rect 8240 4970 8280 4980
rect 8920 4970 9000 4980
rect 9160 4970 9200 4980
rect 3400 4960 4000 4970
rect 4080 4960 4200 4970
rect 4440 4960 4640 4970
rect 4720 4960 5200 4970
rect 5240 4960 5520 4970
rect 5880 4960 5920 4970
rect 5960 4960 6040 4970
rect 6200 4960 6280 4970
rect 6560 4960 7320 4970
rect 8000 4960 8120 4970
rect 8160 4960 8200 4970
rect 8240 4960 8280 4970
rect 8920 4960 9000 4970
rect 9160 4960 9200 4970
rect 3400 4950 4000 4960
rect 4080 4950 4200 4960
rect 4440 4950 4640 4960
rect 4720 4950 5200 4960
rect 5240 4950 5520 4960
rect 5880 4950 5920 4960
rect 5960 4950 6040 4960
rect 6200 4950 6280 4960
rect 6560 4950 7320 4960
rect 8000 4950 8120 4960
rect 8160 4950 8200 4960
rect 8240 4950 8280 4960
rect 8920 4950 9000 4960
rect 9160 4950 9200 4960
rect 3400 4940 4000 4950
rect 4080 4940 4200 4950
rect 4440 4940 4640 4950
rect 4720 4940 5200 4950
rect 5240 4940 5520 4950
rect 5880 4940 5920 4950
rect 5960 4940 6040 4950
rect 6200 4940 6280 4950
rect 6560 4940 7320 4950
rect 8000 4940 8120 4950
rect 8160 4940 8200 4950
rect 8240 4940 8280 4950
rect 8920 4940 9000 4950
rect 9160 4940 9200 4950
rect 3400 4930 3960 4940
rect 4680 4930 4800 4940
rect 4840 4930 5200 4940
rect 5240 4930 5440 4940
rect 6680 4930 7320 4940
rect 7760 4930 7800 4940
rect 8040 4930 8120 4940
rect 8200 4930 8240 4940
rect 8600 4930 8640 4940
rect 8800 4930 8840 4940
rect 9160 4930 9280 4940
rect 3400 4920 3960 4930
rect 4680 4920 4800 4930
rect 4840 4920 5200 4930
rect 5240 4920 5440 4930
rect 6680 4920 7320 4930
rect 7760 4920 7800 4930
rect 8040 4920 8120 4930
rect 8200 4920 8240 4930
rect 8600 4920 8640 4930
rect 8800 4920 8840 4930
rect 9160 4920 9280 4930
rect 3400 4910 3960 4920
rect 4680 4910 4800 4920
rect 4840 4910 5200 4920
rect 5240 4910 5440 4920
rect 6680 4910 7320 4920
rect 7760 4910 7800 4920
rect 8040 4910 8120 4920
rect 8200 4910 8240 4920
rect 8600 4910 8640 4920
rect 8800 4910 8840 4920
rect 9160 4910 9280 4920
rect 3400 4900 3960 4910
rect 4680 4900 4800 4910
rect 4840 4900 5200 4910
rect 5240 4900 5440 4910
rect 6680 4900 7320 4910
rect 7760 4900 7800 4910
rect 8040 4900 8120 4910
rect 8200 4900 8240 4910
rect 8600 4900 8640 4910
rect 8800 4900 8840 4910
rect 9160 4900 9280 4910
rect 3400 4890 3680 4900
rect 3760 4890 3840 4900
rect 4920 4890 5200 4900
rect 5240 4890 5360 4900
rect 6720 4890 7320 4900
rect 7720 4890 7800 4900
rect 7840 4890 7880 4900
rect 7920 4890 7960 4900
rect 8480 4890 8520 4900
rect 8640 4890 8680 4900
rect 8760 4890 8800 4900
rect 9120 4890 9320 4900
rect 9480 4890 9520 4900
rect 9560 4890 9600 4900
rect 9640 4890 9680 4900
rect 3400 4880 3680 4890
rect 3760 4880 3840 4890
rect 4920 4880 5200 4890
rect 5240 4880 5360 4890
rect 6720 4880 7320 4890
rect 7720 4880 7800 4890
rect 7840 4880 7880 4890
rect 7920 4880 7960 4890
rect 8480 4880 8520 4890
rect 8640 4880 8680 4890
rect 8760 4880 8800 4890
rect 9120 4880 9320 4890
rect 9480 4880 9520 4890
rect 9560 4880 9600 4890
rect 9640 4880 9680 4890
rect 3400 4870 3680 4880
rect 3760 4870 3840 4880
rect 4920 4870 5200 4880
rect 5240 4870 5360 4880
rect 6720 4870 7320 4880
rect 7720 4870 7800 4880
rect 7840 4870 7880 4880
rect 7920 4870 7960 4880
rect 8480 4870 8520 4880
rect 8640 4870 8680 4880
rect 8760 4870 8800 4880
rect 9120 4870 9320 4880
rect 9480 4870 9520 4880
rect 9560 4870 9600 4880
rect 9640 4870 9680 4880
rect 3400 4860 3680 4870
rect 3760 4860 3840 4870
rect 4920 4860 5200 4870
rect 5240 4860 5360 4870
rect 6720 4860 7320 4870
rect 7720 4860 7800 4870
rect 7840 4860 7880 4870
rect 7920 4860 7960 4870
rect 8480 4860 8520 4870
rect 8640 4860 8680 4870
rect 8760 4860 8800 4870
rect 9120 4860 9320 4870
rect 9480 4860 9520 4870
rect 9560 4860 9600 4870
rect 9640 4860 9680 4870
rect 3400 4850 3640 4860
rect 5000 4850 5160 4860
rect 5240 4850 5360 4860
rect 6720 4850 7320 4860
rect 7720 4850 7800 4860
rect 7840 4850 7920 4860
rect 8280 4850 8360 4860
rect 8480 4850 8560 4860
rect 9080 4850 9320 4860
rect 9480 4850 9600 4860
rect 9640 4850 9680 4860
rect 3400 4840 3640 4850
rect 5000 4840 5160 4850
rect 5240 4840 5360 4850
rect 6720 4840 7320 4850
rect 7720 4840 7800 4850
rect 7840 4840 7920 4850
rect 8280 4840 8360 4850
rect 8480 4840 8560 4850
rect 9080 4840 9320 4850
rect 9480 4840 9600 4850
rect 9640 4840 9680 4850
rect 3400 4830 3640 4840
rect 5000 4830 5160 4840
rect 5240 4830 5360 4840
rect 6720 4830 7320 4840
rect 7720 4830 7800 4840
rect 7840 4830 7920 4840
rect 8280 4830 8360 4840
rect 8480 4830 8560 4840
rect 9080 4830 9320 4840
rect 9480 4830 9600 4840
rect 9640 4830 9680 4840
rect 3400 4820 3640 4830
rect 5000 4820 5160 4830
rect 5240 4820 5360 4830
rect 6720 4820 7320 4830
rect 7720 4820 7800 4830
rect 7840 4820 7920 4830
rect 8280 4820 8360 4830
rect 8480 4820 8560 4830
rect 9080 4820 9320 4830
rect 9480 4820 9600 4830
rect 9640 4820 9680 4830
rect 3400 4810 3600 4820
rect 5040 4810 5160 4820
rect 5240 4810 5360 4820
rect 6720 4810 7320 4820
rect 8120 4810 8160 4820
rect 8200 4810 8240 4820
rect 8280 4810 8320 4820
rect 9040 4810 9320 4820
rect 9480 4810 9520 4820
rect 3400 4800 3600 4810
rect 5040 4800 5160 4810
rect 5240 4800 5360 4810
rect 6720 4800 7320 4810
rect 8120 4800 8160 4810
rect 8200 4800 8240 4810
rect 8280 4800 8320 4810
rect 9040 4800 9320 4810
rect 9480 4800 9520 4810
rect 3400 4790 3600 4800
rect 5040 4790 5160 4800
rect 5240 4790 5360 4800
rect 6720 4790 7320 4800
rect 8120 4790 8160 4800
rect 8200 4790 8240 4800
rect 8280 4790 8320 4800
rect 9040 4790 9320 4800
rect 9480 4790 9520 4800
rect 3400 4780 3600 4790
rect 5040 4780 5160 4790
rect 5240 4780 5360 4790
rect 6720 4780 7320 4790
rect 8120 4780 8160 4790
rect 8200 4780 8240 4790
rect 8280 4780 8320 4790
rect 9040 4780 9320 4790
rect 9480 4780 9520 4790
rect 3360 4770 3520 4780
rect 5080 4770 5360 4780
rect 5760 4770 5920 4780
rect 6720 4770 7360 4780
rect 8000 4770 8080 4780
rect 8120 4770 8240 4780
rect 8360 4770 8400 4780
rect 8920 4770 8960 4780
rect 9000 4770 9280 4780
rect 3360 4760 3520 4770
rect 5080 4760 5360 4770
rect 5760 4760 5920 4770
rect 6720 4760 7360 4770
rect 8000 4760 8080 4770
rect 8120 4760 8240 4770
rect 8360 4760 8400 4770
rect 8920 4760 8960 4770
rect 9000 4760 9280 4770
rect 3360 4750 3520 4760
rect 5080 4750 5360 4760
rect 5760 4750 5920 4760
rect 6720 4750 7360 4760
rect 8000 4750 8080 4760
rect 8120 4750 8240 4760
rect 8360 4750 8400 4760
rect 8920 4750 8960 4760
rect 9000 4750 9280 4760
rect 3360 4740 3520 4750
rect 5080 4740 5360 4750
rect 5760 4740 5920 4750
rect 6720 4740 7360 4750
rect 8000 4740 8080 4750
rect 8120 4740 8240 4750
rect 8360 4740 8400 4750
rect 8920 4740 8960 4750
rect 9000 4740 9280 4750
rect 3360 4730 3480 4740
rect 5160 4730 5320 4740
rect 5760 4730 5920 4740
rect 6760 4730 7360 4740
rect 8000 4730 8040 4740
rect 8080 4730 8120 4740
rect 8200 4730 8240 4740
rect 8320 4730 8360 4740
rect 8920 4730 9280 4740
rect 9840 4730 9990 4740
rect 3360 4720 3480 4730
rect 5160 4720 5320 4730
rect 5760 4720 5920 4730
rect 6760 4720 7360 4730
rect 8000 4720 8040 4730
rect 8080 4720 8120 4730
rect 8200 4720 8240 4730
rect 8320 4720 8360 4730
rect 8920 4720 9280 4730
rect 9840 4720 9990 4730
rect 3360 4710 3480 4720
rect 5160 4710 5320 4720
rect 5760 4710 5920 4720
rect 6760 4710 7360 4720
rect 8000 4710 8040 4720
rect 8080 4710 8120 4720
rect 8200 4710 8240 4720
rect 8320 4710 8360 4720
rect 8920 4710 9280 4720
rect 9840 4710 9990 4720
rect 3360 4700 3480 4710
rect 5160 4700 5320 4710
rect 5760 4700 5920 4710
rect 6760 4700 7360 4710
rect 8000 4700 8040 4710
rect 8080 4700 8120 4710
rect 8200 4700 8240 4710
rect 8320 4700 8360 4710
rect 8920 4700 9280 4710
rect 9840 4700 9990 4710
rect 3400 4690 3480 4700
rect 5200 4690 5320 4700
rect 6760 4690 7360 4700
rect 7720 4690 7760 4700
rect 7800 4690 7840 4700
rect 7880 4690 7960 4700
rect 8000 4690 8040 4700
rect 8080 4690 8120 4700
rect 8600 4690 8640 4700
rect 9000 4690 9280 4700
rect 9840 4690 9990 4700
rect 3400 4680 3480 4690
rect 5200 4680 5320 4690
rect 6760 4680 7360 4690
rect 7720 4680 7760 4690
rect 7800 4680 7840 4690
rect 7880 4680 7960 4690
rect 8000 4680 8040 4690
rect 8080 4680 8120 4690
rect 8600 4680 8640 4690
rect 9000 4680 9280 4690
rect 9840 4680 9990 4690
rect 3400 4670 3480 4680
rect 5200 4670 5320 4680
rect 6760 4670 7360 4680
rect 7720 4670 7760 4680
rect 7800 4670 7840 4680
rect 7880 4670 7960 4680
rect 8000 4670 8040 4680
rect 8080 4670 8120 4680
rect 8600 4670 8640 4680
rect 9000 4670 9280 4680
rect 9840 4670 9990 4680
rect 3400 4660 3480 4670
rect 5200 4660 5320 4670
rect 6760 4660 7360 4670
rect 7720 4660 7760 4670
rect 7800 4660 7840 4670
rect 7880 4660 7960 4670
rect 8000 4660 8040 4670
rect 8080 4660 8120 4670
rect 8600 4660 8640 4670
rect 9000 4660 9280 4670
rect 9840 4660 9990 4670
rect 3400 4650 3440 4660
rect 5200 4650 5280 4660
rect 6760 4650 7360 4660
rect 7520 4650 7560 4660
rect 7600 4650 7640 4660
rect 7760 4650 7800 4660
rect 8520 4650 8560 4660
rect 8800 4650 8840 4660
rect 9000 4650 9240 4660
rect 9800 4650 9990 4660
rect 3400 4640 3440 4650
rect 5200 4640 5280 4650
rect 6760 4640 7360 4650
rect 7520 4640 7560 4650
rect 7600 4640 7640 4650
rect 7760 4640 7800 4650
rect 8520 4640 8560 4650
rect 8800 4640 8840 4650
rect 9000 4640 9240 4650
rect 9800 4640 9990 4650
rect 3400 4630 3440 4640
rect 5200 4630 5280 4640
rect 6760 4630 7360 4640
rect 7520 4630 7560 4640
rect 7600 4630 7640 4640
rect 7760 4630 7800 4640
rect 8520 4630 8560 4640
rect 8800 4630 8840 4640
rect 9000 4630 9240 4640
rect 9800 4630 9990 4640
rect 3400 4620 3440 4630
rect 5200 4620 5280 4630
rect 6760 4620 7360 4630
rect 7520 4620 7560 4630
rect 7600 4620 7640 4630
rect 7760 4620 7800 4630
rect 8520 4620 8560 4630
rect 8800 4620 8840 4630
rect 9000 4620 9240 4630
rect 9800 4620 9990 4630
rect 3400 4610 3440 4620
rect 5240 4610 5280 4620
rect 6720 4610 7360 4620
rect 7480 4610 7520 4620
rect 7760 4610 7840 4620
rect 8280 4610 8320 4620
rect 8520 4610 8560 4620
rect 9000 4610 9240 4620
rect 9760 4610 9990 4620
rect 3400 4600 3440 4610
rect 5240 4600 5280 4610
rect 6720 4600 7360 4610
rect 7480 4600 7520 4610
rect 7760 4600 7840 4610
rect 8280 4600 8320 4610
rect 8520 4600 8560 4610
rect 9000 4600 9240 4610
rect 9760 4600 9990 4610
rect 3400 4590 3440 4600
rect 5240 4590 5280 4600
rect 6720 4590 7360 4600
rect 7480 4590 7520 4600
rect 7760 4590 7840 4600
rect 8280 4590 8320 4600
rect 8520 4590 8560 4600
rect 9000 4590 9240 4600
rect 9760 4590 9990 4600
rect 3400 4580 3440 4590
rect 5240 4580 5280 4590
rect 6720 4580 7360 4590
rect 7480 4580 7520 4590
rect 7760 4580 7840 4590
rect 8280 4580 8320 4590
rect 8520 4580 8560 4590
rect 9000 4580 9240 4590
rect 9760 4580 9990 4590
rect 3280 4570 3320 4580
rect 3360 4570 3440 4580
rect 5240 4570 5280 4580
rect 5880 4570 6000 4580
rect 6720 4570 7320 4580
rect 7640 4570 7680 4580
rect 8160 4570 8200 4580
rect 8280 4570 8360 4580
rect 8520 4570 8600 4580
rect 8960 4570 9240 4580
rect 9720 4570 9960 4580
rect 3280 4560 3320 4570
rect 3360 4560 3440 4570
rect 5240 4560 5280 4570
rect 5880 4560 6000 4570
rect 6720 4560 7320 4570
rect 7640 4560 7680 4570
rect 8160 4560 8200 4570
rect 8280 4560 8360 4570
rect 8520 4560 8600 4570
rect 8960 4560 9240 4570
rect 9720 4560 9960 4570
rect 3280 4550 3320 4560
rect 3360 4550 3440 4560
rect 5240 4550 5280 4560
rect 5880 4550 6000 4560
rect 6720 4550 7320 4560
rect 7640 4550 7680 4560
rect 8160 4550 8200 4560
rect 8280 4550 8360 4560
rect 8520 4550 8600 4560
rect 8960 4550 9240 4560
rect 9720 4550 9960 4560
rect 3280 4540 3320 4550
rect 3360 4540 3440 4550
rect 5240 4540 5280 4550
rect 5880 4540 6000 4550
rect 6720 4540 7320 4550
rect 7640 4540 7680 4550
rect 8160 4540 8200 4550
rect 8280 4540 8360 4550
rect 8520 4540 8600 4550
rect 8960 4540 9240 4550
rect 9720 4540 9960 4550
rect 3280 4530 3400 4540
rect 5880 4530 6160 4540
rect 6720 4530 7320 4540
rect 7920 4530 7960 4540
rect 8040 4530 8120 4540
rect 8160 4530 8200 4540
rect 8320 4530 8400 4540
rect 8960 4530 9200 4540
rect 9680 4530 9960 4540
rect 3280 4520 3400 4530
rect 5880 4520 6160 4530
rect 6720 4520 7320 4530
rect 7920 4520 7960 4530
rect 8040 4520 8120 4530
rect 8160 4520 8200 4530
rect 8320 4520 8400 4530
rect 8960 4520 9200 4530
rect 9680 4520 9960 4530
rect 3280 4510 3400 4520
rect 5880 4510 6160 4520
rect 6720 4510 7320 4520
rect 7920 4510 7960 4520
rect 8040 4510 8120 4520
rect 8160 4510 8200 4520
rect 8320 4510 8400 4520
rect 8960 4510 9200 4520
rect 9680 4510 9960 4520
rect 3280 4500 3400 4510
rect 5880 4500 6160 4510
rect 6720 4500 7320 4510
rect 7920 4500 7960 4510
rect 8040 4500 8120 4510
rect 8160 4500 8200 4510
rect 8320 4500 8400 4510
rect 8960 4500 9200 4510
rect 9680 4500 9960 4510
rect 3280 4490 3400 4500
rect 5920 4490 6160 4500
rect 6720 4490 7320 4500
rect 7360 4490 7400 4500
rect 7760 4490 7840 4500
rect 7880 4490 7920 4500
rect 7960 4490 8000 4500
rect 8040 4490 8120 4500
rect 8920 4490 9200 4500
rect 9640 4490 9920 4500
rect 3280 4480 3400 4490
rect 5920 4480 6160 4490
rect 6720 4480 7320 4490
rect 7360 4480 7400 4490
rect 7760 4480 7840 4490
rect 7880 4480 7920 4490
rect 7960 4480 8000 4490
rect 8040 4480 8120 4490
rect 8920 4480 9200 4490
rect 9640 4480 9920 4490
rect 3280 4470 3400 4480
rect 5920 4470 6160 4480
rect 6720 4470 7320 4480
rect 7360 4470 7400 4480
rect 7760 4470 7840 4480
rect 7880 4470 7920 4480
rect 7960 4470 8000 4480
rect 8040 4470 8120 4480
rect 8920 4470 9200 4480
rect 9640 4470 9920 4480
rect 3280 4460 3400 4470
rect 5920 4460 6160 4470
rect 6720 4460 7320 4470
rect 7360 4460 7400 4470
rect 7760 4460 7840 4470
rect 7880 4460 7920 4470
rect 7960 4460 8000 4470
rect 8040 4460 8120 4470
rect 8920 4460 9200 4470
rect 9640 4460 9920 4470
rect 3320 4450 3360 4460
rect 6680 4450 7400 4460
rect 7800 4450 7840 4460
rect 7960 4450 8000 4460
rect 8040 4450 8080 4460
rect 8920 4450 9200 4460
rect 9600 4450 9840 4460
rect 3320 4440 3360 4450
rect 6680 4440 7400 4450
rect 7800 4440 7840 4450
rect 7960 4440 8000 4450
rect 8040 4440 8080 4450
rect 8920 4440 9200 4450
rect 9600 4440 9840 4450
rect 3320 4430 3360 4440
rect 6680 4430 7400 4440
rect 7800 4430 7840 4440
rect 7960 4430 8000 4440
rect 8040 4430 8080 4440
rect 8920 4430 9200 4440
rect 9600 4430 9840 4440
rect 3320 4420 3360 4430
rect 6680 4420 7400 4430
rect 7800 4420 7840 4430
rect 7960 4420 8000 4430
rect 8040 4420 8080 4430
rect 8920 4420 9200 4430
rect 9600 4420 9840 4430
rect 3000 4410 3040 4420
rect 3320 4410 3360 4420
rect 6680 4410 7320 4420
rect 7360 4410 7400 4420
rect 7920 4410 8000 4420
rect 8880 4410 9200 4420
rect 9560 4410 9840 4420
rect 3000 4400 3040 4410
rect 3320 4400 3360 4410
rect 6680 4400 7320 4410
rect 7360 4400 7400 4410
rect 7920 4400 8000 4410
rect 8880 4400 9200 4410
rect 9560 4400 9840 4410
rect 3000 4390 3040 4400
rect 3320 4390 3360 4400
rect 6680 4390 7320 4400
rect 7360 4390 7400 4400
rect 7920 4390 8000 4400
rect 8880 4390 9200 4400
rect 9560 4390 9840 4400
rect 3000 4380 3040 4390
rect 3320 4380 3360 4390
rect 6680 4380 7320 4390
rect 7360 4380 7400 4390
rect 7920 4380 8000 4390
rect 8880 4380 9200 4390
rect 9560 4380 9840 4390
rect 3000 4370 3040 4380
rect 5800 4370 5920 4380
rect 6680 4370 7320 4380
rect 8880 4370 9160 4380
rect 9520 4370 9840 4380
rect 3000 4360 3040 4370
rect 5800 4360 5920 4370
rect 6680 4360 7320 4370
rect 8880 4360 9160 4370
rect 9520 4360 9840 4370
rect 3000 4350 3040 4360
rect 5800 4350 5920 4360
rect 6680 4350 7320 4360
rect 8880 4350 9160 4360
rect 9520 4350 9840 4360
rect 3000 4340 3040 4350
rect 5800 4340 5920 4350
rect 6680 4340 7320 4350
rect 8880 4340 9160 4350
rect 9520 4340 9840 4350
rect 4680 4330 4760 4340
rect 5360 4330 5400 4340
rect 6680 4330 7280 4340
rect 8560 4330 8600 4340
rect 8880 4330 9160 4340
rect 9480 4330 9840 4340
rect 4680 4320 4760 4330
rect 5360 4320 5400 4330
rect 6680 4320 7280 4330
rect 8560 4320 8600 4330
rect 8880 4320 9160 4330
rect 9480 4320 9840 4330
rect 4680 4310 4760 4320
rect 5360 4310 5400 4320
rect 6680 4310 7280 4320
rect 8560 4310 8600 4320
rect 8880 4310 9160 4320
rect 9480 4310 9840 4320
rect 4680 4300 4760 4310
rect 5360 4300 5400 4310
rect 6680 4300 7280 4310
rect 8560 4300 8600 4310
rect 8880 4300 9160 4310
rect 9480 4300 9840 4310
rect 4640 4290 4840 4300
rect 5360 4290 5440 4300
rect 6640 4290 7120 4300
rect 8440 4290 8520 4300
rect 8880 4290 9160 4300
rect 9440 4290 9760 4300
rect 9960 4290 9990 4300
rect 4640 4280 4840 4290
rect 5360 4280 5440 4290
rect 6640 4280 7120 4290
rect 8440 4280 8520 4290
rect 8880 4280 9160 4290
rect 9440 4280 9760 4290
rect 9960 4280 9990 4290
rect 4640 4270 4840 4280
rect 5360 4270 5440 4280
rect 6640 4270 7120 4280
rect 8440 4270 8520 4280
rect 8880 4270 9160 4280
rect 9440 4270 9760 4280
rect 9960 4270 9990 4280
rect 4640 4260 4840 4270
rect 5360 4260 5440 4270
rect 6640 4260 7120 4270
rect 8440 4260 8520 4270
rect 8880 4260 9160 4270
rect 9440 4260 9760 4270
rect 9960 4260 9990 4270
rect 4600 4250 4840 4260
rect 5400 4250 5480 4260
rect 5640 4250 5720 4260
rect 6680 4250 7080 4260
rect 8840 4250 9160 4260
rect 9400 4250 9720 4260
rect 4600 4240 4840 4250
rect 5400 4240 5480 4250
rect 5640 4240 5720 4250
rect 6680 4240 7080 4250
rect 8840 4240 9160 4250
rect 9400 4240 9720 4250
rect 4600 4230 4840 4240
rect 5400 4230 5480 4240
rect 5640 4230 5720 4240
rect 6680 4230 7080 4240
rect 8840 4230 9160 4240
rect 9400 4230 9720 4240
rect 4600 4220 4840 4230
rect 5400 4220 5480 4230
rect 5640 4220 5720 4230
rect 6680 4220 7080 4230
rect 8840 4220 9160 4230
rect 9400 4220 9720 4230
rect 4240 4210 4320 4220
rect 5400 4210 5480 4220
rect 5640 4210 5920 4220
rect 6680 4210 7240 4220
rect 7360 4210 7440 4220
rect 8840 4210 9160 4220
rect 9320 4210 9680 4220
rect 9920 4210 9960 4220
rect 4240 4200 4320 4210
rect 5400 4200 5480 4210
rect 5640 4200 5920 4210
rect 6680 4200 7240 4210
rect 7360 4200 7440 4210
rect 8840 4200 9160 4210
rect 9320 4200 9680 4210
rect 9920 4200 9960 4210
rect 4240 4190 4320 4200
rect 5400 4190 5480 4200
rect 5640 4190 5920 4200
rect 6680 4190 7240 4200
rect 7360 4190 7440 4200
rect 8840 4190 9160 4200
rect 9320 4190 9680 4200
rect 9920 4190 9960 4200
rect 4240 4180 4320 4190
rect 5400 4180 5480 4190
rect 5640 4180 5920 4190
rect 6680 4180 7240 4190
rect 7360 4180 7440 4190
rect 8840 4180 9160 4190
rect 9320 4180 9680 4190
rect 9920 4180 9960 4190
rect 4200 4170 4360 4180
rect 5440 4170 5480 4180
rect 5680 4170 5920 4180
rect 6680 4170 7240 4180
rect 7360 4170 7440 4180
rect 8840 4170 9280 4180
rect 9320 4170 9640 4180
rect 9680 4170 9800 4180
rect 9920 4170 9960 4180
rect 4200 4160 4360 4170
rect 5440 4160 5480 4170
rect 5680 4160 5920 4170
rect 6680 4160 7240 4170
rect 7360 4160 7440 4170
rect 8840 4160 9280 4170
rect 9320 4160 9640 4170
rect 9680 4160 9800 4170
rect 9920 4160 9960 4170
rect 4200 4150 4360 4160
rect 5440 4150 5480 4160
rect 5680 4150 5920 4160
rect 6680 4150 7240 4160
rect 7360 4150 7440 4160
rect 8840 4150 9280 4160
rect 9320 4150 9640 4160
rect 9680 4150 9800 4160
rect 9920 4150 9960 4160
rect 4200 4140 4360 4150
rect 5440 4140 5480 4150
rect 5680 4140 5920 4150
rect 6680 4140 7240 4150
rect 7360 4140 7440 4150
rect 8840 4140 9280 4150
rect 9320 4140 9640 4150
rect 9680 4140 9800 4150
rect 9920 4140 9960 4150
rect 4160 4130 4400 4140
rect 5720 4130 5960 4140
rect 6680 4130 7240 4140
rect 8800 4130 9800 4140
rect 4160 4120 4400 4130
rect 5720 4120 5960 4130
rect 6680 4120 7240 4130
rect 8800 4120 9800 4130
rect 4160 4110 4400 4120
rect 5720 4110 5960 4120
rect 6680 4110 7240 4120
rect 8800 4110 9800 4120
rect 4160 4100 4400 4110
rect 5720 4100 5960 4110
rect 6680 4100 7240 4110
rect 8800 4100 9800 4110
rect 4120 4090 4440 4100
rect 4920 4090 5040 4100
rect 5440 4090 5480 4100
rect 5840 4090 5960 4100
rect 6640 4090 7200 4100
rect 8800 4090 9600 4100
rect 9760 4090 9880 4100
rect 4120 4080 4440 4090
rect 4920 4080 5040 4090
rect 5440 4080 5480 4090
rect 5840 4080 5960 4090
rect 6640 4080 7200 4090
rect 8800 4080 9600 4090
rect 9760 4080 9880 4090
rect 4120 4070 4440 4080
rect 4920 4070 5040 4080
rect 5440 4070 5480 4080
rect 5840 4070 5960 4080
rect 6640 4070 7200 4080
rect 8800 4070 9600 4080
rect 9760 4070 9880 4080
rect 4120 4060 4440 4070
rect 4920 4060 5040 4070
rect 5440 4060 5480 4070
rect 5840 4060 5960 4070
rect 6640 4060 7200 4070
rect 8800 4060 9600 4070
rect 9760 4060 9880 4070
rect 4080 4050 4160 4060
rect 4280 4050 4480 4060
rect 4800 4050 4840 4060
rect 4920 4050 5040 4060
rect 5440 4050 5480 4060
rect 6640 4050 7200 4060
rect 8800 4050 9990 4060
rect 4080 4040 4160 4050
rect 4280 4040 4480 4050
rect 4800 4040 4840 4050
rect 4920 4040 5040 4050
rect 5440 4040 5480 4050
rect 6640 4040 7200 4050
rect 8800 4040 9990 4050
rect 4080 4030 4160 4040
rect 4280 4030 4480 4040
rect 4800 4030 4840 4040
rect 4920 4030 5040 4040
rect 5440 4030 5480 4040
rect 6640 4030 7200 4040
rect 8800 4030 9990 4040
rect 4080 4020 4160 4030
rect 4280 4020 4480 4030
rect 4800 4020 4840 4030
rect 4920 4020 5040 4030
rect 5440 4020 5480 4030
rect 6640 4020 7200 4030
rect 8800 4020 9990 4030
rect 4080 4010 4160 4020
rect 4320 4010 4520 4020
rect 4880 4010 5040 4020
rect 5440 4010 5480 4020
rect 6600 4010 7120 4020
rect 8760 4010 9990 4020
rect 4080 4000 4160 4010
rect 4320 4000 4520 4010
rect 4880 4000 5040 4010
rect 5440 4000 5480 4010
rect 6600 4000 7120 4010
rect 8760 4000 9990 4010
rect 4080 3990 4160 4000
rect 4320 3990 4520 4000
rect 4880 3990 5040 4000
rect 5440 3990 5480 4000
rect 6600 3990 7120 4000
rect 8760 3990 9990 4000
rect 4080 3980 4160 3990
rect 4320 3980 4520 3990
rect 4880 3980 5040 3990
rect 5440 3980 5480 3990
rect 6600 3980 7120 3990
rect 8760 3980 9990 3990
rect 4040 3970 4120 3980
rect 4360 3970 4520 3980
rect 4840 3970 5120 3980
rect 6600 3970 7120 3980
rect 8360 3970 8400 3980
rect 8600 3970 8640 3980
rect 8760 3970 9680 3980
rect 9720 3970 9990 3980
rect 4040 3960 4120 3970
rect 4360 3960 4520 3970
rect 4840 3960 5120 3970
rect 6600 3960 7120 3970
rect 8360 3960 8400 3970
rect 8600 3960 8640 3970
rect 8760 3960 9680 3970
rect 9720 3960 9990 3970
rect 4040 3950 4120 3960
rect 4360 3950 4520 3960
rect 4840 3950 5120 3960
rect 6600 3950 7120 3960
rect 8360 3950 8400 3960
rect 8600 3950 8640 3960
rect 8760 3950 9680 3960
rect 9720 3950 9990 3960
rect 4040 3940 4120 3950
rect 4360 3940 4520 3950
rect 4840 3940 5120 3950
rect 6600 3940 7120 3950
rect 8360 3940 8400 3950
rect 8600 3940 8640 3950
rect 8760 3940 9680 3950
rect 9720 3940 9990 3950
rect 3960 3930 4080 3940
rect 4360 3930 4520 3940
rect 4720 3930 5120 3940
rect 6600 3930 7120 3940
rect 8200 3930 8240 3940
rect 8320 3930 8440 3940
rect 8720 3930 9600 3940
rect 9760 3930 9990 3940
rect 3960 3920 4080 3930
rect 4360 3920 4520 3930
rect 4720 3920 5120 3930
rect 6600 3920 7120 3930
rect 8200 3920 8240 3930
rect 8320 3920 8440 3930
rect 8720 3920 9600 3930
rect 9760 3920 9990 3930
rect 3960 3910 4080 3920
rect 4360 3910 4520 3920
rect 4720 3910 5120 3920
rect 6600 3910 7120 3920
rect 8200 3910 8240 3920
rect 8320 3910 8440 3920
rect 8720 3910 9600 3920
rect 9760 3910 9990 3920
rect 3960 3900 4080 3910
rect 4360 3900 4520 3910
rect 4720 3900 5120 3910
rect 6600 3900 7120 3910
rect 8200 3900 8240 3910
rect 8320 3900 8440 3910
rect 8720 3900 9600 3910
rect 9760 3900 9990 3910
rect 3200 3890 3280 3900
rect 3960 3890 4000 3900
rect 4400 3890 4560 3900
rect 4640 3890 5160 3900
rect 6600 3890 7120 3900
rect 8240 3890 8280 3900
rect 8360 3890 8400 3900
rect 8480 3890 8520 3900
rect 8720 3890 9440 3900
rect 9840 3890 9990 3900
rect 3200 3880 3280 3890
rect 3960 3880 4000 3890
rect 4400 3880 4560 3890
rect 4640 3880 5160 3890
rect 6600 3880 7120 3890
rect 8240 3880 8280 3890
rect 8360 3880 8400 3890
rect 8480 3880 8520 3890
rect 8720 3880 9440 3890
rect 9840 3880 9990 3890
rect 3200 3870 3280 3880
rect 3960 3870 4000 3880
rect 4400 3870 4560 3880
rect 4640 3870 5160 3880
rect 6600 3870 7120 3880
rect 8240 3870 8280 3880
rect 8360 3870 8400 3880
rect 8480 3870 8520 3880
rect 8720 3870 9440 3880
rect 9840 3870 9990 3880
rect 3200 3860 3280 3870
rect 3960 3860 4000 3870
rect 4400 3860 4560 3870
rect 4640 3860 5160 3870
rect 6600 3860 7120 3870
rect 8240 3860 8280 3870
rect 8360 3860 8400 3870
rect 8480 3860 8520 3870
rect 8720 3860 9440 3870
rect 9840 3860 9990 3870
rect 3200 3850 3240 3860
rect 3920 3850 3960 3860
rect 4400 3850 4600 3860
rect 4640 3850 5160 3860
rect 6600 3850 7080 3860
rect 8280 3850 8320 3860
rect 8480 3850 8560 3860
rect 8680 3850 9560 3860
rect 9880 3850 9990 3860
rect 3200 3840 3240 3850
rect 3920 3840 3960 3850
rect 4400 3840 4600 3850
rect 4640 3840 5160 3850
rect 6600 3840 7080 3850
rect 8280 3840 8320 3850
rect 8480 3840 8560 3850
rect 8680 3840 9560 3850
rect 9880 3840 9990 3850
rect 3200 3830 3240 3840
rect 3920 3830 3960 3840
rect 4400 3830 4600 3840
rect 4640 3830 5160 3840
rect 6600 3830 7080 3840
rect 8280 3830 8320 3840
rect 8480 3830 8560 3840
rect 8680 3830 9560 3840
rect 9880 3830 9990 3840
rect 3200 3820 3240 3830
rect 3920 3820 3960 3830
rect 4400 3820 4600 3830
rect 4640 3820 5160 3830
rect 6600 3820 7080 3830
rect 8280 3820 8320 3830
rect 8480 3820 8560 3830
rect 8680 3820 9560 3830
rect 9880 3820 9990 3830
rect 3200 3810 3240 3820
rect 4440 3810 5160 3820
rect 6600 3810 7080 3820
rect 8520 3810 8640 3820
rect 8680 3810 9600 3820
rect 9880 3810 9990 3820
rect 3200 3800 3240 3810
rect 4440 3800 5160 3810
rect 6600 3800 7080 3810
rect 8520 3800 8640 3810
rect 8680 3800 9600 3810
rect 9880 3800 9990 3810
rect 3200 3790 3240 3800
rect 4440 3790 5160 3800
rect 6600 3790 7080 3800
rect 8520 3790 8640 3800
rect 8680 3790 9600 3800
rect 9880 3790 9990 3800
rect 3200 3780 3240 3790
rect 4440 3780 5160 3790
rect 6600 3780 7080 3790
rect 8520 3780 8640 3790
rect 8680 3780 9600 3790
rect 9880 3780 9990 3790
rect 4440 3770 4840 3780
rect 4920 3770 5160 3780
rect 6600 3770 7040 3780
rect 8400 3770 8480 3780
rect 8560 3770 9640 3780
rect 9880 3770 9990 3780
rect 4440 3760 4840 3770
rect 4920 3760 5160 3770
rect 6600 3760 7040 3770
rect 8400 3760 8480 3770
rect 8560 3760 9640 3770
rect 9880 3760 9990 3770
rect 4440 3750 4840 3760
rect 4920 3750 5160 3760
rect 6600 3750 7040 3760
rect 8400 3750 8480 3760
rect 8560 3750 9640 3760
rect 9880 3750 9990 3760
rect 4440 3740 4840 3750
rect 4920 3740 5160 3750
rect 6600 3740 7040 3750
rect 8400 3740 8480 3750
rect 8560 3740 9640 3750
rect 9880 3740 9990 3750
rect 4080 3730 4120 3740
rect 4440 3730 4800 3740
rect 6600 3730 7000 3740
rect 8440 3730 8520 3740
rect 8600 3730 9680 3740
rect 4080 3720 4120 3730
rect 4440 3720 4800 3730
rect 6600 3720 7000 3730
rect 8440 3720 8520 3730
rect 8600 3720 9680 3730
rect 4080 3710 4120 3720
rect 4440 3710 4800 3720
rect 6600 3710 7000 3720
rect 8440 3710 8520 3720
rect 8600 3710 9680 3720
rect 4080 3700 4120 3710
rect 4440 3700 4800 3710
rect 6600 3700 7000 3710
rect 8440 3700 8520 3710
rect 8600 3700 9680 3710
rect 4240 3690 4320 3700
rect 4440 3690 4800 3700
rect 6600 3690 6960 3700
rect 8240 3690 8360 3700
rect 8520 3690 8560 3700
rect 8640 3690 9560 3700
rect 9640 3690 9840 3700
rect 9960 3690 9990 3700
rect 4240 3680 4320 3690
rect 4440 3680 4800 3690
rect 6600 3680 6960 3690
rect 8240 3680 8360 3690
rect 8520 3680 8560 3690
rect 8640 3680 9560 3690
rect 9640 3680 9840 3690
rect 9960 3680 9990 3690
rect 4240 3670 4320 3680
rect 4440 3670 4800 3680
rect 6600 3670 6960 3680
rect 8240 3670 8360 3680
rect 8520 3670 8560 3680
rect 8640 3670 9560 3680
rect 9640 3670 9840 3680
rect 9960 3670 9990 3680
rect 4240 3660 4320 3670
rect 4440 3660 4800 3670
rect 6600 3660 6960 3670
rect 8240 3660 8360 3670
rect 8520 3660 8560 3670
rect 8640 3660 9560 3670
rect 9640 3660 9840 3670
rect 9960 3660 9990 3670
rect 4040 3650 4320 3660
rect 4440 3650 4800 3660
rect 6600 3650 6960 3660
rect 8240 3650 8360 3660
rect 8560 3650 9520 3660
rect 9680 3650 9840 3660
rect 9920 3650 9990 3660
rect 4040 3640 4320 3650
rect 4440 3640 4800 3650
rect 6600 3640 6960 3650
rect 8240 3640 8360 3650
rect 8560 3640 9520 3650
rect 9680 3640 9840 3650
rect 9920 3640 9990 3650
rect 4040 3630 4320 3640
rect 4440 3630 4800 3640
rect 6600 3630 6960 3640
rect 8240 3630 8360 3640
rect 8560 3630 9520 3640
rect 9680 3630 9840 3640
rect 9920 3630 9990 3640
rect 4040 3620 4320 3630
rect 4440 3620 4800 3630
rect 6600 3620 6960 3630
rect 8240 3620 8360 3630
rect 8560 3620 9520 3630
rect 9680 3620 9840 3630
rect 9920 3620 9990 3630
rect 4040 3610 4320 3620
rect 4440 3610 4760 3620
rect 4840 3610 4880 3620
rect 6600 3610 6920 3620
rect 8280 3610 8360 3620
rect 8520 3610 9440 3620
rect 9680 3610 9990 3620
rect 4040 3600 4320 3610
rect 4440 3600 4760 3610
rect 4840 3600 4880 3610
rect 6600 3600 6920 3610
rect 8280 3600 8360 3610
rect 8520 3600 9440 3610
rect 9680 3600 9990 3610
rect 4040 3590 4320 3600
rect 4440 3590 4760 3600
rect 4840 3590 4880 3600
rect 6600 3590 6920 3600
rect 8280 3590 8360 3600
rect 8520 3590 9440 3600
rect 9680 3590 9990 3600
rect 4040 3580 4320 3590
rect 4440 3580 4760 3590
rect 4840 3580 4880 3590
rect 6600 3580 6920 3590
rect 8280 3580 8360 3590
rect 8520 3580 9440 3590
rect 9680 3580 9990 3590
rect 4040 3570 4280 3580
rect 4480 3570 4680 3580
rect 4840 3570 5000 3580
rect 6600 3570 6880 3580
rect 8320 3570 8360 3580
rect 8520 3570 9240 3580
rect 9520 3570 9640 3580
rect 9680 3570 9990 3580
rect 4040 3560 4280 3570
rect 4480 3560 4680 3570
rect 4840 3560 5000 3570
rect 6600 3560 6880 3570
rect 8320 3560 8360 3570
rect 8520 3560 9240 3570
rect 9520 3560 9640 3570
rect 9680 3560 9990 3570
rect 4040 3550 4280 3560
rect 4480 3550 4680 3560
rect 4840 3550 5000 3560
rect 6600 3550 6880 3560
rect 8320 3550 8360 3560
rect 8520 3550 9240 3560
rect 9520 3550 9640 3560
rect 9680 3550 9990 3560
rect 4040 3540 4280 3550
rect 4480 3540 4680 3550
rect 4840 3540 5000 3550
rect 6600 3540 6880 3550
rect 8320 3540 8360 3550
rect 8520 3540 9240 3550
rect 9520 3540 9640 3550
rect 9680 3540 9990 3550
rect 4040 3530 4240 3540
rect 4520 3530 4600 3540
rect 4840 3530 5000 3540
rect 6560 3530 6840 3540
rect 8520 3530 9160 3540
rect 9480 3530 9600 3540
rect 9680 3530 9990 3540
rect 4040 3520 4240 3530
rect 4520 3520 4600 3530
rect 4840 3520 5000 3530
rect 6560 3520 6840 3530
rect 8520 3520 9160 3530
rect 9480 3520 9600 3530
rect 9680 3520 9990 3530
rect 4040 3510 4240 3520
rect 4520 3510 4600 3520
rect 4840 3510 5000 3520
rect 6560 3510 6840 3520
rect 8520 3510 9160 3520
rect 9480 3510 9600 3520
rect 9680 3510 9990 3520
rect 4040 3500 4240 3510
rect 4520 3500 4600 3510
rect 4840 3500 5000 3510
rect 6560 3500 6840 3510
rect 8520 3500 9160 3510
rect 9480 3500 9600 3510
rect 9680 3500 9990 3510
rect 2480 3490 2600 3500
rect 4080 3490 4200 3500
rect 4800 3490 4920 3500
rect 6560 3490 6800 3500
rect 8560 3490 9120 3500
rect 9400 3490 9520 3500
rect 9640 3490 9990 3500
rect 2480 3480 2600 3490
rect 4080 3480 4200 3490
rect 4800 3480 4920 3490
rect 6560 3480 6800 3490
rect 8560 3480 9120 3490
rect 9400 3480 9520 3490
rect 9640 3480 9990 3490
rect 2480 3470 2600 3480
rect 4080 3470 4200 3480
rect 4800 3470 4920 3480
rect 6560 3470 6800 3480
rect 8560 3470 9120 3480
rect 9400 3470 9520 3480
rect 9640 3470 9990 3480
rect 2480 3460 2600 3470
rect 4080 3460 4200 3470
rect 4800 3460 4920 3470
rect 6560 3460 6800 3470
rect 8560 3460 9120 3470
rect 9400 3460 9520 3470
rect 9640 3460 9990 3470
rect 2360 3450 2840 3460
rect 4080 3450 4160 3460
rect 4800 3450 4840 3460
rect 5040 3450 5120 3460
rect 6560 3450 6800 3460
rect 8560 3450 9080 3460
rect 9280 3450 9440 3460
rect 9600 3450 9990 3460
rect 2360 3440 2840 3450
rect 4080 3440 4160 3450
rect 4800 3440 4840 3450
rect 5040 3440 5120 3450
rect 6560 3440 6800 3450
rect 8560 3440 9080 3450
rect 9280 3440 9440 3450
rect 9600 3440 9990 3450
rect 2360 3430 2840 3440
rect 4080 3430 4160 3440
rect 4800 3430 4840 3440
rect 5040 3430 5120 3440
rect 6560 3430 6800 3440
rect 8560 3430 9080 3440
rect 9280 3430 9440 3440
rect 9600 3430 9990 3440
rect 2360 3420 2840 3430
rect 4080 3420 4160 3430
rect 4800 3420 4840 3430
rect 5040 3420 5120 3430
rect 6560 3420 6800 3430
rect 8560 3420 9080 3430
rect 9280 3420 9440 3430
rect 9600 3420 9990 3430
rect 2240 3410 2920 3420
rect 5040 3410 5200 3420
rect 6520 3410 6720 3420
rect 8560 3410 9040 3420
rect 9200 3410 9400 3420
rect 9560 3410 9640 3420
rect 9680 3410 9990 3420
rect 2240 3400 2920 3410
rect 5040 3400 5200 3410
rect 6520 3400 6720 3410
rect 8560 3400 9040 3410
rect 9200 3400 9400 3410
rect 9560 3400 9640 3410
rect 9680 3400 9990 3410
rect 2240 3390 2920 3400
rect 5040 3390 5200 3400
rect 6520 3390 6720 3400
rect 8560 3390 9040 3400
rect 9200 3390 9400 3400
rect 9560 3390 9640 3400
rect 9680 3390 9990 3400
rect 2240 3380 2920 3390
rect 5040 3380 5200 3390
rect 6520 3380 6720 3390
rect 8560 3380 9040 3390
rect 9200 3380 9400 3390
rect 9560 3380 9640 3390
rect 9680 3380 9990 3390
rect 2200 3370 3040 3380
rect 5040 3370 5200 3380
rect 6520 3370 6680 3380
rect 8520 3370 9040 3380
rect 9160 3370 9400 3380
rect 9520 3370 9640 3380
rect 9800 3370 9990 3380
rect 2200 3360 3040 3370
rect 5040 3360 5200 3370
rect 6520 3360 6680 3370
rect 8520 3360 9040 3370
rect 9160 3360 9400 3370
rect 9520 3360 9640 3370
rect 9800 3360 9990 3370
rect 2200 3350 3040 3360
rect 5040 3350 5200 3360
rect 6520 3350 6680 3360
rect 8520 3350 9040 3360
rect 9160 3350 9400 3360
rect 9520 3350 9640 3360
rect 9800 3350 9990 3360
rect 2200 3340 3040 3350
rect 5040 3340 5200 3350
rect 6520 3340 6680 3350
rect 8520 3340 9040 3350
rect 9160 3340 9400 3350
rect 9520 3340 9640 3350
rect 9800 3340 9990 3350
rect 2200 3330 3080 3340
rect 4400 3330 4480 3340
rect 5040 3330 5200 3340
rect 6520 3330 6640 3340
rect 8520 3330 8920 3340
rect 9120 3330 9320 3340
rect 9480 3330 9640 3340
rect 9800 3330 9990 3340
rect 2200 3320 3080 3330
rect 4400 3320 4480 3330
rect 5040 3320 5200 3330
rect 6520 3320 6640 3330
rect 8520 3320 8920 3330
rect 9120 3320 9320 3330
rect 9480 3320 9640 3330
rect 9800 3320 9990 3330
rect 2200 3310 3080 3320
rect 4400 3310 4480 3320
rect 5040 3310 5200 3320
rect 6520 3310 6640 3320
rect 8520 3310 8920 3320
rect 9120 3310 9320 3320
rect 9480 3310 9640 3320
rect 9800 3310 9990 3320
rect 2200 3300 3080 3310
rect 4400 3300 4480 3310
rect 5040 3300 5200 3310
rect 6520 3300 6640 3310
rect 8520 3300 8920 3310
rect 9120 3300 9320 3310
rect 9480 3300 9640 3310
rect 9800 3300 9990 3310
rect 2160 3290 3120 3300
rect 5000 3290 5200 3300
rect 6520 3290 6560 3300
rect 8480 3290 8840 3300
rect 9120 3290 9320 3300
rect 9480 3290 9560 3300
rect 9760 3290 9960 3300
rect 2160 3280 3120 3290
rect 5000 3280 5200 3290
rect 6520 3280 6560 3290
rect 8480 3280 8840 3290
rect 9120 3280 9320 3290
rect 9480 3280 9560 3290
rect 9760 3280 9960 3290
rect 2160 3270 3120 3280
rect 5000 3270 5200 3280
rect 6520 3270 6560 3280
rect 8480 3270 8840 3280
rect 9120 3270 9320 3280
rect 9480 3270 9560 3280
rect 9760 3270 9960 3280
rect 2160 3260 3120 3270
rect 5000 3260 5200 3270
rect 6520 3260 6560 3270
rect 8480 3260 8840 3270
rect 9120 3260 9320 3270
rect 9480 3260 9560 3270
rect 9760 3260 9960 3270
rect 2120 3250 3120 3260
rect 5000 3250 5200 3260
rect 8480 3250 8960 3260
rect 9040 3250 9080 3260
rect 9160 3250 9280 3260
rect 9720 3250 9920 3260
rect 2120 3240 3120 3250
rect 5000 3240 5200 3250
rect 8480 3240 8960 3250
rect 9040 3240 9080 3250
rect 9160 3240 9280 3250
rect 9720 3240 9920 3250
rect 2120 3230 3120 3240
rect 5000 3230 5200 3240
rect 8480 3230 8960 3240
rect 9040 3230 9080 3240
rect 9160 3230 9280 3240
rect 9720 3230 9920 3240
rect 2120 3220 3120 3230
rect 5000 3220 5200 3230
rect 8480 3220 8960 3230
rect 9040 3220 9080 3230
rect 9160 3220 9280 3230
rect 9720 3220 9920 3230
rect 2120 3210 3160 3220
rect 5000 3210 5200 3220
rect 8440 3210 9000 3220
rect 9640 3210 9880 3220
rect 2120 3200 3160 3210
rect 5000 3200 5200 3210
rect 8440 3200 9000 3210
rect 9640 3200 9880 3210
rect 2120 3190 3160 3200
rect 5000 3190 5200 3200
rect 8440 3190 9000 3200
rect 9640 3190 9880 3200
rect 2120 3180 3160 3190
rect 5000 3180 5200 3190
rect 8440 3180 9000 3190
rect 9640 3180 9880 3190
rect 2120 3170 3160 3180
rect 5000 3170 5200 3180
rect 8440 3170 8880 3180
rect 9640 3170 9880 3180
rect 2120 3160 3160 3170
rect 5000 3160 5200 3170
rect 8440 3160 8880 3170
rect 9640 3160 9880 3170
rect 2120 3150 3160 3160
rect 5000 3150 5200 3160
rect 8440 3150 8880 3160
rect 9640 3150 9880 3160
rect 2120 3140 3160 3150
rect 5000 3140 5200 3150
rect 8440 3140 8880 3150
rect 9640 3140 9880 3150
rect 2120 3130 3160 3140
rect 5000 3130 5200 3140
rect 8400 3130 8800 3140
rect 9560 3130 9840 3140
rect 2120 3120 3160 3130
rect 5000 3120 5200 3130
rect 8400 3120 8800 3130
rect 9560 3120 9840 3130
rect 2120 3110 3160 3120
rect 5000 3110 5200 3120
rect 8400 3110 8800 3120
rect 9560 3110 9840 3120
rect 2120 3100 3160 3110
rect 5000 3100 5200 3110
rect 8400 3100 8800 3110
rect 9560 3100 9840 3110
rect 2120 3090 3160 3100
rect 3920 3090 3960 3100
rect 5000 3090 5160 3100
rect 8440 3090 8840 3100
rect 9520 3090 9800 3100
rect 2120 3080 3160 3090
rect 3920 3080 3960 3090
rect 5000 3080 5160 3090
rect 8440 3080 8840 3090
rect 9520 3080 9800 3090
rect 2120 3070 3160 3080
rect 3920 3070 3960 3080
rect 5000 3070 5160 3080
rect 8440 3070 8840 3080
rect 9520 3070 9800 3080
rect 2120 3060 3160 3070
rect 3920 3060 3960 3070
rect 5000 3060 5160 3070
rect 8440 3060 8840 3070
rect 9520 3060 9800 3070
rect 2120 3050 3120 3060
rect 3920 3050 4040 3060
rect 4360 3050 4400 3060
rect 5000 3050 5120 3060
rect 8360 3050 8400 3060
rect 8440 3050 8720 3060
rect 9520 3050 9760 3060
rect 9960 3050 9990 3060
rect 2120 3040 3120 3050
rect 3920 3040 4040 3050
rect 4360 3040 4400 3050
rect 5000 3040 5120 3050
rect 8360 3040 8400 3050
rect 8440 3040 8720 3050
rect 9520 3040 9760 3050
rect 9960 3040 9990 3050
rect 2120 3030 3120 3040
rect 3920 3030 4040 3040
rect 4360 3030 4400 3040
rect 5000 3030 5120 3040
rect 8360 3030 8400 3040
rect 8440 3030 8720 3040
rect 9520 3030 9760 3040
rect 9960 3030 9990 3040
rect 2120 3020 3120 3030
rect 3920 3020 4040 3030
rect 4360 3020 4400 3030
rect 5000 3020 5120 3030
rect 8360 3020 8400 3030
rect 8440 3020 8720 3030
rect 9520 3020 9760 3030
rect 9960 3020 9990 3030
rect 2080 3010 3120 3020
rect 3920 3010 4000 3020
rect 8360 3010 8400 3020
rect 8440 3010 8600 3020
rect 9480 3010 9760 3020
rect 9960 3010 9990 3020
rect 2080 3000 3120 3010
rect 3920 3000 4000 3010
rect 8360 3000 8400 3010
rect 8440 3000 8600 3010
rect 9480 3000 9760 3010
rect 9960 3000 9990 3010
rect 2080 2990 3120 3000
rect 3920 2990 4000 3000
rect 8360 2990 8400 3000
rect 8440 2990 8600 3000
rect 9480 2990 9760 3000
rect 9960 2990 9990 3000
rect 2080 2980 3120 2990
rect 3920 2980 4000 2990
rect 8360 2980 8400 2990
rect 8440 2980 8600 2990
rect 9480 2980 9760 2990
rect 9960 2980 9990 2990
rect 2080 2970 3120 2980
rect 3920 2970 4000 2980
rect 4080 2970 4120 2980
rect 8320 2970 8400 2980
rect 8440 2970 8560 2980
rect 9480 2970 9880 2980
rect 9960 2970 9990 2980
rect 2080 2960 3120 2970
rect 3920 2960 4000 2970
rect 4080 2960 4120 2970
rect 8320 2960 8400 2970
rect 8440 2960 8560 2970
rect 9480 2960 9880 2970
rect 9960 2960 9990 2970
rect 2080 2950 3120 2960
rect 3920 2950 4000 2960
rect 4080 2950 4120 2960
rect 8320 2950 8400 2960
rect 8440 2950 8560 2960
rect 9480 2950 9880 2960
rect 9960 2950 9990 2960
rect 2080 2940 3120 2950
rect 3920 2940 4000 2950
rect 4080 2940 4120 2950
rect 8320 2940 8400 2950
rect 8440 2940 8560 2950
rect 9480 2940 9880 2950
rect 9960 2940 9990 2950
rect 2080 2930 3120 2940
rect 4040 2930 4200 2940
rect 8280 2930 8520 2940
rect 9440 2930 9680 2940
rect 9720 2930 9920 2940
rect 9960 2930 9990 2940
rect 2080 2920 3120 2930
rect 4040 2920 4200 2930
rect 8280 2920 8520 2930
rect 9440 2920 9680 2930
rect 9720 2920 9920 2930
rect 9960 2920 9990 2930
rect 2080 2910 3120 2920
rect 4040 2910 4200 2920
rect 8280 2910 8520 2920
rect 9440 2910 9680 2920
rect 9720 2910 9920 2920
rect 9960 2910 9990 2920
rect 2080 2900 3120 2910
rect 4040 2900 4200 2910
rect 8280 2900 8520 2910
rect 9440 2900 9680 2910
rect 9720 2900 9920 2910
rect 9960 2900 9990 2910
rect 2080 2890 3120 2900
rect 4000 2890 4240 2900
rect 8280 2890 8520 2900
rect 9400 2890 9680 2900
rect 9720 2890 9920 2900
rect 2080 2880 3120 2890
rect 4000 2880 4240 2890
rect 8280 2880 8520 2890
rect 9400 2880 9680 2890
rect 9720 2880 9920 2890
rect 2080 2870 3120 2880
rect 4000 2870 4240 2880
rect 8280 2870 8520 2880
rect 9400 2870 9680 2880
rect 9720 2870 9920 2880
rect 2080 2860 3120 2870
rect 4000 2860 4240 2870
rect 8280 2860 8520 2870
rect 9400 2860 9680 2870
rect 9720 2860 9920 2870
rect 2040 2850 3080 2860
rect 4000 2850 4240 2860
rect 7240 2850 7520 2860
rect 8240 2850 8520 2860
rect 9400 2850 9920 2860
rect 2040 2840 3080 2850
rect 4000 2840 4240 2850
rect 7240 2840 7520 2850
rect 8240 2840 8520 2850
rect 9400 2840 9920 2850
rect 2040 2830 3080 2840
rect 4000 2830 4240 2840
rect 7240 2830 7520 2840
rect 8240 2830 8520 2840
rect 9400 2830 9920 2840
rect 2040 2820 3080 2830
rect 4000 2820 4240 2830
rect 7240 2820 7520 2830
rect 8240 2820 8520 2830
rect 9400 2820 9920 2830
rect 2080 2810 2240 2820
rect 2400 2810 2840 2820
rect 4000 2810 4240 2820
rect 7200 2810 7560 2820
rect 8200 2810 8520 2820
rect 9480 2810 9560 2820
rect 9680 2810 9920 2820
rect 2080 2800 2240 2810
rect 2400 2800 2840 2810
rect 4000 2800 4240 2810
rect 7200 2800 7560 2810
rect 8200 2800 8520 2810
rect 9480 2800 9560 2810
rect 9680 2800 9920 2810
rect 2080 2790 2240 2800
rect 2400 2790 2840 2800
rect 4000 2790 4240 2800
rect 7200 2790 7560 2800
rect 8200 2790 8520 2800
rect 9480 2790 9560 2800
rect 9680 2790 9920 2800
rect 2080 2780 2240 2790
rect 2400 2780 2840 2790
rect 4000 2780 4240 2790
rect 7200 2780 7560 2790
rect 8200 2780 8520 2790
rect 9480 2780 9560 2790
rect 9680 2780 9920 2790
rect 2080 2770 2200 2780
rect 2440 2770 2800 2780
rect 3040 2770 3080 2780
rect 3960 2770 4160 2780
rect 4200 2770 4240 2780
rect 7120 2770 7600 2780
rect 8160 2770 8560 2780
rect 9320 2770 9400 2780
rect 9560 2770 9600 2780
rect 9720 2770 9880 2780
rect 2080 2760 2200 2770
rect 2440 2760 2800 2770
rect 3040 2760 3080 2770
rect 3960 2760 4160 2770
rect 4200 2760 4240 2770
rect 7120 2760 7600 2770
rect 8160 2760 8560 2770
rect 9320 2760 9400 2770
rect 9560 2760 9600 2770
rect 9720 2760 9880 2770
rect 2080 2750 2200 2760
rect 2440 2750 2800 2760
rect 3040 2750 3080 2760
rect 3960 2750 4160 2760
rect 4200 2750 4240 2760
rect 7120 2750 7600 2760
rect 8160 2750 8560 2760
rect 9320 2750 9400 2760
rect 9560 2750 9600 2760
rect 9720 2750 9880 2760
rect 2080 2740 2200 2750
rect 2440 2740 2800 2750
rect 3040 2740 3080 2750
rect 3960 2740 4160 2750
rect 4200 2740 4240 2750
rect 7120 2740 7600 2750
rect 8160 2740 8560 2750
rect 9320 2740 9400 2750
rect 9560 2740 9600 2750
rect 9720 2740 9880 2750
rect 2080 2730 2280 2740
rect 2480 2730 2760 2740
rect 2960 2730 3120 2740
rect 3960 2730 4240 2740
rect 7040 2730 7640 2740
rect 8160 2730 8560 2740
rect 9320 2730 9360 2740
rect 9400 2730 9560 2740
rect 9720 2730 9880 2740
rect 2080 2720 2280 2730
rect 2480 2720 2760 2730
rect 2960 2720 3120 2730
rect 3960 2720 4240 2730
rect 7040 2720 7640 2730
rect 8160 2720 8560 2730
rect 9320 2720 9360 2730
rect 9400 2720 9560 2730
rect 9720 2720 9880 2730
rect 2080 2710 2280 2720
rect 2480 2710 2760 2720
rect 2960 2710 3120 2720
rect 3960 2710 4240 2720
rect 7040 2710 7640 2720
rect 8160 2710 8560 2720
rect 9320 2710 9360 2720
rect 9400 2710 9560 2720
rect 9720 2710 9880 2720
rect 2080 2700 2280 2710
rect 2480 2700 2760 2710
rect 2960 2700 3120 2710
rect 3960 2700 4240 2710
rect 7040 2700 7640 2710
rect 8160 2700 8560 2710
rect 9320 2700 9360 2710
rect 9400 2700 9560 2710
rect 9720 2700 9880 2710
rect 2040 2690 2200 2700
rect 2480 2690 2760 2700
rect 3920 2690 4200 2700
rect 6960 2690 7680 2700
rect 8120 2690 8560 2700
rect 9280 2690 9640 2700
rect 9720 2690 9920 2700
rect 2040 2680 2200 2690
rect 2480 2680 2760 2690
rect 3920 2680 4200 2690
rect 6960 2680 7680 2690
rect 8120 2680 8560 2690
rect 9280 2680 9640 2690
rect 9720 2680 9920 2690
rect 2040 2670 2200 2680
rect 2480 2670 2760 2680
rect 3920 2670 4200 2680
rect 6960 2670 7680 2680
rect 8120 2670 8560 2680
rect 9280 2670 9640 2680
rect 9720 2670 9920 2680
rect 2040 2660 2200 2670
rect 2480 2660 2760 2670
rect 3920 2660 4200 2670
rect 6960 2660 7680 2670
rect 8120 2660 8560 2670
rect 9280 2660 9640 2670
rect 9720 2660 9920 2670
rect 2480 2650 2720 2660
rect 3920 2650 4200 2660
rect 6920 2650 7160 2660
rect 7200 2650 7680 2660
rect 8080 2650 8520 2660
rect 8560 2650 8600 2660
rect 9240 2650 9720 2660
rect 9800 2650 9840 2660
rect 2480 2640 2720 2650
rect 3920 2640 4200 2650
rect 6920 2640 7160 2650
rect 7200 2640 7680 2650
rect 8080 2640 8520 2650
rect 8560 2640 8600 2650
rect 9240 2640 9720 2650
rect 9800 2640 9840 2650
rect 2480 2630 2720 2640
rect 3920 2630 4200 2640
rect 6920 2630 7160 2640
rect 7200 2630 7680 2640
rect 8080 2630 8520 2640
rect 8560 2630 8600 2640
rect 9240 2630 9720 2640
rect 9800 2630 9840 2640
rect 2480 2620 2720 2630
rect 3920 2620 4200 2630
rect 6920 2620 7160 2630
rect 7200 2620 7680 2630
rect 8080 2620 8520 2630
rect 8560 2620 8600 2630
rect 9240 2620 9720 2630
rect 9800 2620 9840 2630
rect 2480 2610 2720 2620
rect 3960 2610 4200 2620
rect 6880 2610 7120 2620
rect 7280 2610 7720 2620
rect 8040 2610 8400 2620
rect 8480 2610 8560 2620
rect 9200 2610 9800 2620
rect 2480 2600 2720 2610
rect 3960 2600 4200 2610
rect 6880 2600 7120 2610
rect 7280 2600 7720 2610
rect 8040 2600 8400 2610
rect 8480 2600 8560 2610
rect 9200 2600 9800 2610
rect 2480 2590 2720 2600
rect 3960 2590 4200 2600
rect 6880 2590 7120 2600
rect 7280 2590 7720 2600
rect 8040 2590 8400 2600
rect 8480 2590 8560 2600
rect 9200 2590 9800 2600
rect 2480 2580 2720 2590
rect 3960 2580 4200 2590
rect 6880 2580 7120 2590
rect 7280 2580 7720 2590
rect 8040 2580 8400 2590
rect 8480 2580 8560 2590
rect 9200 2580 9800 2590
rect 2440 2570 2720 2580
rect 4000 2570 4040 2580
rect 4120 2570 4160 2580
rect 6840 2570 7120 2580
rect 7320 2570 7760 2580
rect 8000 2570 8400 2580
rect 9200 2570 9360 2580
rect 9600 2570 9880 2580
rect 2440 2560 2720 2570
rect 4000 2560 4040 2570
rect 4120 2560 4160 2570
rect 6840 2560 7120 2570
rect 7320 2560 7760 2570
rect 8000 2560 8400 2570
rect 9200 2560 9360 2570
rect 9600 2560 9880 2570
rect 2440 2550 2720 2560
rect 4000 2550 4040 2560
rect 4120 2550 4160 2560
rect 6840 2550 7120 2560
rect 7320 2550 7760 2560
rect 8000 2550 8400 2560
rect 9200 2550 9360 2560
rect 9600 2550 9880 2560
rect 2440 2540 2720 2550
rect 4000 2540 4040 2550
rect 4120 2540 4160 2550
rect 6840 2540 7120 2550
rect 7320 2540 7760 2550
rect 8000 2540 8400 2550
rect 9200 2540 9360 2550
rect 9600 2540 9880 2550
rect 2400 2530 2840 2540
rect 2920 2530 3080 2540
rect 6800 2530 7200 2540
rect 7360 2530 7800 2540
rect 7960 2530 8400 2540
rect 9160 2530 9280 2540
rect 9680 2530 9960 2540
rect 2400 2520 2840 2530
rect 2920 2520 3080 2530
rect 6800 2520 7200 2530
rect 7360 2520 7800 2530
rect 7960 2520 8400 2530
rect 9160 2520 9280 2530
rect 9680 2520 9960 2530
rect 2400 2510 2840 2520
rect 2920 2510 3080 2520
rect 6800 2510 7200 2520
rect 7360 2510 7800 2520
rect 7960 2510 8400 2520
rect 9160 2510 9280 2520
rect 9680 2510 9960 2520
rect 2400 2500 2840 2510
rect 2920 2500 3080 2510
rect 6800 2500 7200 2510
rect 7360 2500 7800 2510
rect 7960 2500 8400 2510
rect 9160 2500 9280 2510
rect 9680 2500 9960 2510
rect 1960 2490 2200 2500
rect 2320 2490 3040 2500
rect 3120 2490 3200 2500
rect 6880 2490 7240 2500
rect 7360 2490 7800 2500
rect 7880 2490 8400 2500
rect 9160 2490 9240 2500
rect 9720 2490 9990 2500
rect 1960 2480 2200 2490
rect 2320 2480 3040 2490
rect 3120 2480 3200 2490
rect 6880 2480 7240 2490
rect 7360 2480 7800 2490
rect 7880 2480 8400 2490
rect 9160 2480 9240 2490
rect 9720 2480 9990 2490
rect 1960 2470 2200 2480
rect 2320 2470 3040 2480
rect 3120 2470 3200 2480
rect 6880 2470 7240 2480
rect 7360 2470 7800 2480
rect 7880 2470 8400 2480
rect 9160 2470 9240 2480
rect 9720 2470 9990 2480
rect 1960 2460 2200 2470
rect 2320 2460 3040 2470
rect 3120 2460 3200 2470
rect 6880 2460 7240 2470
rect 7360 2460 7800 2470
rect 7880 2460 8400 2470
rect 9160 2460 9240 2470
rect 9720 2460 9990 2470
rect 1960 2450 2080 2460
rect 2280 2450 3200 2460
rect 6880 2450 7280 2460
rect 7440 2450 8400 2460
rect 9160 2450 9200 2460
rect 9800 2450 9990 2460
rect 1960 2440 2080 2450
rect 2280 2440 3200 2450
rect 6880 2440 7280 2450
rect 7440 2440 8400 2450
rect 9160 2440 9200 2450
rect 9800 2440 9990 2450
rect 1960 2430 2080 2440
rect 2280 2430 3200 2440
rect 6880 2430 7280 2440
rect 7440 2430 8400 2440
rect 9160 2430 9200 2440
rect 9800 2430 9990 2440
rect 1960 2420 2080 2430
rect 2280 2420 3200 2430
rect 6880 2420 7280 2430
rect 7440 2420 8400 2430
rect 9160 2420 9200 2430
rect 9800 2420 9990 2430
rect 1960 2410 3200 2420
rect 6960 2410 7360 2420
rect 7480 2410 8400 2420
rect 9200 2410 9240 2420
rect 9840 2410 9990 2420
rect 1960 2400 3200 2410
rect 6960 2400 7360 2410
rect 7480 2400 8400 2410
rect 9200 2400 9240 2410
rect 9840 2400 9990 2410
rect 1960 2390 3200 2400
rect 6960 2390 7360 2400
rect 7480 2390 8400 2400
rect 9200 2390 9240 2400
rect 9840 2390 9990 2400
rect 1960 2380 3200 2390
rect 6960 2380 7360 2390
rect 7480 2380 8400 2390
rect 9200 2380 9240 2390
rect 9840 2380 9990 2390
rect 1960 2370 3240 2380
rect 7120 2370 7400 2380
rect 7520 2370 8400 2380
rect 8680 2370 8760 2380
rect 9840 2370 9990 2380
rect 1960 2360 3240 2370
rect 7120 2360 7400 2370
rect 7520 2360 8400 2370
rect 8680 2360 8760 2370
rect 9840 2360 9990 2370
rect 1960 2350 3240 2360
rect 7120 2350 7400 2360
rect 7520 2350 8400 2360
rect 8680 2350 8760 2360
rect 9840 2350 9990 2360
rect 1960 2340 3240 2350
rect 7120 2340 7400 2350
rect 7520 2340 8400 2350
rect 8680 2340 8760 2350
rect 9840 2340 9990 2350
rect 1920 2330 3240 2340
rect 7200 2330 7480 2340
rect 7560 2330 8360 2340
rect 8640 2330 8760 2340
rect 8840 2330 8960 2340
rect 9840 2330 9990 2340
rect 1920 2320 3240 2330
rect 7200 2320 7480 2330
rect 7560 2320 8360 2330
rect 8640 2320 8760 2330
rect 8840 2320 8960 2330
rect 9840 2320 9990 2330
rect 1920 2310 3240 2320
rect 7200 2310 7480 2320
rect 7560 2310 8360 2320
rect 8640 2310 8760 2320
rect 8840 2310 8960 2320
rect 9840 2310 9990 2320
rect 1920 2300 3240 2310
rect 7200 2300 7480 2310
rect 7560 2300 8360 2310
rect 8640 2300 8760 2310
rect 8840 2300 8960 2310
rect 9840 2300 9990 2310
rect 1920 2290 3240 2300
rect 7400 2290 7480 2300
rect 7640 2290 8360 2300
rect 8680 2290 8720 2300
rect 9840 2290 9990 2300
rect 1920 2280 3240 2290
rect 7400 2280 7480 2290
rect 7640 2280 8360 2290
rect 8680 2280 8720 2290
rect 9840 2280 9990 2290
rect 1920 2270 3240 2280
rect 7400 2270 7480 2280
rect 7640 2270 8360 2280
rect 8680 2270 8720 2280
rect 9840 2270 9990 2280
rect 1920 2260 3240 2270
rect 7400 2260 7480 2270
rect 7640 2260 8360 2270
rect 8680 2260 8720 2270
rect 9840 2260 9990 2270
rect 1920 2250 2680 2260
rect 2720 2250 3240 2260
rect 7400 2250 7480 2260
rect 7640 2250 8360 2260
rect 8880 2250 9000 2260
rect 9800 2250 9990 2260
rect 1920 2240 2680 2250
rect 2720 2240 3240 2250
rect 7400 2240 7480 2250
rect 7640 2240 8360 2250
rect 8880 2240 9000 2250
rect 9800 2240 9990 2250
rect 1920 2230 2680 2240
rect 2720 2230 3240 2240
rect 7400 2230 7480 2240
rect 7640 2230 8360 2240
rect 8880 2230 9000 2240
rect 9800 2230 9990 2240
rect 1920 2220 2680 2230
rect 2720 2220 3240 2230
rect 7400 2220 7480 2230
rect 7640 2220 8360 2230
rect 8880 2220 9000 2230
rect 9800 2220 9990 2230
rect 1920 2210 2440 2220
rect 2840 2210 3240 2220
rect 7400 2210 7480 2220
rect 7720 2210 8360 2220
rect 9240 2210 9320 2220
rect 9840 2210 9960 2220
rect 1920 2200 2440 2210
rect 2840 2200 3240 2210
rect 7400 2200 7480 2210
rect 7720 2200 8360 2210
rect 9240 2200 9320 2210
rect 9840 2200 9960 2210
rect 1920 2190 2440 2200
rect 2840 2190 3240 2200
rect 7400 2190 7480 2200
rect 7720 2190 8360 2200
rect 9240 2190 9320 2200
rect 9840 2190 9960 2200
rect 1920 2180 2440 2190
rect 2840 2180 3240 2190
rect 7400 2180 7480 2190
rect 7720 2180 8360 2190
rect 9240 2180 9320 2190
rect 9840 2180 9960 2190
rect 1920 2170 2240 2180
rect 2280 2170 2360 2180
rect 2840 2170 3240 2180
rect 7840 2170 8360 2180
rect 9280 2170 9400 2180
rect 9800 2170 9990 2180
rect 1920 2160 2240 2170
rect 2280 2160 2360 2170
rect 2840 2160 3240 2170
rect 7840 2160 8360 2170
rect 9280 2160 9400 2170
rect 9800 2160 9990 2170
rect 1920 2150 2240 2160
rect 2280 2150 2360 2160
rect 2840 2150 3240 2160
rect 7840 2150 8360 2160
rect 9280 2150 9400 2160
rect 9800 2150 9990 2160
rect 1920 2140 2240 2150
rect 2280 2140 2360 2150
rect 2840 2140 3240 2150
rect 7840 2140 8360 2150
rect 9280 2140 9400 2150
rect 9800 2140 9990 2150
rect 1920 2130 2200 2140
rect 2280 2130 2360 2140
rect 2800 2130 3240 2140
rect 7880 2130 8360 2140
rect 9360 2130 9480 2140
rect 9760 2130 9990 2140
rect 1920 2120 2200 2130
rect 2280 2120 2360 2130
rect 2800 2120 3240 2130
rect 7880 2120 8360 2130
rect 9360 2120 9480 2130
rect 9760 2120 9990 2130
rect 1920 2110 2200 2120
rect 2280 2110 2360 2120
rect 2800 2110 3240 2120
rect 7880 2110 8360 2120
rect 9360 2110 9480 2120
rect 9760 2110 9990 2120
rect 1920 2100 2200 2110
rect 2280 2100 2360 2110
rect 2800 2100 3240 2110
rect 7880 2100 8360 2110
rect 9360 2100 9480 2110
rect 9760 2100 9990 2110
rect 1960 2090 2200 2100
rect 2240 2090 3200 2100
rect 7920 2090 8360 2100
rect 9720 2090 9990 2100
rect 1960 2080 2200 2090
rect 2240 2080 3200 2090
rect 7920 2080 8360 2090
rect 9720 2080 9990 2090
rect 1960 2070 2200 2080
rect 2240 2070 3200 2080
rect 7920 2070 8360 2080
rect 9720 2070 9990 2080
rect 1960 2060 2200 2070
rect 2240 2060 3200 2070
rect 7920 2060 8360 2070
rect 9720 2060 9990 2070
rect 2000 2050 2120 2060
rect 2200 2050 3160 2060
rect 8000 2050 8360 2060
rect 9480 2050 9600 2060
rect 9680 2050 9990 2060
rect 2000 2040 2120 2050
rect 2200 2040 3160 2050
rect 8000 2040 8360 2050
rect 9480 2040 9600 2050
rect 9680 2040 9990 2050
rect 2000 2030 2120 2040
rect 2200 2030 3160 2040
rect 8000 2030 8360 2040
rect 9480 2030 9600 2040
rect 9680 2030 9990 2040
rect 2000 2020 2120 2030
rect 2200 2020 3160 2030
rect 8000 2020 8360 2030
rect 9480 2020 9600 2030
rect 9680 2020 9990 2030
rect 2200 2010 3120 2020
rect 8000 2010 8360 2020
rect 9200 2010 9990 2020
rect 2200 2000 3120 2010
rect 8000 2000 8360 2010
rect 9200 2000 9990 2010
rect 2200 1990 3120 2000
rect 8000 1990 8360 2000
rect 9200 1990 9990 2000
rect 2200 1980 3120 1990
rect 8000 1980 8360 1990
rect 9200 1980 9990 1990
rect 2160 1970 3120 1980
rect 7960 1970 8360 1980
rect 9120 1970 9880 1980
rect 9960 1970 9990 1980
rect 2160 1960 3120 1970
rect 7960 1960 8360 1970
rect 9120 1960 9880 1970
rect 9960 1960 9990 1970
rect 2160 1950 3120 1960
rect 7960 1950 8360 1960
rect 9120 1950 9880 1960
rect 9960 1950 9990 1960
rect 2160 1940 3120 1950
rect 7960 1940 8360 1950
rect 9120 1940 9880 1950
rect 9960 1940 9990 1950
rect 2160 1930 2600 1940
rect 2760 1930 3120 1940
rect 7920 1930 8360 1940
rect 8720 1930 8960 1940
rect 9120 1930 9600 1940
rect 9720 1930 9880 1940
rect 2160 1920 2600 1930
rect 2760 1920 3120 1930
rect 7920 1920 8360 1930
rect 8720 1920 8960 1930
rect 9120 1920 9600 1930
rect 9720 1920 9880 1930
rect 2160 1910 2600 1920
rect 2760 1910 3120 1920
rect 7920 1910 8360 1920
rect 8720 1910 8960 1920
rect 9120 1910 9600 1920
rect 9720 1910 9880 1920
rect 2160 1900 2600 1910
rect 2760 1900 3120 1910
rect 7920 1900 8360 1910
rect 8720 1900 8960 1910
rect 9120 1900 9600 1910
rect 9720 1900 9880 1910
rect 2160 1890 2400 1900
rect 3000 1890 3120 1900
rect 7920 1890 8360 1900
rect 8640 1890 9000 1900
rect 9200 1890 9680 1900
rect 9760 1890 9990 1900
rect 2160 1880 2400 1890
rect 3000 1880 3120 1890
rect 7920 1880 8360 1890
rect 8640 1880 9000 1890
rect 9200 1880 9680 1890
rect 9760 1880 9990 1890
rect 2160 1870 2400 1880
rect 3000 1870 3120 1880
rect 7920 1870 8360 1880
rect 8640 1870 9000 1880
rect 9200 1870 9680 1880
rect 9760 1870 9990 1880
rect 2160 1860 2400 1870
rect 3000 1860 3120 1870
rect 7920 1860 8360 1870
rect 8640 1860 9000 1870
rect 9200 1860 9680 1870
rect 9760 1860 9990 1870
rect 2160 1850 2200 1860
rect 2960 1850 3120 1860
rect 7920 1850 8360 1860
rect 8640 1850 8960 1860
rect 9400 1850 9680 1860
rect 9800 1850 9960 1860
rect 2160 1840 2200 1850
rect 2960 1840 3120 1850
rect 7920 1840 8360 1850
rect 8640 1840 8960 1850
rect 9400 1840 9680 1850
rect 9800 1840 9960 1850
rect 2160 1830 2200 1840
rect 2960 1830 3120 1840
rect 7920 1830 8360 1840
rect 8640 1830 8960 1840
rect 9400 1830 9680 1840
rect 9800 1830 9960 1840
rect 2160 1820 2200 1830
rect 2960 1820 3120 1830
rect 7920 1820 8360 1830
rect 8640 1820 8960 1830
rect 9400 1820 9680 1830
rect 9800 1820 9960 1830
rect 2120 1810 2200 1820
rect 2920 1810 3160 1820
rect 7920 1810 8360 1820
rect 8640 1810 8920 1820
rect 9320 1810 9400 1820
rect 9440 1810 9680 1820
rect 9800 1810 9920 1820
rect 2120 1800 2200 1810
rect 2920 1800 3160 1810
rect 7920 1800 8360 1810
rect 8640 1800 8920 1810
rect 9320 1800 9400 1810
rect 9440 1800 9680 1810
rect 9800 1800 9920 1810
rect 2120 1790 2200 1800
rect 2920 1790 3160 1800
rect 7920 1790 8360 1800
rect 8640 1790 8920 1800
rect 9320 1790 9400 1800
rect 9440 1790 9680 1800
rect 9800 1790 9920 1800
rect 2120 1780 2200 1790
rect 2920 1780 3160 1790
rect 7920 1780 8360 1790
rect 8640 1780 8920 1790
rect 9320 1780 9400 1790
rect 9440 1780 9680 1790
rect 9800 1780 9920 1790
rect 2040 1770 2200 1780
rect 2240 1770 2360 1780
rect 2760 1770 3160 1780
rect 4080 1770 4200 1780
rect 7040 1770 7120 1780
rect 7920 1770 8360 1780
rect 8600 1770 8920 1780
rect 9240 1770 9680 1780
rect 9800 1770 9920 1780
rect 9960 1770 9990 1780
rect 2040 1760 2200 1770
rect 2240 1760 2360 1770
rect 2760 1760 3160 1770
rect 4080 1760 4200 1770
rect 7040 1760 7120 1770
rect 7920 1760 8360 1770
rect 8600 1760 8920 1770
rect 9240 1760 9680 1770
rect 9800 1760 9920 1770
rect 9960 1760 9990 1770
rect 2040 1750 2200 1760
rect 2240 1750 2360 1760
rect 2760 1750 3160 1760
rect 4080 1750 4200 1760
rect 7040 1750 7120 1760
rect 7920 1750 8360 1760
rect 8600 1750 8920 1760
rect 9240 1750 9680 1760
rect 9800 1750 9920 1760
rect 9960 1750 9990 1760
rect 2040 1740 2200 1750
rect 2240 1740 2360 1750
rect 2760 1740 3160 1750
rect 4080 1740 4200 1750
rect 7040 1740 7120 1750
rect 7920 1740 8360 1750
rect 8600 1740 8920 1750
rect 9240 1740 9680 1750
rect 9800 1740 9920 1750
rect 9960 1740 9990 1750
rect 2040 1730 2440 1740
rect 2680 1730 3160 1740
rect 4080 1730 4160 1740
rect 7000 1730 7120 1740
rect 7960 1730 8320 1740
rect 8600 1730 8880 1740
rect 9240 1730 9680 1740
rect 9800 1730 9880 1740
rect 9960 1730 9990 1740
rect 2040 1720 2440 1730
rect 2680 1720 3160 1730
rect 4080 1720 4160 1730
rect 7000 1720 7120 1730
rect 7960 1720 8320 1730
rect 8600 1720 8880 1730
rect 9240 1720 9680 1730
rect 9800 1720 9880 1730
rect 9960 1720 9990 1730
rect 2040 1710 2440 1720
rect 2680 1710 3160 1720
rect 4080 1710 4160 1720
rect 7000 1710 7120 1720
rect 7960 1710 8320 1720
rect 8600 1710 8880 1720
rect 9240 1710 9680 1720
rect 9800 1710 9880 1720
rect 9960 1710 9990 1720
rect 2040 1700 2440 1710
rect 2680 1700 3160 1710
rect 4080 1700 4160 1710
rect 7000 1700 7120 1710
rect 7960 1700 8320 1710
rect 8600 1700 8880 1710
rect 9240 1700 9680 1710
rect 9800 1700 9880 1710
rect 9960 1700 9990 1710
rect 2040 1690 2480 1700
rect 2680 1690 3120 1700
rect 7000 1690 7120 1700
rect 7960 1690 8320 1700
rect 8600 1690 8840 1700
rect 9080 1690 9120 1700
rect 9240 1690 9720 1700
rect 9800 1690 9880 1700
rect 9920 1690 9990 1700
rect 2040 1680 2480 1690
rect 2680 1680 3120 1690
rect 7000 1680 7120 1690
rect 7960 1680 8320 1690
rect 8600 1680 8840 1690
rect 9080 1680 9120 1690
rect 9240 1680 9720 1690
rect 9800 1680 9880 1690
rect 9920 1680 9990 1690
rect 2040 1670 2480 1680
rect 2680 1670 3120 1680
rect 7000 1670 7120 1680
rect 7960 1670 8320 1680
rect 8600 1670 8840 1680
rect 9080 1670 9120 1680
rect 9240 1670 9720 1680
rect 9800 1670 9880 1680
rect 9920 1670 9990 1680
rect 2040 1660 2480 1670
rect 2680 1660 3120 1670
rect 7000 1660 7120 1670
rect 7960 1660 8320 1670
rect 8600 1660 8840 1670
rect 9080 1660 9120 1670
rect 9240 1660 9720 1670
rect 9800 1660 9880 1670
rect 9920 1660 9990 1670
rect 2080 1650 2400 1660
rect 2760 1650 3080 1660
rect 7000 1650 7160 1660
rect 7960 1650 8320 1660
rect 8640 1650 8840 1660
rect 9080 1650 9120 1660
rect 9240 1650 9840 1660
rect 9880 1650 9990 1660
rect 2080 1640 2400 1650
rect 2760 1640 3080 1650
rect 7000 1640 7160 1650
rect 7960 1640 8320 1650
rect 8640 1640 8840 1650
rect 9080 1640 9120 1650
rect 9240 1640 9840 1650
rect 9880 1640 9990 1650
rect 2080 1630 2400 1640
rect 2760 1630 3080 1640
rect 7000 1630 7160 1640
rect 7960 1630 8320 1640
rect 8640 1630 8840 1640
rect 9080 1630 9120 1640
rect 9240 1630 9840 1640
rect 9880 1630 9990 1640
rect 2080 1620 2400 1630
rect 2760 1620 3080 1630
rect 7000 1620 7160 1630
rect 7960 1620 8320 1630
rect 8640 1620 8840 1630
rect 9080 1620 9120 1630
rect 9240 1620 9840 1630
rect 9880 1620 9990 1630
rect 2080 1610 2360 1620
rect 2720 1610 3040 1620
rect 7000 1610 7120 1620
rect 7960 1610 8320 1620
rect 8640 1610 8680 1620
rect 8720 1610 8760 1620
rect 9080 1610 9120 1620
rect 9200 1610 9840 1620
rect 9880 1610 9990 1620
rect 2080 1600 2360 1610
rect 2720 1600 3040 1610
rect 7000 1600 7120 1610
rect 7960 1600 8320 1610
rect 8640 1600 8680 1610
rect 8720 1600 8760 1610
rect 9080 1600 9120 1610
rect 9200 1600 9840 1610
rect 9880 1600 9990 1610
rect 2080 1590 2360 1600
rect 2720 1590 3040 1600
rect 7000 1590 7120 1600
rect 7960 1590 8320 1600
rect 8640 1590 8680 1600
rect 8720 1590 8760 1600
rect 9080 1590 9120 1600
rect 9200 1590 9840 1600
rect 9880 1590 9990 1600
rect 2080 1580 2360 1590
rect 2720 1580 3040 1590
rect 7000 1580 7120 1590
rect 7960 1580 8320 1590
rect 8640 1580 8680 1590
rect 8720 1580 8760 1590
rect 9080 1580 9120 1590
rect 9200 1580 9840 1590
rect 9880 1580 9990 1590
rect 2120 1570 2440 1580
rect 2520 1570 2960 1580
rect 4280 1570 4320 1580
rect 7000 1570 7160 1580
rect 8000 1570 8280 1580
rect 8600 1570 8680 1580
rect 9080 1570 9720 1580
rect 2120 1560 2440 1570
rect 2520 1560 2960 1570
rect 4280 1560 4320 1570
rect 7000 1560 7160 1570
rect 8000 1560 8280 1570
rect 8600 1560 8680 1570
rect 9080 1560 9720 1570
rect 2120 1550 2440 1560
rect 2520 1550 2960 1560
rect 4280 1550 4320 1560
rect 7000 1550 7160 1560
rect 8000 1550 8280 1560
rect 8600 1550 8680 1560
rect 9080 1550 9720 1560
rect 2120 1540 2440 1550
rect 2520 1540 2960 1550
rect 4280 1540 4320 1550
rect 7000 1540 7160 1550
rect 8000 1540 8280 1550
rect 8600 1540 8680 1550
rect 9080 1540 9720 1550
rect 2200 1530 2920 1540
rect 4240 1530 4320 1540
rect 7000 1530 7200 1540
rect 8000 1530 8280 1540
rect 8640 1530 8680 1540
rect 9080 1530 9720 1540
rect 9840 1530 9880 1540
rect 2200 1520 2920 1530
rect 4240 1520 4320 1530
rect 7000 1520 7200 1530
rect 8000 1520 8280 1530
rect 8640 1520 8680 1530
rect 9080 1520 9720 1530
rect 9840 1520 9880 1530
rect 2200 1510 2920 1520
rect 4240 1510 4320 1520
rect 7000 1510 7200 1520
rect 8000 1510 8280 1520
rect 8640 1510 8680 1520
rect 9080 1510 9720 1520
rect 9840 1510 9880 1520
rect 2200 1500 2920 1510
rect 4240 1500 4320 1510
rect 7000 1500 7200 1510
rect 8000 1500 8280 1510
rect 8640 1500 8680 1510
rect 9080 1500 9720 1510
rect 9840 1500 9880 1510
rect 2200 1490 2880 1500
rect 4240 1490 4360 1500
rect 6960 1490 7240 1500
rect 8000 1490 8280 1500
rect 8600 1490 8720 1500
rect 9080 1490 9120 1500
rect 9200 1490 9680 1500
rect 9800 1490 9880 1500
rect 9920 1490 9990 1500
rect 2200 1480 2880 1490
rect 4240 1480 4360 1490
rect 6960 1480 7240 1490
rect 8000 1480 8280 1490
rect 8600 1480 8720 1490
rect 9080 1480 9120 1490
rect 9200 1480 9680 1490
rect 9800 1480 9880 1490
rect 9920 1480 9990 1490
rect 2200 1470 2880 1480
rect 4240 1470 4360 1480
rect 6960 1470 7240 1480
rect 8000 1470 8280 1480
rect 8600 1470 8720 1480
rect 9080 1470 9120 1480
rect 9200 1470 9680 1480
rect 9800 1470 9880 1480
rect 9920 1470 9990 1480
rect 2200 1460 2880 1470
rect 4240 1460 4360 1470
rect 6960 1460 7240 1470
rect 8000 1460 8280 1470
rect 8600 1460 8720 1470
rect 9080 1460 9120 1470
rect 9200 1460 9680 1470
rect 9800 1460 9880 1470
rect 9920 1460 9990 1470
rect 2240 1450 2840 1460
rect 4280 1450 4360 1460
rect 6880 1450 7240 1460
rect 8000 1450 8240 1460
rect 8600 1450 8680 1460
rect 9120 1450 9560 1460
rect 9800 1450 9990 1460
rect 2240 1440 2840 1450
rect 4280 1440 4360 1450
rect 6880 1440 7240 1450
rect 8000 1440 8240 1450
rect 8600 1440 8680 1450
rect 9120 1440 9560 1450
rect 9800 1440 9990 1450
rect 2240 1430 2840 1440
rect 4280 1430 4360 1440
rect 6880 1430 7240 1440
rect 8000 1430 8240 1440
rect 8600 1430 8680 1440
rect 9120 1430 9560 1440
rect 9800 1430 9990 1440
rect 2240 1420 2840 1430
rect 4280 1420 4360 1430
rect 6880 1420 7240 1430
rect 8000 1420 8240 1430
rect 8600 1420 8680 1430
rect 9120 1420 9560 1430
rect 9800 1420 9990 1430
rect 2280 1410 2800 1420
rect 4320 1410 4360 1420
rect 6840 1410 7280 1420
rect 8000 1410 8200 1420
rect 9120 1410 9200 1420
rect 9280 1410 9600 1420
rect 9760 1410 9920 1420
rect 2280 1400 2800 1410
rect 4320 1400 4360 1410
rect 6840 1400 7280 1410
rect 8000 1400 8200 1410
rect 9120 1400 9200 1410
rect 9280 1400 9600 1410
rect 9760 1400 9920 1410
rect 2280 1390 2800 1400
rect 4320 1390 4360 1400
rect 6840 1390 7280 1400
rect 8000 1390 8200 1400
rect 9120 1390 9200 1400
rect 9280 1390 9600 1400
rect 9760 1390 9920 1400
rect 2280 1380 2800 1390
rect 4320 1380 4360 1390
rect 6840 1380 7280 1390
rect 8000 1380 8200 1390
rect 9120 1380 9200 1390
rect 9280 1380 9600 1390
rect 9760 1380 9920 1390
rect 2360 1370 2760 1380
rect 4320 1370 4400 1380
rect 6840 1370 7280 1380
rect 8000 1370 8160 1380
rect 9120 1370 9160 1380
rect 9280 1370 9640 1380
rect 9760 1370 9800 1380
rect 9840 1370 9960 1380
rect 2360 1360 2760 1370
rect 4320 1360 4400 1370
rect 6840 1360 7280 1370
rect 8000 1360 8160 1370
rect 9120 1360 9160 1370
rect 9280 1360 9640 1370
rect 9760 1360 9800 1370
rect 9840 1360 9960 1370
rect 2360 1350 2760 1360
rect 4320 1350 4400 1360
rect 6840 1350 7280 1360
rect 8000 1350 8160 1360
rect 9120 1350 9160 1360
rect 9280 1350 9640 1360
rect 9760 1350 9800 1360
rect 9840 1350 9960 1360
rect 2360 1340 2760 1350
rect 4320 1340 4400 1350
rect 6840 1340 7280 1350
rect 8000 1340 8160 1350
rect 9120 1340 9160 1350
rect 9280 1340 9640 1350
rect 9760 1340 9800 1350
rect 9840 1340 9960 1350
rect 2440 1330 2680 1340
rect 3520 1330 3640 1340
rect 4280 1330 4400 1340
rect 6840 1330 7320 1340
rect 9280 1330 9640 1340
rect 9720 1330 9760 1340
rect 9840 1330 9960 1340
rect 2440 1320 2680 1330
rect 3520 1320 3640 1330
rect 4280 1320 4400 1330
rect 6840 1320 7320 1330
rect 9280 1320 9640 1330
rect 9720 1320 9760 1330
rect 9840 1320 9960 1330
rect 2440 1310 2680 1320
rect 3520 1310 3640 1320
rect 4280 1310 4400 1320
rect 6840 1310 7320 1320
rect 9280 1310 9640 1320
rect 9720 1310 9760 1320
rect 9840 1310 9960 1320
rect 2440 1300 2680 1310
rect 3520 1300 3640 1310
rect 4280 1300 4400 1310
rect 6840 1300 7320 1310
rect 9280 1300 9640 1310
rect 9720 1300 9760 1310
rect 9840 1300 9960 1310
rect 3520 1290 3720 1300
rect 4240 1290 4400 1300
rect 6840 1290 7280 1300
rect 9320 1290 9640 1300
rect 9840 1290 9960 1300
rect 3520 1280 3720 1290
rect 4240 1280 4400 1290
rect 6840 1280 7280 1290
rect 9320 1280 9640 1290
rect 9840 1280 9960 1290
rect 3520 1270 3720 1280
rect 4240 1270 4400 1280
rect 6840 1270 7280 1280
rect 9320 1270 9640 1280
rect 9840 1270 9960 1280
rect 3520 1260 3720 1270
rect 4240 1260 4400 1270
rect 6840 1260 7280 1270
rect 9320 1260 9640 1270
rect 9840 1260 9960 1270
rect 3680 1250 3760 1260
rect 4200 1250 4440 1260
rect 6840 1250 7320 1260
rect 9320 1250 9600 1260
rect 9680 1250 9720 1260
rect 9840 1250 9920 1260
rect 3680 1240 3760 1250
rect 4200 1240 4440 1250
rect 6840 1240 7320 1250
rect 9320 1240 9600 1250
rect 9680 1240 9720 1250
rect 9840 1240 9920 1250
rect 3680 1230 3760 1240
rect 4200 1230 4440 1240
rect 6840 1230 7320 1240
rect 9320 1230 9600 1240
rect 9680 1230 9720 1240
rect 9840 1230 9920 1240
rect 3680 1220 3760 1230
rect 4200 1220 4440 1230
rect 6840 1220 7320 1230
rect 9320 1220 9600 1230
rect 9680 1220 9720 1230
rect 9840 1220 9920 1230
rect 3720 1210 3800 1220
rect 4240 1210 4440 1220
rect 6840 1210 7320 1220
rect 9360 1210 9520 1220
rect 9560 1210 9600 1220
rect 9840 1210 9920 1220
rect 3720 1200 3800 1210
rect 4240 1200 4440 1210
rect 6840 1200 7320 1210
rect 9360 1200 9520 1210
rect 9560 1200 9600 1210
rect 9840 1200 9920 1210
rect 3720 1190 3800 1200
rect 4240 1190 4440 1200
rect 6840 1190 7320 1200
rect 9360 1190 9520 1200
rect 9560 1190 9600 1200
rect 9840 1190 9920 1200
rect 3720 1180 3800 1190
rect 4240 1180 4440 1190
rect 6840 1180 7320 1190
rect 9360 1180 9520 1190
rect 9560 1180 9600 1190
rect 9840 1180 9920 1190
rect 3760 1170 3880 1180
rect 4240 1170 4440 1180
rect 6720 1170 6760 1180
rect 6840 1170 7320 1180
rect 9400 1170 9520 1180
rect 9560 1170 9600 1180
rect 9640 1170 9680 1180
rect 9840 1170 9990 1180
rect 3760 1160 3880 1170
rect 4240 1160 4440 1170
rect 6720 1160 6760 1170
rect 6840 1160 7320 1170
rect 9400 1160 9520 1170
rect 9560 1160 9600 1170
rect 9640 1160 9680 1170
rect 9840 1160 9990 1170
rect 3760 1150 3880 1160
rect 4240 1150 4440 1160
rect 6720 1150 6760 1160
rect 6840 1150 7320 1160
rect 9400 1150 9520 1160
rect 9560 1150 9600 1160
rect 9640 1150 9680 1160
rect 9840 1150 9990 1160
rect 3760 1140 3880 1150
rect 4240 1140 4440 1150
rect 6720 1140 6760 1150
rect 6840 1140 7320 1150
rect 9400 1140 9520 1150
rect 9560 1140 9600 1150
rect 9640 1140 9680 1150
rect 9840 1140 9990 1150
rect 3760 1130 3920 1140
rect 4240 1130 4440 1140
rect 6640 1130 6760 1140
rect 6840 1130 7320 1140
rect 9400 1130 9520 1140
rect 9640 1130 9720 1140
rect 9960 1130 9990 1140
rect 3760 1120 3920 1130
rect 4240 1120 4440 1130
rect 6640 1120 6760 1130
rect 6840 1120 7320 1130
rect 9400 1120 9520 1130
rect 9640 1120 9720 1130
rect 9960 1120 9990 1130
rect 3760 1110 3920 1120
rect 4240 1110 4440 1120
rect 6640 1110 6760 1120
rect 6840 1110 7320 1120
rect 9400 1110 9520 1120
rect 9640 1110 9720 1120
rect 9960 1110 9990 1120
rect 3760 1100 3920 1110
rect 4240 1100 4440 1110
rect 6640 1100 6760 1110
rect 6840 1100 7320 1110
rect 9400 1100 9520 1110
rect 9640 1100 9720 1110
rect 9960 1100 9990 1110
rect 3840 1090 3960 1100
rect 4240 1090 4480 1100
rect 6560 1090 6800 1100
rect 6840 1090 7320 1100
rect 9440 1090 9520 1100
rect 9600 1090 9720 1100
rect 3840 1080 3960 1090
rect 4240 1080 4480 1090
rect 6560 1080 6800 1090
rect 6840 1080 7320 1090
rect 9440 1080 9520 1090
rect 9600 1080 9720 1090
rect 3840 1070 3960 1080
rect 4240 1070 4480 1080
rect 6560 1070 6800 1080
rect 6840 1070 7320 1080
rect 9440 1070 9520 1080
rect 9600 1070 9720 1080
rect 3840 1060 3960 1070
rect 4240 1060 4480 1070
rect 6560 1060 6800 1070
rect 6840 1060 7320 1070
rect 9440 1060 9520 1070
rect 9600 1060 9720 1070
rect 3880 1050 4040 1060
rect 4240 1050 4520 1060
rect 6560 1050 6800 1060
rect 6880 1050 7320 1060
rect 9160 1050 9240 1060
rect 9320 1050 9360 1060
rect 9440 1050 9520 1060
rect 9560 1050 9720 1060
rect 3880 1040 4040 1050
rect 4240 1040 4520 1050
rect 6560 1040 6800 1050
rect 6880 1040 7320 1050
rect 9160 1040 9240 1050
rect 9320 1040 9360 1050
rect 9440 1040 9520 1050
rect 9560 1040 9720 1050
rect 3880 1030 4040 1040
rect 4240 1030 4520 1040
rect 6560 1030 6800 1040
rect 6880 1030 7320 1040
rect 9160 1030 9240 1040
rect 9320 1030 9360 1040
rect 9440 1030 9520 1040
rect 9560 1030 9720 1040
rect 3880 1020 4040 1030
rect 4240 1020 4520 1030
rect 6560 1020 6800 1030
rect 6880 1020 7320 1030
rect 9160 1020 9240 1030
rect 9320 1020 9360 1030
rect 9440 1020 9520 1030
rect 9560 1020 9720 1030
rect 3880 1010 4120 1020
rect 4240 1010 4680 1020
rect 6520 1010 6800 1020
rect 6880 1010 7320 1020
rect 9160 1010 9480 1020
rect 9560 1010 9720 1020
rect 9840 1010 9920 1020
rect 9960 1010 9990 1020
rect 3880 1000 4120 1010
rect 4240 1000 4680 1010
rect 6520 1000 6800 1010
rect 6880 1000 7320 1010
rect 9160 1000 9480 1010
rect 9560 1000 9720 1010
rect 9840 1000 9920 1010
rect 9960 1000 9990 1010
rect 3880 990 4120 1000
rect 4240 990 4680 1000
rect 6520 990 6800 1000
rect 6880 990 7320 1000
rect 9160 990 9480 1000
rect 9560 990 9720 1000
rect 9840 990 9920 1000
rect 9960 990 9990 1000
rect 3880 980 4120 990
rect 4240 980 4680 990
rect 6520 980 6800 990
rect 6880 980 7320 990
rect 9160 980 9480 990
rect 9560 980 9720 990
rect 9840 980 9920 990
rect 9960 980 9990 990
rect 3880 970 4760 980
rect 6560 970 6800 980
rect 6880 970 7320 980
rect 9240 970 9480 980
rect 9520 970 9990 980
rect 3880 960 4760 970
rect 6560 960 6800 970
rect 6880 960 7320 970
rect 9240 960 9480 970
rect 9520 960 9990 970
rect 3880 950 4760 960
rect 6560 950 6800 960
rect 6880 950 7320 960
rect 9240 950 9480 960
rect 9520 950 9990 960
rect 3880 940 4760 950
rect 6560 940 6800 950
rect 6880 940 7320 950
rect 9240 940 9480 950
rect 9520 940 9990 950
rect 3880 930 4800 940
rect 6560 930 6800 940
rect 6880 930 7320 940
rect 9200 930 9440 940
rect 9520 930 9990 940
rect 3880 920 4800 930
rect 6560 920 6800 930
rect 6880 920 7320 930
rect 9200 920 9440 930
rect 9520 920 9990 930
rect 3880 910 4800 920
rect 6560 910 6800 920
rect 6880 910 7320 920
rect 9200 910 9440 920
rect 9520 910 9990 920
rect 3880 900 4800 910
rect 6560 900 6800 910
rect 6880 900 7320 910
rect 9200 900 9440 910
rect 9520 900 9990 910
rect 4040 890 4840 900
rect 6560 890 6800 900
rect 6880 890 7280 900
rect 9200 890 9440 900
rect 9480 890 9520 900
rect 9560 890 9990 900
rect 4040 880 4840 890
rect 6560 880 6800 890
rect 6880 880 7280 890
rect 9200 880 9440 890
rect 9480 880 9520 890
rect 9560 880 9990 890
rect 4040 870 4840 880
rect 6560 870 6800 880
rect 6880 870 7280 880
rect 9200 870 9440 880
rect 9480 870 9520 880
rect 9560 870 9990 880
rect 4040 860 4840 870
rect 6560 860 6800 870
rect 6880 860 7280 870
rect 9200 860 9440 870
rect 9480 860 9520 870
rect 9560 860 9990 870
rect 2440 850 2480 860
rect 2520 850 2560 860
rect 4040 850 4240 860
rect 4280 850 4880 860
rect 6560 850 6840 860
rect 6880 850 7280 860
rect 9200 850 9400 860
rect 9480 850 9990 860
rect 2440 840 2480 850
rect 2520 840 2560 850
rect 4040 840 4240 850
rect 4280 840 4880 850
rect 6560 840 6840 850
rect 6880 840 7280 850
rect 9200 840 9400 850
rect 9480 840 9990 850
rect 2440 830 2480 840
rect 2520 830 2560 840
rect 4040 830 4240 840
rect 4280 830 4880 840
rect 6560 830 6840 840
rect 6880 830 7280 840
rect 9200 830 9400 840
rect 9480 830 9990 840
rect 2440 820 2480 830
rect 2520 820 2560 830
rect 4040 820 4240 830
rect 4280 820 4880 830
rect 6560 820 6840 830
rect 6880 820 7280 830
rect 9200 820 9400 830
rect 9480 820 9990 830
rect 2360 810 2440 820
rect 2480 810 2560 820
rect 4040 810 4280 820
rect 4360 810 4880 820
rect 6600 810 6840 820
rect 6880 810 7280 820
rect 9200 810 9360 820
rect 9440 810 9990 820
rect 2360 800 2440 810
rect 2480 800 2560 810
rect 4040 800 4280 810
rect 4360 800 4880 810
rect 6600 800 6840 810
rect 6880 800 7280 810
rect 9200 800 9360 810
rect 9440 800 9990 810
rect 2360 790 2440 800
rect 2480 790 2560 800
rect 4040 790 4280 800
rect 4360 790 4880 800
rect 6600 790 6840 800
rect 6880 790 7280 800
rect 9200 790 9360 800
rect 9440 790 9990 800
rect 2360 780 2440 790
rect 2480 780 2560 790
rect 4040 780 4280 790
rect 4360 780 4880 790
rect 6600 780 6840 790
rect 6880 780 7280 790
rect 9200 780 9360 790
rect 9440 780 9990 790
rect 2320 770 2480 780
rect 3720 770 3760 780
rect 3800 770 3840 780
rect 4040 770 4320 780
rect 4360 770 4920 780
rect 6600 770 6840 780
rect 6880 770 7280 780
rect 9240 770 9360 780
rect 9400 770 9990 780
rect 2320 760 2480 770
rect 3720 760 3760 770
rect 3800 760 3840 770
rect 4040 760 4320 770
rect 4360 760 4920 770
rect 6600 760 6840 770
rect 6880 760 7280 770
rect 9240 760 9360 770
rect 9400 760 9990 770
rect 2320 750 2480 760
rect 3720 750 3760 760
rect 3800 750 3840 760
rect 4040 750 4320 760
rect 4360 750 4920 760
rect 6600 750 6840 760
rect 6880 750 7280 760
rect 9240 750 9360 760
rect 9400 750 9990 760
rect 2320 740 2480 750
rect 3720 740 3760 750
rect 3800 740 3840 750
rect 4040 740 4320 750
rect 4360 740 4920 750
rect 6600 740 6840 750
rect 6880 740 7280 750
rect 9240 740 9360 750
rect 9400 740 9990 750
rect 2240 730 2400 740
rect 3480 730 3920 740
rect 4200 730 4720 740
rect 4800 730 4920 740
rect 6600 730 6840 740
rect 6920 730 7280 740
rect 9240 730 9320 740
rect 9400 730 9990 740
rect 2240 720 2400 730
rect 3480 720 3920 730
rect 4200 720 4720 730
rect 4800 720 4920 730
rect 6600 720 6840 730
rect 6920 720 7280 730
rect 9240 720 9320 730
rect 9400 720 9990 730
rect 2240 710 2400 720
rect 3480 710 3920 720
rect 4200 710 4720 720
rect 4800 710 4920 720
rect 6600 710 6840 720
rect 6920 710 7280 720
rect 9240 710 9320 720
rect 9400 710 9990 720
rect 2240 700 2400 710
rect 3480 700 3920 710
rect 4200 700 4720 710
rect 4800 700 4920 710
rect 6600 700 6840 710
rect 6920 700 7280 710
rect 9240 700 9320 710
rect 9400 700 9990 710
rect 2240 690 2320 700
rect 3360 690 4040 700
rect 4200 690 4720 700
rect 4840 690 4920 700
rect 6640 690 6840 700
rect 6920 690 7240 700
rect 9240 690 9320 700
rect 9360 690 9990 700
rect 2240 680 2320 690
rect 3360 680 4040 690
rect 4200 680 4720 690
rect 4840 680 4920 690
rect 6640 680 6840 690
rect 6920 680 7240 690
rect 9240 680 9320 690
rect 9360 680 9990 690
rect 2240 670 2320 680
rect 3360 670 4040 680
rect 4200 670 4720 680
rect 4840 670 4920 680
rect 6640 670 6840 680
rect 6920 670 7240 680
rect 9240 670 9320 680
rect 9360 670 9990 680
rect 2240 660 2320 670
rect 3360 660 4040 670
rect 4200 660 4720 670
rect 4840 660 4920 670
rect 6640 660 6840 670
rect 6920 660 7240 670
rect 9240 660 9320 670
rect 9360 660 9990 670
rect 3280 650 4080 660
rect 4120 650 4680 660
rect 4840 650 4920 660
rect 6680 650 6840 660
rect 6960 650 7240 660
rect 9240 650 9280 660
rect 9360 650 9600 660
rect 9720 650 9990 660
rect 3280 640 4080 650
rect 4120 640 4680 650
rect 4840 640 4920 650
rect 6680 640 6840 650
rect 6960 640 7240 650
rect 9240 640 9280 650
rect 9360 640 9600 650
rect 9720 640 9990 650
rect 3280 630 4080 640
rect 4120 630 4680 640
rect 4840 630 4920 640
rect 6680 630 6840 640
rect 6960 630 7240 640
rect 9240 630 9280 640
rect 9360 630 9600 640
rect 9720 630 9990 640
rect 3280 620 4080 630
rect 4120 620 4680 630
rect 4840 620 4920 630
rect 6680 620 6840 630
rect 6960 620 7240 630
rect 9240 620 9280 630
rect 9360 620 9600 630
rect 9720 620 9990 630
rect 480 610 560 620
rect 3200 610 4040 620
rect 4080 610 4520 620
rect 4560 610 4680 620
rect 4800 610 4920 620
rect 6720 610 6880 620
rect 7000 610 7200 620
rect 9320 610 9990 620
rect 480 600 560 610
rect 3200 600 4040 610
rect 4080 600 4520 610
rect 4560 600 4680 610
rect 4800 600 4920 610
rect 6720 600 6880 610
rect 7000 600 7200 610
rect 9320 600 9990 610
rect 480 590 560 600
rect 3200 590 4040 600
rect 4080 590 4520 600
rect 4560 590 4680 600
rect 4800 590 4920 600
rect 6720 590 6880 600
rect 7000 590 7200 600
rect 9320 590 9990 600
rect 480 580 560 590
rect 3200 580 4040 590
rect 4080 580 4520 590
rect 4560 580 4680 590
rect 4800 580 4920 590
rect 6720 580 6880 590
rect 7000 580 7200 590
rect 9320 580 9990 590
rect 360 570 600 580
rect 3120 570 4360 580
rect 4560 570 4640 580
rect 4800 570 4840 580
rect 4880 570 4920 580
rect 6720 570 6880 580
rect 7040 570 7160 580
rect 9320 570 9990 580
rect 360 560 600 570
rect 3120 560 4360 570
rect 4560 560 4640 570
rect 4800 560 4840 570
rect 4880 560 4920 570
rect 6720 560 6880 570
rect 7040 560 7160 570
rect 9320 560 9990 570
rect 360 550 600 560
rect 3120 550 4360 560
rect 4560 550 4640 560
rect 4800 550 4840 560
rect 4880 550 4920 560
rect 6720 550 6880 560
rect 7040 550 7160 560
rect 9320 550 9990 560
rect 360 540 600 550
rect 3120 540 4360 550
rect 4560 540 4640 550
rect 4800 540 4840 550
rect 4880 540 4920 550
rect 6720 540 6880 550
rect 7040 540 7160 550
rect 9320 540 9990 550
rect 360 530 520 540
rect 1280 530 1480 540
rect 3000 530 4240 540
rect 4800 530 4960 540
rect 6760 530 6880 540
rect 7080 530 7120 540
rect 9280 530 9920 540
rect 360 520 520 530
rect 1280 520 1480 530
rect 3000 520 4240 530
rect 4800 520 4960 530
rect 6760 520 6880 530
rect 7080 520 7120 530
rect 9280 520 9920 530
rect 360 510 520 520
rect 1280 510 1480 520
rect 3000 510 4240 520
rect 4800 510 4960 520
rect 6760 510 6880 520
rect 7080 510 7120 520
rect 9280 510 9920 520
rect 360 500 520 510
rect 1280 500 1480 510
rect 3000 500 4240 510
rect 4800 500 4960 510
rect 6760 500 6880 510
rect 7080 500 7120 510
rect 9280 500 9920 510
rect 400 490 440 500
rect 1200 490 1520 500
rect 2880 490 4200 500
rect 4800 490 4880 500
rect 4920 490 4960 500
rect 6760 490 6880 500
rect 9240 490 9880 500
rect 9960 490 9990 500
rect 400 480 440 490
rect 1200 480 1520 490
rect 2880 480 4200 490
rect 4800 480 4880 490
rect 4920 480 4960 490
rect 6760 480 6880 490
rect 9240 480 9880 490
rect 9960 480 9990 490
rect 400 470 440 480
rect 1200 470 1520 480
rect 2880 470 4200 480
rect 4800 470 4880 480
rect 4920 470 4960 480
rect 6760 470 6880 480
rect 9240 470 9880 480
rect 9960 470 9990 480
rect 400 460 440 470
rect 1200 460 1520 470
rect 2880 460 4200 470
rect 4800 460 4880 470
rect 4920 460 4960 470
rect 6760 460 6880 470
rect 9240 460 9880 470
rect 9960 460 9990 470
rect 120 450 280 460
rect 1160 450 1560 460
rect 2040 450 2240 460
rect 2720 450 4160 460
rect 4760 450 4880 460
rect 4920 450 4960 460
rect 9240 450 9280 460
rect 9360 450 9990 460
rect 120 440 280 450
rect 1160 440 1560 450
rect 2040 440 2240 450
rect 2720 440 4160 450
rect 4760 440 4880 450
rect 4920 440 4960 450
rect 9240 440 9280 450
rect 9360 440 9990 450
rect 120 430 280 440
rect 1160 430 1560 440
rect 2040 430 2240 440
rect 2720 430 4160 440
rect 4760 430 4880 440
rect 4920 430 4960 440
rect 9240 430 9280 440
rect 9360 430 9990 440
rect 120 420 280 430
rect 1160 420 1560 430
rect 2040 420 2240 430
rect 2720 420 4160 430
rect 4760 420 4880 430
rect 4920 420 4960 430
rect 9240 420 9280 430
rect 9360 420 9990 430
rect 80 410 280 420
rect 1120 410 4160 420
rect 4760 410 4960 420
rect 9200 410 9280 420
rect 9400 410 9990 420
rect 80 400 280 410
rect 1120 400 4160 410
rect 4760 400 4960 410
rect 9200 400 9280 410
rect 9400 400 9990 410
rect 80 390 280 400
rect 1120 390 4160 400
rect 4760 390 4960 400
rect 9200 390 9280 400
rect 9400 390 9990 400
rect 80 380 280 390
rect 1120 380 4160 390
rect 4760 380 4960 390
rect 9200 380 9280 390
rect 9400 380 9990 390
rect 80 370 280 380
rect 1080 370 4120 380
rect 4760 370 4920 380
rect 9200 370 9240 380
rect 9440 370 9990 380
rect 80 360 280 370
rect 1080 360 4120 370
rect 4760 360 4920 370
rect 9200 360 9240 370
rect 9440 360 9990 370
rect 80 350 280 360
rect 1080 350 4120 360
rect 4760 350 4920 360
rect 9200 350 9240 360
rect 9440 350 9990 360
rect 80 340 280 350
rect 1080 340 4120 350
rect 4760 340 4920 350
rect 9200 340 9240 350
rect 9440 340 9990 350
rect 40 330 80 340
rect 120 330 240 340
rect 1040 330 4080 340
rect 9160 330 9200 340
rect 9440 330 9990 340
rect 40 320 80 330
rect 120 320 240 330
rect 1040 320 4080 330
rect 9160 320 9200 330
rect 9440 320 9990 330
rect 40 310 80 320
rect 120 310 240 320
rect 1040 310 4080 320
rect 9160 310 9200 320
rect 9440 310 9990 320
rect 40 300 80 310
rect 120 300 240 310
rect 1040 300 4080 310
rect 9160 300 9200 310
rect 9440 300 9990 310
rect 520 290 560 300
rect 1040 290 4080 300
rect 9120 290 9200 300
rect 9480 290 9990 300
rect 520 280 560 290
rect 1040 280 4080 290
rect 9120 280 9200 290
rect 9480 280 9990 290
rect 520 270 560 280
rect 1040 270 4080 280
rect 9120 270 9200 280
rect 9480 270 9990 280
rect 520 260 560 270
rect 1040 260 4080 270
rect 9120 260 9200 270
rect 9480 260 9990 270
rect 1040 250 4080 260
rect 4960 250 5000 260
rect 9120 250 9160 260
rect 9480 250 9800 260
rect 9840 250 9990 260
rect 1040 240 4080 250
rect 4960 240 5000 250
rect 9120 240 9160 250
rect 9480 240 9800 250
rect 9840 240 9990 250
rect 1040 230 4080 240
rect 4960 230 5000 240
rect 9120 230 9160 240
rect 9480 230 9800 240
rect 9840 230 9990 240
rect 1040 220 4080 230
rect 4960 220 5000 230
rect 9120 220 9160 230
rect 9480 220 9800 230
rect 9840 220 9990 230
rect 1040 210 4120 220
rect 4920 210 5000 220
rect 9080 210 9120 220
rect 9360 210 9720 220
rect 1040 200 4120 210
rect 4920 200 5000 210
rect 9080 200 9120 210
rect 9360 200 9720 210
rect 1040 190 4120 200
rect 4920 190 5000 200
rect 9080 190 9120 200
rect 9360 190 9720 200
rect 1040 180 4120 190
rect 4920 180 5000 190
rect 9080 180 9120 190
rect 9360 180 9720 190
rect 1040 170 4160 180
rect 4960 170 5000 180
rect 9080 170 9120 180
rect 9360 170 9720 180
rect 1040 160 4160 170
rect 4960 160 5000 170
rect 9080 160 9120 170
rect 9360 160 9720 170
rect 1040 150 4160 160
rect 4960 150 5000 160
rect 9080 150 9120 160
rect 9360 150 9720 160
rect 1040 140 4160 150
rect 4960 140 5000 150
rect 9080 140 9120 150
rect 9360 140 9720 150
rect 1040 130 4200 140
rect 4960 130 5000 140
rect 8840 130 8920 140
rect 9400 130 9720 140
rect 1040 120 4200 130
rect 4960 120 5000 130
rect 8840 120 8920 130
rect 9400 120 9720 130
rect 1040 110 4200 120
rect 4960 110 5000 120
rect 8840 110 8920 120
rect 9400 110 9720 120
rect 1040 100 4200 110
rect 4960 100 5000 110
rect 8840 100 8920 110
rect 9400 100 9720 110
rect 1040 90 4240 100
rect 4960 90 5040 100
rect 8800 90 8920 100
rect 9080 90 9120 100
rect 9480 90 9560 100
rect 9600 90 9680 100
rect 1040 80 4240 90
rect 4960 80 5040 90
rect 8800 80 8920 90
rect 9080 80 9120 90
rect 9480 80 9560 90
rect 9600 80 9680 90
rect 1040 70 4240 80
rect 4960 70 5040 80
rect 8800 70 8920 80
rect 9080 70 9120 80
rect 9480 70 9560 80
rect 9600 70 9680 80
rect 1040 60 4240 70
rect 4960 60 5040 70
rect 8800 60 8920 70
rect 9080 60 9120 70
rect 9480 60 9560 70
rect 9600 60 9680 70
rect 0 50 40 60
rect 1040 50 4320 60
rect 4960 50 5040 60
rect 8760 50 8920 60
rect 9040 50 9080 60
rect 9120 50 9160 60
rect 0 40 40 50
rect 1040 40 4320 50
rect 4960 40 5040 50
rect 8760 40 8920 50
rect 9040 40 9080 50
rect 9120 40 9160 50
rect 0 30 40 40
rect 1040 30 4320 40
rect 4960 30 5040 40
rect 8760 30 8920 40
rect 9040 30 9080 40
rect 9120 30 9160 40
rect 0 20 40 30
rect 1040 20 4320 30
rect 4960 20 5040 30
rect 8760 20 8920 30
rect 9040 20 9080 30
rect 9120 20 9160 30
rect 1040 10 4360 20
rect 4960 10 5040 20
rect 8720 10 8880 20
rect 9040 10 9080 20
rect 9120 10 9160 20
rect 9960 10 9990 20
rect 1040 0 4360 10
rect 4960 0 5040 10
rect 8720 0 8880 10
rect 9040 0 9080 10
rect 9120 0 9160 10
rect 9960 0 9990 10
<< end >>
